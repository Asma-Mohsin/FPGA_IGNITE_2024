magic
tech sky130A
magscale 1 2
timestamp 1732544675
<< viali >>
rect 1869 43401 1903 43435
rect 2789 43401 2823 43435
rect 3157 43401 3191 43435
rect 4629 43401 4663 43435
rect 5549 43401 5583 43435
rect 6101 43401 6135 43435
rect 6377 43401 6411 43435
rect 6837 43401 6871 43435
rect 7389 43401 7423 43435
rect 7757 43401 7791 43435
rect 8309 43401 8343 43435
rect 8677 43401 8711 43435
rect 9229 43401 9263 43435
rect 9781 43401 9815 43435
rect 10517 43401 10551 43435
rect 15209 43401 15243 43435
rect 20085 43401 20119 43435
rect 21005 43401 21039 43435
rect 22017 43401 22051 43435
rect 22385 43401 22419 43435
rect 23489 43401 23523 43435
rect 4537 43333 4571 43367
rect 6745 43333 6779 43367
rect 8033 43333 8067 43367
rect 12449 43333 12483 43367
rect 12817 43333 12851 43367
rect 13737 43333 13771 43367
rect 14197 43333 14231 43367
rect 14749 43333 14783 43367
rect 15117 43333 15151 43367
rect 15577 43333 15611 43367
rect 16313 43333 16347 43367
rect 16773 43333 16807 43367
rect 1593 43265 1627 43299
rect 1777 43265 1811 43299
rect 2513 43265 2547 43299
rect 3065 43265 3099 43299
rect 3985 43265 4019 43299
rect 5273 43265 5307 43299
rect 5917 43265 5951 43299
rect 6561 43265 6595 43299
rect 7205 43265 7239 43299
rect 7573 43265 7607 43299
rect 8493 43265 8527 43299
rect 9045 43265 9079 43299
rect 9505 43265 9539 43299
rect 9965 43265 9999 43299
rect 10333 43265 10367 43299
rect 10701 43265 10735 43299
rect 11069 43265 11103 43299
rect 11529 43265 11563 43299
rect 12081 43265 12115 43299
rect 15853 43265 15887 43299
rect 17509 43265 17543 43299
rect 17785 43265 17819 43299
rect 18061 43265 18095 43299
rect 18337 43265 18371 43299
rect 18613 43265 18647 43299
rect 18889 43265 18923 43299
rect 19441 43265 19475 43299
rect 19717 43265 19751 43299
rect 19901 43265 19935 43299
rect 20361 43265 20395 43299
rect 20913 43265 20947 43299
rect 21373 43265 21407 43299
rect 21833 43265 21867 43299
rect 22293 43265 22327 43299
rect 22845 43265 22879 43299
rect 23397 43265 23431 43299
rect 23949 43265 23983 43299
rect 16497 43197 16531 43231
rect 20637 43197 20671 43231
rect 3801 43129 3835 43163
rect 10149 43129 10183 43163
rect 14933 43129 14967 43163
rect 18153 43129 18187 43163
rect 18705 43129 18739 43163
rect 21557 43129 21591 43163
rect 1409 43061 1443 43095
rect 4261 43061 4295 43095
rect 10885 43061 10919 43095
rect 11253 43061 11287 43095
rect 11713 43061 11747 43095
rect 12265 43061 12299 43095
rect 12541 43061 12575 43095
rect 12909 43061 12943 43095
rect 13829 43061 13863 43095
rect 14289 43061 14323 43095
rect 15669 43061 15703 43095
rect 16037 43061 16071 43095
rect 16865 43061 16899 43095
rect 17325 43061 17359 43095
rect 17601 43061 17635 43095
rect 17877 43061 17911 43095
rect 18429 43061 18463 43095
rect 19257 43061 19291 43095
rect 19533 43061 19567 43095
rect 22937 43061 22971 43095
rect 24133 43061 24167 43095
rect 2237 42857 2271 42891
rect 3341 42857 3375 42891
rect 6101 42857 6135 42891
rect 6837 42857 6871 42891
rect 7389 42857 7423 42891
rect 10333 42857 10367 42891
rect 10609 42857 10643 42891
rect 18889 42857 18923 42891
rect 13185 42789 13219 42823
rect 21097 42789 21131 42823
rect 1777 42721 1811 42755
rect 4353 42721 4387 42755
rect 5365 42721 5399 42755
rect 8677 42721 8711 42755
rect 9781 42721 9815 42755
rect 22937 42721 22971 42755
rect 23489 42721 23523 42755
rect 2145 42653 2179 42687
rect 4537 42653 4571 42687
rect 5089 42653 5123 42687
rect 5549 42653 5583 42687
rect 7757 42653 7791 42687
rect 8401 42653 8435 42687
rect 9137 42653 9171 42687
rect 10057 42653 10091 42687
rect 10517 42653 10551 42687
rect 10793 42653 10827 42687
rect 11621 42653 11655 42687
rect 11897 42653 11931 42687
rect 12725 42653 12759 42687
rect 13001 42653 13035 42687
rect 14105 42653 14139 42687
rect 14381 42653 14415 42687
rect 14657 42653 14691 42687
rect 15301 42653 15335 42687
rect 15577 42653 15611 42687
rect 16497 42653 16531 42687
rect 16589 42653 16623 42687
rect 17141 42653 17175 42687
rect 17417 42653 17451 42687
rect 17693 42653 17727 42687
rect 17969 42653 18003 42687
rect 18245 42653 18279 42687
rect 18521 42653 18555 42687
rect 18797 42649 18831 42683
rect 19073 42653 19107 42687
rect 21281 42653 21315 42687
rect 21925 42653 21959 42687
rect 22477 42653 22511 42687
rect 24133 42653 24167 42687
rect 1501 42585 1535 42619
rect 2697 42585 2731 42619
rect 3249 42585 3283 42619
rect 4077 42585 4111 42619
rect 6009 42585 6043 42619
rect 6745 42585 6779 42619
rect 7297 42585 7331 42619
rect 9505 42585 9539 42619
rect 19257 42585 19291 42619
rect 21557 42585 21591 42619
rect 22109 42585 22143 42619
rect 22661 42585 22695 42619
rect 23213 42585 23247 42619
rect 23765 42585 23799 42619
rect 2789 42517 2823 42551
rect 4721 42517 4755 42551
rect 5733 42517 5767 42551
rect 7941 42517 7975 42551
rect 8953 42517 8987 42551
rect 10241 42517 10275 42551
rect 11805 42517 11839 42551
rect 12081 42517 12115 42551
rect 12909 42517 12943 42551
rect 14289 42517 14323 42551
rect 14565 42517 14599 42551
rect 14841 42517 14875 42551
rect 15485 42517 15519 42551
rect 15761 42517 15795 42551
rect 16313 42517 16347 42551
rect 16773 42517 16807 42551
rect 16957 42517 16991 42551
rect 17233 42517 17267 42551
rect 17509 42517 17543 42551
rect 17785 42517 17819 42551
rect 18061 42517 18095 42551
rect 18337 42517 18371 42551
rect 18613 42517 18647 42551
rect 20545 42517 20579 42551
rect 1593 42313 1627 42347
rect 2513 42313 2547 42347
rect 3433 42313 3467 42347
rect 3709 42313 3743 42347
rect 4169 42313 4203 42347
rect 4997 42313 5031 42347
rect 6009 42313 6043 42347
rect 8493 42313 8527 42347
rect 8953 42313 8987 42347
rect 9229 42313 9263 42347
rect 9689 42313 9723 42347
rect 9965 42313 9999 42347
rect 19717 42313 19751 42347
rect 19993 42313 20027 42347
rect 20821 42313 20855 42347
rect 21833 42313 21867 42347
rect 23121 42313 23155 42347
rect 23673 42313 23707 42347
rect 1501 42245 1535 42279
rect 16773 42245 16807 42279
rect 17141 42245 17175 42279
rect 17509 42245 17543 42279
rect 17877 42245 17911 42279
rect 18245 42245 18279 42279
rect 18613 42245 18647 42279
rect 18981 42245 19015 42279
rect 19349 42245 19383 42279
rect 2053 42177 2087 42211
rect 2697 42177 2731 42211
rect 2789 42177 2823 42211
rect 3617 42177 3651 42211
rect 3893 42177 3927 42211
rect 3985 42177 4019 42211
rect 4721 42177 4755 42211
rect 4813 42177 4847 42211
rect 5457 42177 5491 42211
rect 5917 42177 5951 42211
rect 6193 42177 6227 42211
rect 6561 42177 6595 42211
rect 7113 42177 7147 42211
rect 7389 42177 7423 42211
rect 7665 42177 7699 42211
rect 7941 42177 7975 42211
rect 8217 42177 8251 42211
rect 8401 42177 8435 42211
rect 9137 42177 9171 42211
rect 9413 42177 9447 42211
rect 9873 42177 9907 42211
rect 10149 42177 10183 42211
rect 16221 42177 16255 42211
rect 19901 42177 19935 42211
rect 20177 42177 20211 42211
rect 20453 42177 20487 42211
rect 20729 42177 20763 42211
rect 21005 42177 21039 42211
rect 21281 42177 21315 42211
rect 21649 42177 21683 42211
rect 22017 42177 22051 42211
rect 22293 42177 22327 42211
rect 22845 42177 22879 42211
rect 23397 42177 23431 42211
rect 24041 42177 24075 42211
rect 22569 42109 22603 42143
rect 2973 42041 3007 42075
rect 4537 42041 4571 42075
rect 6377 42041 6411 42075
rect 16405 42041 16439 42075
rect 17325 42041 17359 42075
rect 18061 42041 18095 42075
rect 18429 42041 18463 42075
rect 20545 42041 20579 42075
rect 2145 41973 2179 42007
rect 5733 41973 5767 42007
rect 6929 41973 6963 42007
rect 7205 41973 7239 42007
rect 7481 41973 7515 42007
rect 7757 41973 7791 42007
rect 8033 41973 8067 42007
rect 16865 41973 16899 42007
rect 17601 41973 17635 42007
rect 18705 41973 18739 42007
rect 19073 41973 19107 42007
rect 19441 41973 19475 42007
rect 20269 41973 20303 42007
rect 24317 41973 24351 42007
rect 1593 41769 1627 41803
rect 2697 41769 2731 41803
rect 2881 41769 2915 41803
rect 3157 41769 3191 41803
rect 3433 41769 3467 41803
rect 3801 41769 3835 41803
rect 4445 41769 4479 41803
rect 4721 41769 4755 41803
rect 5457 41769 5491 41803
rect 5825 41769 5859 41803
rect 6193 41769 6227 41803
rect 7205 41769 7239 41803
rect 7573 41769 7607 41803
rect 8401 41769 8435 41803
rect 17969 41769 18003 41803
rect 18429 41769 18463 41803
rect 18797 41769 18831 41803
rect 19625 41769 19659 41803
rect 20269 41769 20303 41803
rect 20729 41769 20763 41803
rect 21189 41769 21223 41803
rect 23029 41769 23063 41803
rect 24133 41769 24167 41803
rect 8125 41701 8159 41735
rect 19349 41701 19383 41735
rect 19993 41701 20027 41735
rect 23581 41701 23615 41735
rect 9689 41633 9723 41667
rect 1501 41565 1535 41599
rect 2513 41565 2547 41599
rect 3065 41565 3099 41599
rect 3341 41565 3375 41599
rect 3617 41565 3651 41599
rect 3985 41565 4019 41599
rect 4261 41565 4295 41599
rect 4629 41565 4663 41599
rect 4905 41565 4939 41599
rect 5365 41565 5399 41599
rect 5641 41565 5675 41599
rect 6009 41565 6043 41599
rect 6377 41565 6411 41599
rect 6745 41565 6779 41599
rect 7389 41565 7423 41599
rect 7757 41565 7791 41599
rect 8033 41565 8067 41599
rect 8309 41565 8343 41599
rect 8585 41565 8619 41599
rect 9963 41565 9997 41599
rect 18153 41565 18187 41599
rect 18337 41565 18371 41599
rect 18981 41565 19015 41599
rect 19533 41565 19567 41599
rect 19809 41565 19843 41599
rect 20177 41565 20211 41599
rect 20453 41565 20487 41599
rect 20545 41561 20579 41595
rect 21097 41565 21131 41599
rect 21373 41565 21407 41599
rect 21649 41565 21683 41599
rect 21925 41565 21959 41599
rect 22753 41565 22787 41599
rect 23305 41565 23339 41599
rect 2053 41497 2087 41531
rect 22201 41497 22235 41531
rect 23857 41497 23891 41531
rect 2145 41429 2179 41463
rect 4077 41429 4111 41463
rect 5181 41429 5215 41463
rect 6561 41429 6595 41463
rect 7113 41429 7147 41463
rect 7849 41429 7883 41463
rect 10701 41429 10735 41463
rect 20913 41429 20947 41463
rect 21465 41429 21499 41463
rect 21741 41429 21775 41463
rect 22477 41429 22511 41463
rect 2513 41225 2547 41259
rect 2789 41225 2823 41259
rect 3065 41225 3099 41259
rect 7757 41225 7791 41259
rect 19533 41225 19567 41259
rect 20085 41225 20119 41259
rect 20637 41225 20671 41259
rect 20913 41225 20947 41259
rect 21465 41225 21499 41259
rect 22385 41225 22419 41259
rect 23121 41225 23155 41259
rect 24225 41225 24259 41259
rect 2237 41157 2271 41191
rect 1409 41089 1443 41123
rect 2697 41089 2731 41123
rect 2973 41089 3007 41123
rect 3249 41089 3283 41123
rect 3799 41089 3833 41123
rect 5179 41089 5213 41123
rect 7941 41089 7975 41123
rect 8843 41119 8877 41153
rect 10331 41089 10365 41123
rect 19257 41089 19291 41123
rect 19717 41089 19751 41123
rect 19993 41089 20027 41123
rect 20269 41089 20303 41123
rect 20545 41089 20579 41123
rect 20821 41089 20855 41123
rect 21097 41089 21131 41123
rect 21373 41089 21407 41123
rect 21649 41089 21683 41123
rect 22017 41089 22051 41123
rect 22293 41089 22327 41123
rect 22569 41089 22603 41123
rect 22845 41089 22879 41123
rect 23397 41089 23431 41123
rect 23949 41089 23983 41123
rect 3525 41021 3559 41055
rect 4905 41021 4939 41055
rect 8585 41021 8619 41055
rect 10057 41021 10091 41055
rect 20361 40953 20395 40987
rect 21189 40953 21223 40987
rect 22109 40953 22143 40987
rect 4537 40885 4571 40919
rect 5917 40885 5951 40919
rect 9597 40885 9631 40919
rect 11069 40885 11103 40919
rect 19073 40885 19107 40919
rect 19809 40885 19843 40919
rect 21833 40885 21867 40919
rect 23673 40885 23707 40919
rect 3433 40681 3467 40715
rect 20545 40681 20579 40715
rect 20821 40681 20855 40715
rect 21373 40681 21407 40715
rect 21649 40681 21683 40715
rect 22201 40681 22235 40715
rect 22753 40681 22787 40715
rect 23029 40681 23063 40715
rect 23489 40681 23523 40715
rect 10517 40613 10551 40647
rect 19993 40613 20027 40647
rect 20269 40613 20303 40647
rect 22477 40613 22511 40647
rect 3801 40545 3835 40579
rect 10057 40545 10091 40579
rect 10910 40545 10944 40579
rect 11069 40545 11103 40579
rect 3617 40477 3651 40511
rect 4075 40477 4109 40511
rect 5549 40477 5583 40511
rect 5823 40477 5857 40511
rect 6929 40477 6963 40511
rect 7203 40477 7237 40511
rect 9873 40477 9907 40511
rect 10793 40477 10827 40511
rect 11805 40477 11839 40511
rect 12063 40447 12097 40481
rect 13369 40477 13403 40511
rect 19349 40477 19383 40511
rect 19809 40477 19843 40511
rect 20177 40477 20211 40511
rect 20453 40477 20487 40511
rect 20729 40477 20763 40511
rect 21005 40477 21039 40511
rect 21281 40477 21315 40511
rect 21557 40477 21591 40511
rect 21833 40477 21867 40511
rect 22109 40477 22143 40511
rect 22385 40477 22419 40511
rect 22661 40477 22695 40511
rect 22937 40477 22971 40511
rect 23213 40477 23247 40511
rect 23673 40477 23707 40511
rect 1409 40409 1443 40443
rect 2237 40409 2271 40443
rect 2421 40409 2455 40443
rect 3249 40409 3283 40443
rect 23857 40409 23891 40443
rect 24225 40409 24259 40443
rect 4813 40341 4847 40375
rect 6561 40341 6595 40375
rect 7941 40341 7975 40375
rect 11713 40341 11747 40375
rect 12817 40341 12851 40375
rect 19441 40341 19475 40375
rect 19625 40341 19659 40375
rect 21097 40341 21131 40375
rect 21925 40341 21959 40375
rect 7481 40137 7515 40171
rect 19809 40137 19843 40171
rect 20085 40137 20119 40171
rect 20913 40137 20947 40171
rect 21189 40137 21223 40171
rect 1685 40069 1719 40103
rect 7849 40069 7883 40103
rect 8585 40069 8619 40103
rect 9137 40069 9171 40103
rect 9413 40069 9447 40103
rect 9505 40069 9539 40103
rect 10241 40069 10275 40103
rect 19257 40069 19291 40103
rect 1409 40001 1443 40035
rect 2235 40011 2269 40045
rect 3341 40001 3375 40035
rect 5147 40001 5181 40035
rect 7757 40001 7791 40035
rect 8217 40001 8251 40035
rect 9873 40001 9907 40035
rect 11069 40001 11103 40035
rect 12725 40001 12759 40035
rect 19993 40001 20027 40035
rect 20269 40001 20303 40035
rect 20537 40001 20571 40035
rect 20821 40001 20855 40035
rect 21097 40001 21131 40035
rect 21373 40001 21407 40035
rect 21649 40001 21683 40035
rect 22017 40001 22051 40035
rect 22293 40001 22327 40035
rect 22569 40001 22603 40035
rect 22845 40001 22879 40035
rect 23121 40001 23155 40035
rect 23397 40001 23431 40035
rect 23857 40001 23891 40035
rect 24133 40001 24167 40035
rect 1961 39933 1995 39967
rect 3525 39933 3559 39967
rect 4445 39933 4479 39967
rect 4905 39933 4939 39967
rect 11805 39933 11839 39967
rect 11989 39933 12023 39967
rect 12842 39933 12876 39967
rect 13001 39933 13035 39967
rect 12449 39865 12483 39899
rect 19441 39865 19475 39899
rect 20637 39865 20671 39899
rect 22661 39865 22695 39899
rect 23213 39865 23247 39899
rect 2973 39797 3007 39831
rect 4077 39797 4111 39831
rect 5917 39797 5951 39831
rect 8769 39797 8803 39831
rect 10425 39797 10459 39831
rect 13645 39797 13679 39831
rect 20361 39797 20395 39831
rect 21465 39797 21499 39831
rect 21833 39797 21867 39831
rect 22109 39797 22143 39831
rect 22385 39797 22419 39831
rect 22937 39797 22971 39831
rect 23673 39797 23707 39831
rect 24409 39797 24443 39831
rect 8401 39593 8435 39627
rect 10517 39593 10551 39627
rect 13369 39593 13403 39627
rect 20729 39593 20763 39627
rect 21557 39593 21591 39627
rect 21833 39593 21867 39627
rect 22385 39593 22419 39627
rect 22845 39593 22879 39627
rect 3249 39525 3283 39559
rect 5273 39525 5307 39559
rect 6101 39525 6135 39559
rect 23213 39525 23247 39559
rect 5457 39457 5491 39491
rect 6494 39457 6528 39491
rect 6653 39457 6687 39491
rect 7389 39457 7423 39491
rect 12357 39457 12391 39491
rect 2237 39389 2271 39423
rect 4353 39389 4387 39423
rect 5641 39389 5675 39423
rect 6377 39389 6411 39423
rect 7663 39389 7697 39423
rect 9505 39389 9539 39423
rect 9779 39389 9813 39423
rect 12599 39389 12633 39423
rect 20913 39389 20947 39423
rect 21281 39389 21315 39423
rect 21741 39389 21775 39423
rect 22017 39389 22051 39423
rect 22293 39389 22327 39423
rect 22569 39389 22603 39423
rect 23029 39389 23063 39423
rect 23397 39389 23431 39423
rect 23857 39389 23891 39423
rect 23949 39389 23983 39423
rect 1501 39321 1535 39355
rect 1685 39321 1719 39355
rect 2329 39321 2363 39355
rect 2697 39321 2731 39355
rect 3065 39321 3099 39355
rect 4261 39321 4295 39355
rect 4721 39321 4755 39355
rect 1961 39253 1995 39287
rect 3985 39253 4019 39287
rect 5089 39253 5123 39287
rect 7297 39253 7331 39287
rect 21097 39253 21131 39287
rect 22109 39253 22143 39287
rect 23673 39253 23707 39287
rect 24133 39253 24167 39287
rect 20453 39049 20487 39083
rect 20729 39049 20763 39083
rect 23397 39049 23431 39083
rect 23673 39049 23707 39083
rect 24133 38981 24167 39015
rect 1959 38913 1993 38947
rect 3065 38913 3099 38947
rect 4077 38913 4111 38947
rect 4629 38913 4663 38947
rect 4905 38913 4939 38947
rect 8399 38913 8433 38947
rect 11771 38913 11805 38947
rect 20637 38897 20671 38931
rect 20913 38913 20947 38947
rect 21649 38913 21683 38947
rect 22089 38913 22123 38947
rect 23581 38913 23615 38947
rect 23857 38913 23891 38947
rect 1685 38845 1719 38879
rect 3801 38845 3835 38879
rect 4353 38845 4387 38879
rect 8125 38845 8159 38879
rect 11529 38845 11563 38879
rect 21833 38845 21867 38879
rect 23213 38777 23247 38811
rect 2697 38709 2731 38743
rect 9137 38709 9171 38743
rect 12541 38709 12575 38743
rect 21465 38709 21499 38743
rect 24409 38709 24443 38743
rect 13277 38505 13311 38539
rect 19901 38505 19935 38539
rect 22477 38505 22511 38539
rect 23305 38505 23339 38539
rect 23673 38505 23707 38539
rect 6009 38437 6043 38471
rect 12081 38437 12115 38471
rect 23029 38437 23063 38471
rect 6402 38369 6436 38403
rect 9137 38369 9171 38403
rect 11621 38369 11655 38403
rect 12474 38369 12508 38403
rect 3801 38301 3835 38335
rect 4059 38271 4093 38305
rect 5365 38301 5399 38335
rect 5549 38301 5583 38335
rect 6285 38301 6319 38335
rect 6561 38301 6595 38335
rect 9411 38301 9445 38335
rect 11437 38301 11471 38335
rect 12357 38301 12391 38335
rect 12633 38301 12667 38335
rect 20085 38301 20119 38335
rect 22109 38301 22143 38335
rect 22661 38301 22695 38335
rect 22753 38301 22787 38335
rect 22937 38301 22971 38335
rect 23213 38301 23247 38335
rect 23489 38301 23523 38335
rect 23857 38301 23891 38335
rect 23949 38301 23983 38335
rect 1409 38233 1443 38267
rect 2237 38233 2271 38267
rect 2421 38233 2455 38267
rect 3157 38233 3191 38267
rect 4813 38165 4847 38199
rect 7205 38165 7239 38199
rect 10149 38165 10183 38199
rect 22201 38165 22235 38199
rect 22937 38165 22971 38199
rect 24133 38165 24167 38199
rect 7389 37961 7423 37995
rect 8953 37961 8987 37995
rect 13093 37961 13127 37995
rect 21465 37961 21499 37995
rect 23857 37961 23891 37995
rect 1685 37893 1719 37927
rect 3525 37893 3559 37927
rect 3893 37893 3927 37927
rect 4629 37893 4663 37927
rect 5825 37893 5859 37927
rect 9229 37893 9263 37927
rect 9321 37893 9355 37927
rect 23765 37893 23799 37927
rect 1409 37825 1443 37859
rect 2203 37825 2237 37859
rect 3801 37825 3835 37859
rect 4261 37825 4295 37859
rect 4997 37825 5031 37859
rect 5549 37825 5583 37859
rect 6651 37825 6685 37859
rect 9689 37825 9723 37859
rect 10071 37825 10105 37859
rect 12081 37825 12115 37859
rect 12355 37825 12389 37859
rect 21649 37825 21683 37859
rect 22107 37825 22141 37859
rect 23397 37825 23431 37859
rect 24041 37825 24075 37859
rect 24225 37825 24259 37859
rect 1961 37757 1995 37791
rect 5273 37757 5307 37791
rect 6377 37757 6411 37791
rect 21833 37757 21867 37791
rect 23213 37757 23247 37791
rect 2973 37689 3007 37723
rect 22845 37689 22879 37723
rect 23673 37689 23707 37723
rect 4813 37621 4847 37655
rect 10241 37621 10275 37655
rect 24409 37621 24443 37655
rect 21649 37417 21683 37451
rect 21925 37417 21959 37451
rect 22569 37417 22603 37451
rect 22845 37417 22879 37451
rect 8217 37281 8251 37315
rect 8401 37281 8435 37315
rect 24133 37281 24167 37315
rect 2513 37213 2547 37247
rect 3801 37213 3835 37247
rect 4721 37213 4755 37247
rect 4995 37213 5029 37247
rect 6561 37213 6595 37247
rect 6819 37183 6853 37217
rect 7941 37213 7975 37247
rect 8033 37213 8067 37247
rect 8309 37213 8343 37247
rect 8493 37213 8527 37247
rect 10057 37213 10091 37247
rect 10315 37183 10349 37217
rect 20729 37213 20763 37247
rect 21833 37213 21867 37247
rect 22109 37213 22143 37247
rect 22753 37213 22787 37247
rect 23029 37213 23063 37247
rect 23305 37213 23339 37247
rect 23581 37213 23615 37247
rect 1409 37145 1443 37179
rect 2237 37145 2271 37179
rect 2789 37145 2823 37179
rect 3157 37145 3191 37179
rect 4077 37145 4111 37179
rect 23857 37145 23891 37179
rect 3433 37077 3467 37111
rect 5733 37077 5767 37111
rect 7573 37077 7607 37111
rect 8217 37077 8251 37111
rect 11069 37077 11103 37111
rect 20545 37077 20579 37111
rect 23121 37077 23155 37111
rect 23397 37077 23431 37111
rect 5917 36873 5951 36907
rect 7021 36873 7055 36907
rect 19625 36873 19659 36907
rect 20361 36873 20395 36907
rect 20913 36873 20947 36907
rect 23949 36873 23983 36907
rect 1593 36805 1627 36839
rect 3433 36805 3467 36839
rect 3709 36805 3743 36839
rect 3801 36805 3835 36839
rect 23673 36805 23707 36839
rect 2143 36737 2177 36771
rect 4169 36737 4203 36771
rect 4551 36737 4585 36771
rect 5179 36737 5213 36771
rect 6929 36737 6963 36771
rect 7389 36737 7423 36771
rect 7755 36737 7789 36771
rect 11771 36737 11805 36771
rect 17785 36737 17819 36771
rect 19165 36737 19199 36771
rect 19809 36741 19843 36775
rect 20269 36737 20303 36771
rect 20545 36737 20579 36771
rect 20821 36737 20855 36771
rect 21097 36737 21131 36771
rect 23029 36737 23063 36771
rect 23305 36737 23339 36771
rect 24133 36737 24167 36771
rect 24225 36737 24259 36771
rect 1869 36669 1903 36703
rect 4905 36669 4939 36703
rect 7481 36669 7515 36703
rect 11529 36669 11563 36703
rect 1777 36601 1811 36635
rect 2881 36601 2915 36635
rect 18981 36601 19015 36635
rect 20085 36601 20119 36635
rect 23121 36601 23155 36635
rect 4721 36533 4755 36567
rect 7205 36533 7239 36567
rect 8493 36533 8527 36567
rect 12541 36533 12575 36567
rect 17601 36533 17635 36567
rect 20637 36533 20671 36567
rect 22845 36533 22879 36567
rect 24409 36533 24443 36567
rect 4721 36329 4755 36363
rect 7021 36329 7055 36363
rect 22385 36329 22419 36363
rect 23397 36329 23431 36363
rect 5733 36261 5767 36295
rect 10977 36261 11011 36295
rect 6147 36193 6181 36227
rect 6285 36193 6319 36227
rect 8953 36193 8987 36227
rect 11529 36193 11563 36227
rect 1501 36125 1535 36159
rect 1775 36125 1809 36159
rect 2881 36125 2915 36159
rect 3801 36125 3835 36159
rect 5089 36125 5123 36159
rect 5273 36125 5307 36159
rect 6009 36125 6043 36159
rect 6929 36125 6963 36159
rect 7205 36125 7239 36159
rect 9195 36125 9229 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 11253 36125 11287 36159
rect 11391 36125 11425 36159
rect 17141 36125 17175 36159
rect 18797 36125 18831 36159
rect 21189 36125 21223 36159
rect 21833 36125 21867 36159
rect 22569 36125 22603 36159
rect 23581 36125 23615 36159
rect 23857 36125 23891 36159
rect 3157 36057 3191 36091
rect 4077 36057 4111 36091
rect 4445 36057 4479 36091
rect 12173 36057 12207 36091
rect 17386 36057 17420 36091
rect 24225 36057 24259 36091
rect 2513 35989 2547 36023
rect 9965 35989 9999 36023
rect 18521 35989 18555 36023
rect 18613 35989 18647 36023
rect 21005 35989 21039 36023
rect 21649 35989 21683 36023
rect 3341 35785 3375 35819
rect 6193 35785 6227 35819
rect 11713 35785 11747 35819
rect 14197 35785 14231 35819
rect 21833 35785 21867 35819
rect 23121 35785 23155 35819
rect 23489 35785 23523 35819
rect 8217 35717 8251 35751
rect 8585 35717 8619 35751
rect 9321 35717 9355 35751
rect 11989 35717 12023 35751
rect 12081 35717 12115 35751
rect 12817 35717 12851 35751
rect 19257 35717 19291 35751
rect 1685 35649 1719 35683
rect 2697 35649 2731 35683
rect 3433 35649 3467 35683
rect 4537 35649 4571 35683
rect 8493 35649 8527 35683
rect 8953 35649 8987 35683
rect 9963 35649 9997 35683
rect 12449 35649 12483 35683
rect 13459 35649 13493 35683
rect 17843 35649 17877 35683
rect 18981 35649 19015 35683
rect 19349 35649 19383 35683
rect 19533 35649 19567 35683
rect 21281 35649 21315 35683
rect 22017 35649 22051 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 23305 35649 23339 35683
rect 23673 35649 23707 35683
rect 23949 35649 23983 35683
rect 24133 35649 24167 35683
rect 1501 35581 1535 35615
rect 2421 35581 2455 35615
rect 2538 35581 2572 35615
rect 3617 35581 3651 35615
rect 4353 35581 4387 35615
rect 5273 35581 5307 35615
rect 5390 35581 5424 35615
rect 5549 35581 5583 35615
rect 9689 35581 9723 35615
rect 13185 35581 13219 35615
rect 17601 35581 17635 35615
rect 19073 35581 19107 35615
rect 19257 35581 19291 35615
rect 19441 35581 19475 35615
rect 2145 35513 2179 35547
rect 4997 35513 5031 35547
rect 9505 35513 9539 35547
rect 18613 35513 18647 35547
rect 21097 35513 21131 35547
rect 22661 35513 22695 35547
rect 7757 35445 7791 35479
rect 10701 35445 10735 35479
rect 13001 35445 13035 35479
rect 22385 35445 22419 35479
rect 23765 35445 23799 35479
rect 24409 35445 24443 35479
rect 6469 35241 6503 35275
rect 12817 35241 12851 35275
rect 18245 35241 18279 35275
rect 23213 35241 23247 35275
rect 3341 35173 3375 35207
rect 10517 35173 10551 35207
rect 19901 35173 19935 35207
rect 2329 35105 2363 35139
rect 10057 35105 10091 35139
rect 10793 35105 10827 35139
rect 11805 35105 11839 35139
rect 15669 35105 15703 35139
rect 1409 35037 1443 35071
rect 2571 35037 2605 35071
rect 4261 35037 4295 35071
rect 5457 35037 5491 35071
rect 5731 35037 5765 35071
rect 9873 35037 9907 35071
rect 10931 35037 10965 35071
rect 11069 35037 11103 35071
rect 12079 35037 12113 35071
rect 14105 35037 14139 35071
rect 14379 35037 14413 35071
rect 15943 35037 15977 35071
rect 18153 35037 18187 35071
rect 19717 35037 19751 35071
rect 20085 35013 20119 35047
rect 21005 35037 21039 35071
rect 23397 35037 23431 35071
rect 23673 35037 23707 35071
rect 23949 35037 23983 35071
rect 1685 34969 1719 35003
rect 4353 34969 4387 35003
rect 4721 34969 4755 35003
rect 11713 34969 11747 35003
rect 3985 34901 4019 34935
rect 5089 34901 5123 34935
rect 5273 34901 5307 34935
rect 15117 34901 15151 34935
rect 16681 34901 16715 34935
rect 19533 34901 19567 34935
rect 20821 34901 20855 34935
rect 23489 34901 23523 34935
rect 24133 34901 24167 34935
rect 2421 34697 2455 34731
rect 4537 34697 4571 34731
rect 9045 34697 9079 34731
rect 11069 34697 11103 34731
rect 15209 34697 15243 34731
rect 16957 34697 16991 34731
rect 18797 34697 18831 34731
rect 21465 34697 21499 34731
rect 23673 34697 23707 34731
rect 3065 34629 3099 34663
rect 24133 34629 24167 34663
rect 1683 34561 1717 34595
rect 2789 34561 2823 34595
rect 3799 34561 3833 34595
rect 4905 34561 4939 34595
rect 5181 34561 5215 34595
rect 6651 34561 6685 34595
rect 8769 34561 8803 34595
rect 9321 34561 9355 34595
rect 9505 34561 9539 34595
rect 9597 34561 9631 34595
rect 10299 34561 10333 34595
rect 14471 34561 14505 34595
rect 16681 34561 16715 34595
rect 17049 34561 17083 34595
rect 17325 34561 17359 34595
rect 17509 34561 17543 34595
rect 18981 34561 19015 34595
rect 19073 34561 19107 34595
rect 19340 34561 19374 34595
rect 20545 34561 20579 34595
rect 21005 34561 21039 34595
rect 21649 34561 21683 34595
rect 22091 34591 22125 34625
rect 23397 34561 23431 34595
rect 23857 34561 23891 34595
rect 1409 34493 1443 34527
rect 3525 34493 3559 34527
rect 6377 34493 6411 34527
rect 9045 34493 9079 34527
rect 10057 34493 10091 34527
rect 14197 34493 14231 34527
rect 16957 34493 16991 34527
rect 17417 34493 17451 34527
rect 20637 34493 20671 34527
rect 21833 34493 21867 34527
rect 24409 34493 24443 34527
rect 16773 34425 16807 34459
rect 17141 34425 17175 34459
rect 23213 34425 23247 34459
rect 7389 34357 7423 34391
rect 8861 34357 8895 34391
rect 9413 34357 9447 34391
rect 9689 34357 9723 34391
rect 20453 34357 20487 34391
rect 20821 34357 20855 34391
rect 22845 34357 22879 34391
rect 9965 34153 9999 34187
rect 17325 34153 17359 34187
rect 21097 34153 21131 34187
rect 22385 34153 22419 34187
rect 7481 34085 7515 34119
rect 13553 34085 13587 34119
rect 20637 34085 20671 34119
rect 23121 34085 23155 34119
rect 3065 34017 3099 34051
rect 4537 34017 4571 34051
rect 7895 34017 7929 34051
rect 15945 34017 15979 34051
rect 19625 34017 19659 34051
rect 21281 34017 21315 34051
rect 21465 34017 21499 34051
rect 1409 33949 1443 33983
rect 1683 33949 1717 33983
rect 2789 33949 2823 33983
rect 3801 33949 3835 33983
rect 4779 33949 4813 33983
rect 6837 33949 6871 33983
rect 7021 33949 7055 33983
rect 7757 33949 7791 33983
rect 8033 33949 8067 33983
rect 8953 33949 8987 33983
rect 9195 33949 9229 33983
rect 12541 33949 12575 33983
rect 12815 33949 12849 33983
rect 14105 33949 14139 33983
rect 14347 33949 14381 33983
rect 16187 33949 16221 33983
rect 17509 33949 17543 33983
rect 17877 33949 17911 33983
rect 18153 33949 18187 33983
rect 19899 33949 19933 33983
rect 21005 33949 21039 33983
rect 21373 33949 21407 33983
rect 21557 33949 21591 33983
rect 22569 33949 22603 33983
rect 22845 33949 22879 33983
rect 23305 33949 23339 33983
rect 23581 33949 23615 33983
rect 23857 33949 23891 33983
rect 23949 33949 23983 33983
rect 4077 33881 4111 33915
rect 2421 33813 2455 33847
rect 5549 33813 5583 33847
rect 8677 33813 8711 33847
rect 15117 33813 15151 33847
rect 16957 33813 16991 33847
rect 17693 33813 17727 33847
rect 18245 33813 18279 33847
rect 21281 33813 21315 33847
rect 22661 33813 22695 33847
rect 23397 33813 23431 33847
rect 23673 33813 23707 33847
rect 24133 33813 24167 33847
rect 3065 33609 3099 33643
rect 4353 33609 4387 33643
rect 8861 33609 8895 33643
rect 9137 33609 9171 33643
rect 16957 33609 16991 33643
rect 23213 33609 23247 33643
rect 3341 33541 3375 33575
rect 4169 33541 4203 33575
rect 13645 33541 13679 33575
rect 24133 33541 24167 33575
rect 1743 33473 1777 33507
rect 3433 33473 3467 33507
rect 3801 33473 3835 33507
rect 5147 33473 5181 33507
rect 8125 33473 8159 33507
rect 9045 33473 9079 33507
rect 9321 33473 9355 33507
rect 9779 33473 9813 33507
rect 11805 33473 11839 33507
rect 11989 33473 12023 33507
rect 15451 33473 15485 33507
rect 17141 33473 17175 33507
rect 17233 33473 17267 33507
rect 17489 33473 17523 33507
rect 18705 33473 18739 33507
rect 19073 33473 19107 33507
rect 19257 33473 19291 33507
rect 19533 33473 19567 33507
rect 21649 33473 21683 33507
rect 21833 33473 21867 33507
rect 22089 33473 22123 33507
rect 23305 33473 23339 33507
rect 23673 33473 23707 33507
rect 23857 33473 23891 33507
rect 1501 33405 1535 33439
rect 4905 33405 4939 33439
rect 6929 33405 6963 33439
rect 7113 33405 7147 33439
rect 7849 33405 7883 33439
rect 7987 33405 8021 33439
rect 8769 33405 8803 33439
rect 9505 33405 9539 33439
rect 12725 33405 12759 33439
rect 12842 33405 12876 33439
rect 13001 33405 13035 33439
rect 15209 33405 15243 33439
rect 18797 33405 18831 33439
rect 18981 33405 19015 33439
rect 19165 33405 19199 33439
rect 23581 33405 23615 33439
rect 23765 33405 23799 33439
rect 2513 33337 2547 33371
rect 7573 33337 7607 33371
rect 12449 33337 12483 33371
rect 18613 33337 18647 33371
rect 19349 33337 19383 33371
rect 5917 33269 5951 33303
rect 10517 33269 10551 33303
rect 16221 33269 16255 33303
rect 18889 33269 18923 33303
rect 21465 33269 21499 33303
rect 23397 33269 23431 33303
rect 23489 33269 23523 33303
rect 24409 33269 24443 33303
rect 3341 33065 3375 33099
rect 4537 33065 4571 33099
rect 8217 33065 8251 33099
rect 12909 33065 12943 33099
rect 15945 33065 15979 33099
rect 18613 33065 18647 33099
rect 22293 33065 22327 33099
rect 10609 32997 10643 33031
rect 14749 32997 14783 33031
rect 21925 32997 21959 33031
rect 23673 32997 23707 33031
rect 2329 32929 2363 32963
rect 3985 32929 4019 32963
rect 7205 32929 7239 32963
rect 10149 32929 10183 32963
rect 11023 32929 11057 32963
rect 11897 32929 11931 32963
rect 15163 32929 15197 32963
rect 17601 32929 17635 32963
rect 1409 32861 1443 32895
rect 2603 32861 2637 32895
rect 3801 32861 3835 32895
rect 5273 32861 5307 32895
rect 5365 32861 5399 32895
rect 7463 32831 7497 32865
rect 9965 32861 9999 32895
rect 10885 32861 10919 32895
rect 11161 32861 11195 32895
rect 12139 32861 12173 32895
rect 14105 32861 14139 32895
rect 14289 32861 14323 32895
rect 15025 32861 15059 32895
rect 15301 32861 15335 32895
rect 17843 32861 17877 32895
rect 22101 32861 22135 32895
rect 22201 32863 22235 32897
rect 23029 32861 23063 32895
rect 23581 32861 23615 32895
rect 23857 32861 23891 32895
rect 23949 32861 23983 32895
rect 1685 32793 1719 32827
rect 5733 32793 5767 32827
rect 11805 32793 11839 32827
rect 4997 32725 5031 32759
rect 6101 32725 6135 32759
rect 6285 32725 6319 32759
rect 22845 32725 22879 32759
rect 23397 32725 23431 32759
rect 24133 32725 24167 32759
rect 11069 32521 11103 32555
rect 14105 32521 14139 32555
rect 15209 32521 15243 32555
rect 15393 32521 15427 32555
rect 22661 32521 22695 32555
rect 23673 32521 23707 32555
rect 3893 32453 3927 32487
rect 14340 32453 14374 32487
rect 14473 32453 14507 32487
rect 19432 32453 19466 32487
rect 2446 32385 2480 32419
rect 3341 32385 3375 32419
rect 8307 32385 8341 32419
rect 10057 32385 10091 32419
rect 10315 32415 10349 32449
rect 14841 32385 14875 32419
rect 19165 32385 19199 32419
rect 22017 32385 22051 32419
rect 22569 32385 22603 32419
rect 22845 32385 22879 32419
rect 23305 32385 23339 32419
rect 23581 32385 23615 32419
rect 23857 32385 23891 32419
rect 24133 32385 24167 32419
rect 24225 32385 24259 32419
rect 1409 32317 1443 32351
rect 1593 32317 1627 32351
rect 2053 32317 2087 32351
rect 2329 32317 2363 32351
rect 2605 32317 2639 32351
rect 3249 32317 3283 32351
rect 3617 32317 3651 32351
rect 4629 32317 4663 32351
rect 8033 32317 8067 32351
rect 21833 32249 21867 32283
rect 23397 32249 23431 32283
rect 9045 32181 9079 32215
rect 20545 32181 20579 32215
rect 22385 32181 22419 32215
rect 23121 32181 23155 32215
rect 23949 32181 23983 32215
rect 24409 32181 24443 32215
rect 2421 31977 2455 32011
rect 4721 31977 4755 32011
rect 15117 31977 15151 32011
rect 17417 31977 17451 32011
rect 23489 31977 23523 32011
rect 16221 31909 16255 31943
rect 19533 31909 19567 31943
rect 20637 31909 20671 31943
rect 20913 31909 20947 31943
rect 21189 31909 21223 31943
rect 21649 31909 21683 31943
rect 3065 31841 3099 31875
rect 14105 31841 14139 31875
rect 15761 31841 15795 31875
rect 16497 31841 16531 31875
rect 16614 31841 16648 31875
rect 16773 31841 16807 31875
rect 1409 31773 1443 31807
rect 1683 31773 1717 31807
rect 2789 31773 2823 31807
rect 3801 31773 3835 31807
rect 4905 31773 4939 31807
rect 5825 31773 5859 31807
rect 6099 31773 6133 31807
rect 11069 31773 11103 31807
rect 11343 31773 11377 31807
rect 13093 31773 13127 31807
rect 14379 31773 14413 31807
rect 15577 31773 15611 31807
rect 19717 31773 19751 31807
rect 20085 31773 20119 31807
rect 20177 31773 20211 31807
rect 20821 31773 20855 31807
rect 21097 31773 21131 31807
rect 21373 31773 21407 31807
rect 21833 31773 21867 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24225 31773 24259 31807
rect 4077 31705 4111 31739
rect 6837 31637 6871 31671
rect 12081 31637 12115 31671
rect 13185 31637 13219 31671
rect 3893 31433 3927 31467
rect 8677 31433 8711 31467
rect 4169 31365 4203 31399
rect 4445 31365 4479 31399
rect 4537 31365 4571 31399
rect 5273 31365 5307 31399
rect 6561 31365 6595 31399
rect 6837 31365 6871 31399
rect 6929 31365 6963 31399
rect 7665 31365 7699 31399
rect 8953 31365 8987 31399
rect 9045 31365 9079 31399
rect 9781 31365 9815 31399
rect 12265 31365 12299 31399
rect 1683 31307 1717 31341
rect 3065 31297 3099 31331
rect 3709 31297 3743 31331
rect 4905 31297 4939 31331
rect 7297 31297 7331 31331
rect 9413 31297 9447 31331
rect 11621 31297 11655 31331
rect 12783 31297 12817 31331
rect 13921 31297 13955 31331
rect 14105 31297 14139 31331
rect 15375 31327 15409 31361
rect 16681 31297 16715 31331
rect 16955 31297 16989 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 19807 31297 19841 31331
rect 21097 31297 21131 31331
rect 21465 31297 21499 31331
rect 22477 31297 22511 31331
rect 23121 31297 23155 31331
rect 23765 31297 23799 31331
rect 24133 31297 24167 31331
rect 24225 31297 24259 31331
rect 1409 31229 1443 31263
rect 2789 31229 2823 31263
rect 12541 31229 12575 31263
rect 15117 31229 15151 31263
rect 19533 31229 19567 31263
rect 20913 31229 20947 31263
rect 5457 31161 5491 31195
rect 7849 31161 7883 31195
rect 9965 31161 9999 31195
rect 12449 31161 12483 31195
rect 13553 31161 13587 31195
rect 18061 31161 18095 31195
rect 20545 31161 20579 31195
rect 22293 31161 22327 31195
rect 22937 31161 22971 31195
rect 23581 31161 23615 31195
rect 2421 31093 2455 31127
rect 11713 31093 11747 31127
rect 14013 31093 14047 31127
rect 16129 31093 16163 31127
rect 17693 31093 17727 31127
rect 18613 31093 18647 31127
rect 21373 31093 21407 31127
rect 23949 31093 23983 31127
rect 24409 31093 24443 31127
rect 3341 30889 3375 30923
rect 5273 30889 5307 30923
rect 7389 30889 7423 30923
rect 9965 30889 9999 30923
rect 12541 30889 12575 30923
rect 12817 30889 12851 30923
rect 17601 30889 17635 30923
rect 19349 30889 19383 30923
rect 20729 30889 20763 30923
rect 23121 30889 23155 30923
rect 16405 30821 16439 30855
rect 19073 30821 19107 30855
rect 19901 30821 19935 30855
rect 22845 30821 22879 30855
rect 23489 30821 23523 30855
rect 6377 30753 6411 30787
rect 8953 30753 8987 30787
rect 10517 30753 10551 30787
rect 11161 30753 11195 30787
rect 11437 30753 11471 30787
rect 11554 30753 11588 30787
rect 11713 30753 11747 30787
rect 15117 30753 15151 30787
rect 16798 30753 16832 30787
rect 16957 30753 16991 30787
rect 17693 30753 17727 30787
rect 19533 30753 19567 30787
rect 19717 30753 19751 30787
rect 2329 30685 2363 30719
rect 2603 30685 2637 30719
rect 3801 30685 3835 30719
rect 4261 30685 4295 30719
rect 4535 30685 4569 30719
rect 6651 30685 6685 30719
rect 9227 30685 9261 30719
rect 10701 30685 10735 30719
rect 12357 30685 12391 30719
rect 12725 30685 12759 30719
rect 13001 30685 13035 30719
rect 14105 30685 14139 30719
rect 14473 30685 14507 30719
rect 14933 30685 14967 30719
rect 15761 30685 15795 30719
rect 15945 30685 15979 30719
rect 16681 30685 16715 30719
rect 17949 30685 17983 30719
rect 19257 30685 19291 30719
rect 19625 30685 19659 30719
rect 19809 30685 19843 30719
rect 20085 30685 20119 30719
rect 20637 30685 20671 30719
rect 20821 30685 20855 30719
rect 22293 30685 22327 30719
rect 23029 30685 23063 30719
rect 23305 30685 23339 30719
rect 23673 30685 23707 30719
rect 1501 30617 1535 30651
rect 1685 30617 1719 30651
rect 19533 30617 19567 30651
rect 23857 30617 23891 30651
rect 24225 30617 24259 30651
rect 3985 30549 4019 30583
rect 22109 30549 22143 30583
rect 3893 30345 3927 30379
rect 10977 30345 11011 30379
rect 23765 30345 23799 30379
rect 3341 30277 3375 30311
rect 24133 30277 24167 30311
rect 2421 30209 2455 30243
rect 2697 30209 2731 30243
rect 3433 30209 3467 30243
rect 3709 30209 3743 30243
rect 4443 30209 4477 30243
rect 7111 30209 7145 30243
rect 9965 30209 9999 30243
rect 10239 30209 10273 30243
rect 13921 30209 13955 30243
rect 14195 30209 14229 30243
rect 17969 30209 18003 30243
rect 18227 30239 18261 30273
rect 20525 30209 20559 30243
rect 22107 30209 22141 30243
rect 23397 30209 23431 30243
rect 23673 30209 23707 30243
rect 23949 30209 23983 30243
rect 1501 30141 1535 30175
rect 1685 30141 1719 30175
rect 2145 30141 2179 30175
rect 2559 30141 2593 30175
rect 4169 30141 4203 30175
rect 6837 30141 6871 30175
rect 20269 30141 20303 30175
rect 21833 30141 21867 30175
rect 18981 30073 19015 30107
rect 23489 30073 23523 30107
rect 3617 30005 3651 30039
rect 5181 30005 5215 30039
rect 7849 30005 7883 30039
rect 14933 30005 14967 30039
rect 21649 30005 21683 30039
rect 22845 30005 22879 30039
rect 23213 30005 23247 30039
rect 24409 30005 24443 30039
rect 2697 29801 2731 29835
rect 3249 29801 3283 29835
rect 3617 29801 3651 29835
rect 8769 29801 8803 29835
rect 12357 29801 12391 29835
rect 17417 29801 17451 29835
rect 7573 29733 7607 29767
rect 11161 29733 11195 29767
rect 13461 29733 13495 29767
rect 16221 29733 16255 29767
rect 23305 29733 23339 29767
rect 23581 29733 23615 29767
rect 4077 29665 4111 29699
rect 7849 29665 7883 29699
rect 7987 29665 8021 29699
rect 10701 29665 10735 29699
rect 11437 29665 11471 29699
rect 11575 29665 11609 29699
rect 11713 29665 11747 29699
rect 14197 29665 14231 29699
rect 15761 29665 15795 29699
rect 16497 29665 16531 29699
rect 16773 29665 16807 29699
rect 21741 29665 21775 29699
rect 22109 29665 22143 29699
rect 22293 29665 22327 29699
rect 22477 29665 22511 29699
rect 1685 29597 1719 29631
rect 1959 29597 1993 29631
rect 3433 29597 3467 29631
rect 3801 29597 3835 29631
rect 5273 29597 5307 29631
rect 6929 29597 6963 29631
rect 7113 29597 7147 29631
rect 8125 29597 8159 29631
rect 10517 29597 10551 29631
rect 12449 29597 12483 29631
rect 12723 29597 12757 29631
rect 14439 29597 14473 29631
rect 15577 29597 15611 29631
rect 16614 29597 16648 29631
rect 21189 29597 21223 29631
rect 21649 29597 21683 29631
rect 22017 29597 22051 29631
rect 22385 29597 22419 29631
rect 22569 29597 22603 29631
rect 23489 29597 23523 29631
rect 23765 29597 23799 29631
rect 23949 29597 23983 29631
rect 3157 29529 3191 29563
rect 5365 29529 5399 29563
rect 5733 29529 5767 29563
rect 22293 29529 22327 29563
rect 4997 29461 5031 29495
rect 6101 29461 6135 29495
rect 6285 29461 6319 29495
rect 15209 29461 15243 29495
rect 21005 29461 21039 29495
rect 24133 29461 24167 29495
rect 5917 29257 5951 29291
rect 8401 29257 8435 29291
rect 10885 29257 10919 29291
rect 11713 29257 11747 29291
rect 14289 29257 14323 29291
rect 23121 29257 23155 29291
rect 1869 29189 1903 29223
rect 2053 29189 2087 29223
rect 11621 29189 11655 29223
rect 14657 29189 14691 29223
rect 15393 29189 15427 29223
rect 1501 29121 1535 29155
rect 2479 29121 2513 29155
rect 3617 29121 3651 29155
rect 5179 29121 5213 29155
rect 7389 29121 7423 29155
rect 7663 29121 7697 29155
rect 9229 29121 9263 29155
rect 9471 29131 9505 29165
rect 10609 29121 10643 29155
rect 12815 29121 12849 29155
rect 14565 29121 14599 29155
rect 15025 29121 15059 29155
rect 16955 29121 16989 29155
rect 18889 29121 18923 29155
rect 19147 29151 19181 29185
rect 20269 29121 20303 29155
rect 20453 29121 20487 29155
rect 23305 29121 23339 29155
rect 23581 29121 23615 29155
rect 23857 29121 23891 29155
rect 24133 29121 24167 29155
rect 1685 29053 1719 29087
rect 2237 29053 2271 29087
rect 4905 29053 4939 29087
rect 10885 29053 10919 29087
rect 12541 29053 12575 29087
rect 16681 29053 16715 29087
rect 3249 28985 3283 29019
rect 3801 28985 3835 29019
rect 10241 28985 10275 29019
rect 10701 28985 10735 29019
rect 15577 28985 15611 29019
rect 23397 28985 23431 29019
rect 23673 28985 23707 29019
rect 13553 28917 13587 28951
rect 17693 28917 17727 28951
rect 19901 28917 19935 28951
rect 20361 28917 20395 28951
rect 24409 28917 24443 28951
rect 2237 28713 2271 28747
rect 11161 28713 11195 28747
rect 11437 28713 11471 28747
rect 18889 28713 18923 28747
rect 23489 28713 23523 28747
rect 10517 28645 10551 28679
rect 10793 28645 10827 28679
rect 18429 28645 18463 28679
rect 23213 28645 23247 28679
rect 2329 28577 2363 28611
rect 16681 28577 16715 28611
rect 16957 28577 16991 28611
rect 17233 28577 17267 28611
rect 19349 28577 19383 28611
rect 19717 28577 19751 28611
rect 19901 28577 19935 28611
rect 1777 28509 1811 28543
rect 2053 28509 2087 28543
rect 2603 28509 2637 28543
rect 3893 28509 3927 28543
rect 4167 28509 4201 28543
rect 8953 28509 8987 28543
rect 9227 28509 9261 28543
rect 10701 28509 10735 28543
rect 10977 28509 11011 28543
rect 11069 28509 11103 28543
rect 11345 28509 11379 28543
rect 11529 28509 11563 28543
rect 11713 28509 11747 28543
rect 11987 28509 12021 28543
rect 14105 28509 14139 28543
rect 14379 28509 14413 28543
rect 16037 28509 16071 28543
rect 16221 28509 16255 28543
rect 17074 28509 17108 28543
rect 17877 28509 17911 28543
rect 18613 28509 18647 28543
rect 19073 28509 19107 28543
rect 19257 28509 19291 28543
rect 19625 28509 19659 28543
rect 19993 28509 20027 28543
rect 20267 28509 20301 28543
rect 22845 28509 22879 28543
rect 23397 28509 23431 28543
rect 23673 28509 23707 28543
rect 23949 28509 23983 28543
rect 1501 28441 1535 28475
rect 1593 28373 1627 28407
rect 1961 28373 1995 28407
rect 3341 28373 3375 28407
rect 4905 28373 4939 28407
rect 9965 28373 9999 28407
rect 12725 28373 12759 28407
rect 15117 28373 15151 28407
rect 19901 28373 19935 28407
rect 21005 28373 21039 28407
rect 22661 28373 22695 28407
rect 24133 28373 24167 28407
rect 1593 28169 1627 28203
rect 2513 28169 2547 28203
rect 4077 28169 4111 28203
rect 5825 28169 5859 28203
rect 16221 28169 16255 28203
rect 23489 28169 23523 28203
rect 2789 28101 2823 28135
rect 3157 28101 3191 28135
rect 3893 28101 3927 28135
rect 4537 28101 4571 28135
rect 5273 28101 5307 28135
rect 5641 28101 5675 28135
rect 19708 28101 19742 28135
rect 1501 28033 1535 28067
rect 2329 28033 2363 28067
rect 3065 28033 3099 28067
rect 3525 28033 3559 28067
rect 4813 28033 4847 28067
rect 4905 28033 4939 28067
rect 6651 28033 6685 28067
rect 10331 28043 10365 28077
rect 14013 28033 14047 28067
rect 15451 28033 15485 28067
rect 17877 28033 17911 28067
rect 18133 28033 18167 28067
rect 20913 28033 20947 28067
rect 21281 28033 21315 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22293 28033 22327 28067
rect 22845 28033 22879 28067
rect 23121 28033 23155 28067
rect 23397 28033 23431 28067
rect 23673 28033 23707 28067
rect 23949 28033 23983 28067
rect 24133 28033 24167 28067
rect 6377 27965 6411 27999
rect 10057 27965 10091 27999
rect 12817 27965 12851 27999
rect 13001 27965 13035 27999
rect 13737 27965 13771 27999
rect 13854 27965 13888 27999
rect 15209 27965 15243 27999
rect 19441 27965 19475 27999
rect 21189 27965 21223 27999
rect 21925 27965 21959 27999
rect 13461 27897 13495 27931
rect 19257 27897 19291 27931
rect 21005 27897 21039 27931
rect 21373 27897 21407 27931
rect 22937 27897 22971 27931
rect 23213 27897 23247 27931
rect 7389 27829 7423 27863
rect 11069 27829 11103 27863
rect 14657 27829 14691 27863
rect 20821 27829 20855 27863
rect 21097 27829 21131 27863
rect 22109 27829 22143 27863
rect 22661 27829 22695 27863
rect 23765 27829 23799 27863
rect 24409 27829 24443 27863
rect 22569 27625 22603 27659
rect 23581 27625 23615 27659
rect 5825 27557 5859 27591
rect 10425 27557 10459 27591
rect 19993 27557 20027 27591
rect 20913 27557 20947 27591
rect 22753 27557 22787 27591
rect 23121 27557 23155 27591
rect 1409 27489 1443 27523
rect 22937 27489 22971 27523
rect 23397 27489 23431 27523
rect 1683 27421 1717 27455
rect 2789 27421 2823 27455
rect 4813 27421 4847 27455
rect 5087 27421 5121 27455
rect 7113 27421 7147 27455
rect 9505 27421 9539 27455
rect 11529 27421 11563 27455
rect 11787 27391 11821 27425
rect 15209 27421 15243 27455
rect 16221 27421 16255 27455
rect 16479 27421 16513 27455
rect 17601 27421 17635 27455
rect 17843 27421 17877 27455
rect 20177 27421 20211 27455
rect 21097 27421 21131 27455
rect 21189 27421 21223 27455
rect 22661 27421 22695 27455
rect 23029 27421 23063 27455
rect 23305 27421 23339 27455
rect 23489 27421 23523 27455
rect 23765 27421 23799 27455
rect 23949 27421 23983 27455
rect 6653 27353 6687 27387
rect 6745 27353 6779 27387
rect 9413 27353 9447 27387
rect 9873 27353 9907 27387
rect 10241 27353 10275 27387
rect 21434 27353 21468 27387
rect 2421 27285 2455 27319
rect 2973 27285 3007 27319
rect 6377 27285 6411 27319
rect 7481 27285 7515 27319
rect 7665 27285 7699 27319
rect 9137 27285 9171 27319
rect 12541 27285 12575 27319
rect 15025 27285 15059 27319
rect 17233 27285 17267 27319
rect 18613 27285 18647 27319
rect 22937 27285 22971 27319
rect 24133 27285 24167 27319
rect 2053 27081 2087 27115
rect 3157 27081 3191 27115
rect 3341 27081 3375 27115
rect 3709 27081 3743 27115
rect 5549 27081 5583 27115
rect 8769 27081 8803 27115
rect 14657 27081 14691 27115
rect 22845 27081 22879 27115
rect 23305 27081 23339 27115
rect 23949 27081 23983 27115
rect 2329 26945 2363 26979
rect 2421 26945 2455 26979
rect 2789 26945 2823 26979
rect 3525 26945 3559 26979
rect 4795 26975 4829 27009
rect 8031 26945 8065 26979
rect 12817 26945 12851 26979
rect 13854 26945 13888 26979
rect 14749 26945 14783 26979
rect 15023 26945 15057 26979
rect 16865 26945 16899 26979
rect 17877 26945 17911 26979
rect 21833 26945 21867 26979
rect 22107 26945 22141 26979
rect 23489 26945 23523 26979
rect 23765 26945 23799 26979
rect 24133 26945 24167 26979
rect 24225 26945 24259 26979
rect 4537 26877 4571 26911
rect 7757 26877 7791 26911
rect 13001 26877 13035 26911
rect 13461 26877 13495 26911
rect 13737 26877 13771 26911
rect 14013 26877 14047 26911
rect 16681 26877 16715 26911
rect 17325 26877 17359 26911
rect 17601 26877 17635 26911
rect 17739 26877 17773 26911
rect 23581 26809 23615 26843
rect 15761 26741 15795 26775
rect 18521 26741 18555 26775
rect 24409 26741 24443 26775
rect 2605 26537 2639 26571
rect 3249 26537 3283 26571
rect 3985 26537 4019 26571
rect 11069 26537 11103 26571
rect 16773 26537 16807 26571
rect 22753 26537 22787 26571
rect 3157 26469 3191 26503
rect 9873 26469 9907 26503
rect 15945 26469 15979 26503
rect 19073 26469 19107 26503
rect 1593 26401 1627 26435
rect 6561 26401 6595 26435
rect 9229 26401 9263 26435
rect 10266 26401 10300 26435
rect 16313 26401 16347 26435
rect 17693 26401 17727 26435
rect 1851 26303 1885 26337
rect 2973 26333 3007 26367
rect 3433 26333 3467 26367
rect 3801 26333 3835 26367
rect 6835 26333 6869 26367
rect 9413 26333 9447 26367
rect 10149 26333 10183 26367
rect 10425 26333 10459 26367
rect 11805 26333 11839 26367
rect 11897 26333 11931 26367
rect 14933 26333 14967 26367
rect 15207 26333 15241 26367
rect 16497 26333 16531 26367
rect 17960 26333 17994 26367
rect 19441 26333 19475 26367
rect 22937 26333 22971 26367
rect 23489 26333 23523 26367
rect 23673 26333 23707 26367
rect 12265 26265 12299 26299
rect 16865 26265 16899 26299
rect 23857 26265 23891 26299
rect 24225 26265 24259 26299
rect 7573 26197 7607 26231
rect 11529 26197 11563 26231
rect 12633 26197 12667 26231
rect 12817 26197 12851 26231
rect 19257 26197 19291 26231
rect 23673 26197 23707 26231
rect 2513 25993 2547 26027
rect 3065 25993 3099 26027
rect 3341 25993 3375 26027
rect 15669 25993 15703 26027
rect 16037 25993 16071 26027
rect 22385 25993 22419 26027
rect 23489 25993 23523 26027
rect 23949 25993 23983 26027
rect 7113 25925 7147 25959
rect 7849 25925 7883 25959
rect 8217 25925 8251 25959
rect 24133 25925 24167 25959
rect 1501 25857 1535 25891
rect 1775 25857 1809 25891
rect 2881 25857 2915 25891
rect 3157 25857 3191 25891
rect 3707 25857 3741 25891
rect 5087 25857 5121 25891
rect 6837 25857 6871 25891
rect 7389 25857 7423 25891
rect 7481 25857 7515 25891
rect 11529 25857 11563 25891
rect 11803 25857 11837 25891
rect 13277 25857 13311 25891
rect 14013 25857 14047 25891
rect 14289 25857 14323 25891
rect 14933 25857 14967 25891
rect 15485 25857 15519 25891
rect 15577 25857 15611 25891
rect 15853 25857 15887 25891
rect 16037 25857 16071 25891
rect 18855 25857 18889 25891
rect 19993 25857 20027 25891
rect 20361 25857 20395 25891
rect 20545 25857 20579 25891
rect 21373 25857 21407 25891
rect 21557 25857 21591 25891
rect 22569 25857 22603 25891
rect 23029 25857 23063 25891
rect 23673 25857 23707 25891
rect 23765 25857 23799 25891
rect 3433 25789 3467 25823
rect 4813 25789 4847 25823
rect 9045 25789 9079 25823
rect 9229 25789 9263 25823
rect 9965 25789 9999 25823
rect 10082 25789 10116 25823
rect 10241 25789 10275 25823
rect 13093 25789 13127 25823
rect 13737 25789 13771 25823
rect 14151 25789 14185 25823
rect 18613 25789 18647 25823
rect 20269 25789 20303 25823
rect 20453 25789 20487 25823
rect 9689 25721 9723 25755
rect 10885 25721 10919 25755
rect 15301 25721 15335 25755
rect 19625 25721 19659 25755
rect 4445 25653 4479 25687
rect 5825 25653 5859 25687
rect 8401 25653 8435 25687
rect 12541 25653 12575 25687
rect 20085 25653 20119 25687
rect 20177 25653 20211 25687
rect 21465 25653 21499 25687
rect 23121 25653 23155 25687
rect 24409 25653 24443 25687
rect 1593 25449 1627 25483
rect 8309 25449 8343 25483
rect 10517 25449 10551 25483
rect 19349 25449 19383 25483
rect 21373 25449 21407 25483
rect 23489 25449 23523 25483
rect 3341 25381 3375 25415
rect 19625 25381 19659 25415
rect 23213 25381 23247 25415
rect 2329 25313 2363 25347
rect 5457 25313 5491 25347
rect 7297 25313 7331 25347
rect 16681 25313 16715 25347
rect 16865 25313 16899 25347
rect 17325 25313 17359 25347
rect 17718 25313 17752 25347
rect 20361 25313 20395 25347
rect 23673 25313 23707 25347
rect 1409 25245 1443 25279
rect 1685 25245 1719 25279
rect 2145 25245 2179 25279
rect 2571 25245 2605 25279
rect 4721 25245 4755 25279
rect 5731 25245 5765 25279
rect 7571 25245 7605 25279
rect 9505 25245 9539 25279
rect 9779 25245 9813 25279
rect 11713 25245 11747 25279
rect 11805 25245 11839 25279
rect 17601 25245 17635 25279
rect 17877 25245 17911 25279
rect 19257 25245 19291 25279
rect 19809 25245 19843 25279
rect 20619 25215 20653 25249
rect 21833 25245 21867 25279
rect 23397 25245 23431 25279
rect 4261 25177 4295 25211
rect 4353 25177 4387 25211
rect 12173 25177 12207 25211
rect 22100 25177 22134 25211
rect 23857 25177 23891 25211
rect 24225 25177 24259 25211
rect 1869 25109 1903 25143
rect 1961 25109 1995 25143
rect 3985 25109 4019 25143
rect 5089 25109 5123 25143
rect 5273 25109 5307 25143
rect 6469 25109 6503 25143
rect 11437 25109 11471 25143
rect 12541 25109 12575 25143
rect 12725 25109 12759 25143
rect 18521 25109 18555 25143
rect 23673 25109 23707 25143
rect 1593 24905 1627 24939
rect 3985 24905 4019 24939
rect 17693 24905 17727 24939
rect 21833 24905 21867 24939
rect 23489 24905 23523 24939
rect 2881 24837 2915 24871
rect 3617 24837 3651 24871
rect 1409 24769 1443 24803
rect 1685 24769 1719 24803
rect 1961 24769 1995 24803
rect 2237 24769 2271 24803
rect 3157 24769 3191 24803
rect 3249 24769 3283 24803
rect 4353 24769 4387 24803
rect 6193 24769 6227 24803
rect 8767 24769 8801 24803
rect 12447 24769 12481 24803
rect 16955 24769 16989 24803
rect 18061 24769 18095 24803
rect 18303 24769 18337 24803
rect 20157 24769 20191 24803
rect 21373 24769 21407 24803
rect 22017 24769 22051 24803
rect 22719 24769 22753 24803
rect 24133 24769 24167 24803
rect 4537 24701 4571 24735
rect 5273 24701 5307 24735
rect 5411 24701 5445 24735
rect 5549 24701 5583 24735
rect 8493 24701 8527 24735
rect 12173 24701 12207 24735
rect 16681 24701 16715 24735
rect 19901 24701 19935 24735
rect 21649 24701 21683 24735
rect 22477 24701 22511 24735
rect 2145 24633 2179 24667
rect 4997 24633 5031 24667
rect 9505 24633 9539 24667
rect 21281 24633 21315 24667
rect 1869 24565 1903 24599
rect 2421 24565 2455 24599
rect 4169 24565 4203 24599
rect 13185 24565 13219 24599
rect 19073 24565 19107 24599
rect 21465 24565 21499 24599
rect 21557 24565 21591 24599
rect 24409 24565 24443 24599
rect 2881 24361 2915 24395
rect 7021 24361 7055 24395
rect 17969 24361 18003 24395
rect 19533 24361 19567 24395
rect 21005 24361 21039 24395
rect 23397 24361 23431 24395
rect 5825 24293 5859 24327
rect 7113 24293 7147 24327
rect 23857 24293 23891 24327
rect 5181 24225 5215 24259
rect 6218 24225 6252 24259
rect 6377 24225 6411 24259
rect 10609 24225 10643 24259
rect 12633 24225 12667 24259
rect 15025 24225 15059 24259
rect 15209 24225 15243 24259
rect 15669 24225 15703 24259
rect 16221 24225 16255 24259
rect 16957 24225 16991 24259
rect 1961 24157 1995 24191
rect 5365 24157 5399 24191
rect 6101 24157 6135 24191
rect 7297 24157 7331 24191
rect 7481 24157 7515 24191
rect 7941 24157 7975 24191
rect 8953 24157 8987 24191
rect 9227 24157 9261 24191
rect 10883 24157 10917 24191
rect 12907 24157 12941 24191
rect 15945 24157 15979 24191
rect 16062 24157 16096 24191
rect 17199 24157 17233 24191
rect 19717 24157 19751 24191
rect 19809 24157 19843 24191
rect 19993 24157 20027 24191
rect 20545 24157 20579 24191
rect 20913 24157 20947 24191
rect 23581 24157 23615 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 1593 24089 1627 24123
rect 1869 24089 1903 24123
rect 2329 24089 2363 24123
rect 2697 24089 2731 24123
rect 7573 24021 7607 24055
rect 7757 24021 7791 24055
rect 9965 24021 9999 24055
rect 11621 24021 11655 24055
rect 13645 24021 13679 24055
rect 16865 24021 16899 24055
rect 19901 24021 19935 24055
rect 20361 24021 20395 24055
rect 24133 24021 24167 24055
rect 3525 23817 3559 23851
rect 4077 23817 4111 23851
rect 9965 23817 9999 23851
rect 15669 23817 15703 23851
rect 19257 23817 19291 23851
rect 22845 23817 22879 23851
rect 8861 23749 8895 23783
rect 9137 23749 9171 23783
rect 9229 23749 9263 23783
rect 24133 23749 24167 23783
rect 2787 23681 2821 23715
rect 3893 23681 3927 23715
rect 6929 23681 6963 23715
rect 7203 23681 7237 23715
rect 8309 23681 8343 23715
rect 8493 23681 8527 23715
rect 9597 23681 9631 23715
rect 11897 23681 11931 23715
rect 12633 23681 12667 23715
rect 13691 23681 13725 23715
rect 13829 23681 13863 23715
rect 14899 23681 14933 23715
rect 16221 23681 16255 23715
rect 17877 23681 17911 23715
rect 18133 23681 18167 23715
rect 19623 23691 19657 23725
rect 23029 23681 23063 23715
rect 23213 23681 23247 23715
rect 23397 23681 23431 23715
rect 23489 23681 23523 23715
rect 23949 23681 23983 23715
rect 1409 23613 1443 23647
rect 1685 23613 1719 23647
rect 2513 23613 2547 23647
rect 12817 23613 12851 23647
rect 13277 23613 13311 23647
rect 13553 23613 13587 23647
rect 14657 23613 14691 23647
rect 19349 23613 19383 23647
rect 10149 23545 10183 23579
rect 23765 23545 23799 23579
rect 7941 23477 7975 23511
rect 8401 23477 8435 23511
rect 12081 23477 12115 23511
rect 14473 23477 14507 23511
rect 20361 23477 20395 23511
rect 23305 23477 23339 23511
rect 23581 23477 23615 23511
rect 24409 23477 24443 23511
rect 2421 23273 2455 23307
rect 2973 23273 3007 23307
rect 23765 23273 23799 23307
rect 18429 23205 18463 23239
rect 7941 23137 7975 23171
rect 14105 23137 14139 23171
rect 19349 23137 19383 23171
rect 19717 23137 19751 23171
rect 19901 23137 19935 23171
rect 1409 23069 1443 23103
rect 1683 23069 1717 23103
rect 2789 23069 2823 23103
rect 3065 23069 3099 23103
rect 7849 23069 7883 23103
rect 8217 23069 8251 23103
rect 10885 23069 10919 23103
rect 10977 23069 11011 23103
rect 11345 23069 11379 23103
rect 14379 23069 14413 23103
rect 18613 23069 18647 23103
rect 19257 23069 19291 23103
rect 19625 23069 19659 23103
rect 20637 23069 20671 23103
rect 22109 23069 22143 23103
rect 22385 23069 22419 23103
rect 22652 23069 22686 23103
rect 23949 23069 23983 23103
rect 8125 23001 8159 23035
rect 10149 23001 10183 23035
rect 11713 23001 11747 23035
rect 20882 23001 20916 23035
rect 3249 22933 3283 22967
rect 10609 22933 10643 22967
rect 11897 22933 11931 22967
rect 15117 22933 15151 22967
rect 19901 22933 19935 22967
rect 22017 22933 22051 22967
rect 22201 22933 22235 22967
rect 24133 22933 24167 22967
rect 3801 22729 3835 22763
rect 9689 22729 9723 22763
rect 11069 22729 11103 22763
rect 21097 22729 21131 22763
rect 24225 22729 24259 22763
rect 1667 22623 1701 22657
rect 2789 22593 2823 22627
rect 3063 22593 3097 22627
rect 4169 22593 4203 22627
rect 4443 22593 4477 22627
rect 6619 22593 6653 22627
rect 8935 22623 8969 22657
rect 10331 22593 10365 22627
rect 16865 22593 16899 22627
rect 17739 22593 17773 22627
rect 21281 22593 21315 22627
rect 21465 22593 21499 22627
rect 21649 22593 21683 22627
rect 21833 22593 21867 22627
rect 22107 22603 22141 22637
rect 23213 22593 23247 22627
rect 23487 22593 23521 22627
rect 1409 22525 1443 22559
rect 6377 22525 6411 22559
rect 8677 22525 8711 22559
rect 10057 22525 10091 22559
rect 16681 22525 16715 22559
rect 17601 22525 17635 22559
rect 17877 22525 17911 22559
rect 17325 22457 17359 22491
rect 2421 22389 2455 22423
rect 5181 22389 5215 22423
rect 7389 22389 7423 22423
rect 14841 22389 14875 22423
rect 18521 22389 18555 22423
rect 21557 22389 21591 22423
rect 22845 22389 22879 22423
rect 3065 22185 3099 22219
rect 3985 22185 4019 22219
rect 11069 22185 11103 22219
rect 22109 22185 22143 22219
rect 23213 22185 23247 22219
rect 6009 22117 6043 22151
rect 6561 22117 6595 22151
rect 12909 22117 12943 22151
rect 17325 22117 17359 22151
rect 22385 22117 22419 22151
rect 6653 22049 6687 22083
rect 14749 22049 14783 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 22293 22049 22327 22083
rect 23397 22049 23431 22083
rect 2145 21981 2179 22015
rect 2513 21981 2547 22015
rect 3249 21981 3283 22015
rect 3801 21981 3835 22015
rect 4997 21981 5031 22015
rect 5089 21981 5123 22015
rect 6927 21981 6961 22015
rect 10057 21981 10091 22015
rect 10331 21981 10365 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 15142 21981 15176 22015
rect 16313 21981 16347 22015
rect 16587 21981 16621 22015
rect 18429 21981 18463 22015
rect 19257 21981 19291 22015
rect 19524 21981 19558 22015
rect 20821 21981 20855 22015
rect 21005 21981 21039 22015
rect 22017 21981 22051 22015
rect 22569 21981 22603 22015
rect 23121 21981 23155 22015
rect 23581 21981 23615 22015
rect 24225 21981 24259 22015
rect 1777 21913 1811 21947
rect 2053 21913 2087 21947
rect 5457 21913 5491 21947
rect 11897 21913 11931 21947
rect 11989 21913 12023 21947
rect 12357 21913 12391 21947
rect 23949 21913 23983 21947
rect 2881 21845 2915 21879
rect 3433 21845 3467 21879
rect 4721 21845 4755 21879
rect 5825 21845 5859 21879
rect 7665 21845 7699 21879
rect 11621 21845 11655 21879
rect 12725 21845 12759 21879
rect 15945 21845 15979 21879
rect 18245 21845 18279 21879
rect 20637 21845 20671 21879
rect 21005 21845 21039 21879
rect 22293 21845 22327 21879
rect 23397 21845 23431 21879
rect 24041 21845 24075 21879
rect 2421 21641 2455 21675
rect 2973 21641 3007 21675
rect 5733 21641 5767 21675
rect 9597 21641 9631 21675
rect 9781 21641 9815 21675
rect 12817 21641 12851 21675
rect 14289 21641 14323 21675
rect 20913 21641 20947 21675
rect 22017 21641 22051 21675
rect 24409 21641 24443 21675
rect 6561 21573 6595 21607
rect 6837 21573 6871 21607
rect 6929 21573 6963 21607
rect 7665 21573 7699 21607
rect 8493 21573 8527 21607
rect 24133 21573 24167 21607
rect 1409 21505 1443 21539
rect 1667 21535 1701 21569
rect 2789 21505 2823 21539
rect 3065 21505 3099 21539
rect 4721 21505 4755 21539
rect 4995 21505 5029 21539
rect 7297 21505 7331 21539
rect 8769 21505 8803 21539
rect 8861 21505 8895 21539
rect 9229 21505 9263 21539
rect 12047 21505 12081 21539
rect 13551 21505 13585 21539
rect 15375 21505 15409 21539
rect 16681 21505 16715 21539
rect 17601 21505 17635 21539
rect 17877 21505 17911 21539
rect 18521 21505 18555 21539
rect 18797 21505 18831 21539
rect 18889 21505 18923 21539
rect 19809 21505 19843 21539
rect 20143 21505 20177 21539
rect 21281 21505 21315 21539
rect 21833 21505 21867 21539
rect 23397 21505 23431 21539
rect 23581 21505 23615 21539
rect 23673 21505 23707 21539
rect 11805 21437 11839 21471
rect 13277 21437 13311 21471
rect 15117 21437 15151 21471
rect 16865 21437 16899 21471
rect 17718 21437 17752 21471
rect 19901 21437 19935 21471
rect 21557 21437 21591 21471
rect 3249 21369 3283 21403
rect 7849 21369 7883 21403
rect 17325 21369 17359 21403
rect 18613 21369 18647 21403
rect 21465 21369 21499 21403
rect 15025 21301 15059 21335
rect 16129 21301 16163 21335
rect 18981 21301 19015 21335
rect 19625 21301 19659 21335
rect 21373 21301 21407 21335
rect 23489 21301 23523 21335
rect 23857 21301 23891 21335
rect 2513 21097 2547 21131
rect 8493 21097 8527 21131
rect 9965 21097 9999 21131
rect 17969 21097 18003 21131
rect 20453 21097 20487 21131
rect 2789 21029 2823 21063
rect 20729 21029 20763 21063
rect 10333 20961 10367 20995
rect 14749 20961 14783 20995
rect 15393 20961 15427 20995
rect 15669 20961 15703 20995
rect 15945 20961 15979 20995
rect 16957 20961 16991 20995
rect 18889 20961 18923 20995
rect 22569 20961 22603 20995
rect 1409 20893 1443 20927
rect 1685 20893 1719 20927
rect 2329 20893 2363 20927
rect 2605 20893 2639 20927
rect 3801 20893 3835 20927
rect 4075 20893 4109 20927
rect 7481 20893 7515 20927
rect 7723 20893 7757 20927
rect 8953 20893 8987 20927
rect 9195 20893 9229 20927
rect 10575 20893 10609 20927
rect 11989 20893 12023 20927
rect 12231 20893 12265 20927
rect 14933 20893 14967 20927
rect 15786 20893 15820 20927
rect 17199 20893 17233 20927
rect 18705 20893 18739 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 20361 20893 20395 20927
rect 20913 20893 20947 20927
rect 22825 20893 22859 20927
rect 24041 20893 24075 20927
rect 18981 20825 19015 20859
rect 19073 20825 19107 20859
rect 19349 20825 19383 20859
rect 4813 20757 4847 20791
rect 11345 20757 11379 20791
rect 13001 20757 13035 20791
rect 16589 20757 16623 20791
rect 23949 20757 23983 20791
rect 24133 20757 24167 20791
rect 15393 20553 15427 20587
rect 18797 20553 18831 20587
rect 23765 20553 23799 20587
rect 9965 20485 9999 20519
rect 10701 20485 10735 20519
rect 11069 20485 11103 20519
rect 1683 20417 1717 20451
rect 3918 20417 3952 20451
rect 4077 20417 4111 20451
rect 4813 20417 4847 20451
rect 5087 20417 5121 20451
rect 10241 20417 10275 20451
rect 10333 20417 10367 20451
rect 12357 20417 12391 20451
rect 13394 20417 13428 20451
rect 13553 20417 13587 20451
rect 14381 20417 14415 20451
rect 14623 20417 14657 20451
rect 17785 20417 17819 20451
rect 18059 20417 18093 20451
rect 22385 20417 22419 20451
rect 22661 20417 22695 20451
rect 23011 20447 23045 20481
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 1409 20349 1443 20383
rect 2881 20349 2915 20383
rect 3065 20349 3099 20383
rect 3801 20349 3835 20383
rect 12541 20349 12575 20383
rect 13001 20349 13035 20383
rect 13277 20349 13311 20383
rect 22753 20349 22787 20383
rect 24409 20349 24443 20383
rect 3525 20281 3559 20315
rect 22201 20281 22235 20315
rect 2421 20213 2455 20247
rect 4721 20213 4755 20247
rect 5825 20213 5859 20247
rect 11253 20213 11287 20247
rect 14197 20213 14231 20247
rect 22477 20213 22511 20247
rect 24317 20213 24351 20247
rect 1593 20009 1627 20043
rect 3341 20009 3375 20043
rect 3985 20009 4019 20043
rect 7665 20009 7699 20043
rect 11161 20009 11195 20043
rect 13553 20009 13587 20043
rect 22109 20009 22143 20043
rect 23949 20009 23983 20043
rect 2329 19873 2363 19907
rect 6653 19873 6687 19907
rect 12541 19873 12575 19907
rect 15853 19873 15887 19907
rect 16313 19873 16347 19907
rect 16589 19873 16623 19907
rect 22201 19873 22235 19907
rect 1501 19805 1535 19839
rect 2603 19805 2637 19839
rect 3801 19805 3835 19839
rect 4905 19805 4939 19839
rect 5917 19805 5951 19839
rect 6927 19805 6961 19839
rect 8217 19805 8251 19839
rect 10149 19805 10183 19839
rect 10423 19805 10457 19839
rect 12815 19805 12849 19839
rect 15669 19805 15703 19839
rect 16727 19805 16761 19839
rect 16865 19805 16899 19839
rect 19073 19805 19107 19839
rect 19257 19805 19291 19839
rect 20729 19805 20763 19839
rect 20985 19805 21019 19839
rect 22443 19805 22477 19839
rect 23673 19805 23707 19839
rect 5135 19737 5169 19771
rect 5457 19737 5491 19771
rect 5549 19737 5583 19771
rect 6285 19737 6319 19771
rect 19502 19737 19536 19771
rect 6469 19669 6503 19703
rect 17509 19669 17543 19703
rect 18889 19669 18923 19703
rect 20637 19669 20671 19703
rect 23213 19669 23247 19703
rect 1593 19465 1627 19499
rect 3065 19465 3099 19499
rect 3525 19465 3559 19499
rect 5917 19465 5951 19499
rect 7113 19465 7147 19499
rect 17693 19465 17727 19499
rect 20177 19465 20211 19499
rect 20821 19465 20855 19499
rect 21189 19465 21223 19499
rect 22385 19465 22419 19499
rect 8217 19397 8251 19431
rect 23581 19397 23615 19431
rect 24133 19397 24167 19431
rect 1409 19329 1443 19363
rect 1959 19329 1993 19363
rect 3249 19329 3283 19363
rect 3341 19329 3375 19363
rect 4905 19329 4939 19363
rect 5179 19329 5213 19363
rect 7389 19329 7423 19363
rect 7481 19329 7515 19363
rect 7849 19329 7883 19363
rect 8861 19329 8895 19363
rect 9135 19329 9169 19363
rect 11803 19329 11837 19363
rect 13461 19329 13495 19363
rect 13735 19329 13769 19363
rect 16681 19329 16715 19363
rect 16939 19359 16973 19393
rect 19165 19329 19199 19363
rect 19407 19329 19441 19363
rect 20545 19329 20579 19363
rect 20913 19329 20947 19363
rect 21097 19329 21131 19363
rect 21373 19329 21407 19363
rect 21833 19329 21867 19363
rect 21925 19329 21959 19363
rect 22109 19329 22143 19363
rect 22477 19329 22511 19363
rect 22661 19329 22695 19363
rect 23397 19329 23431 19363
rect 1685 19261 1719 19295
rect 11529 19261 11563 19295
rect 16497 19261 16531 19295
rect 20821 19261 20855 19295
rect 21005 19261 21039 19295
rect 22201 19261 22235 19295
rect 22385 19261 22419 19295
rect 22569 19261 22603 19295
rect 24409 19261 24443 19295
rect 8401 19193 8435 19227
rect 23213 19193 23247 19227
rect 2697 19125 2731 19159
rect 9873 19125 9907 19159
rect 12541 19125 12575 19159
rect 14473 19125 14507 19159
rect 20637 19125 20671 19159
rect 23857 19125 23891 19159
rect 8125 18921 8159 18955
rect 17049 18921 17083 18955
rect 19717 18921 19751 18955
rect 3249 18853 3283 18887
rect 4813 18853 4847 18887
rect 10425 18853 10459 18887
rect 14749 18853 14783 18887
rect 19993 18853 20027 18887
rect 23581 18853 23615 18887
rect 1593 18785 1627 18819
rect 7113 18785 7147 18819
rect 14105 18785 14139 18819
rect 15025 18785 15059 18819
rect 15142 18785 15176 18819
rect 16037 18785 16071 18819
rect 22845 18785 22879 18819
rect 1867 18717 1901 18751
rect 3801 18717 3835 18751
rect 4059 18707 4093 18741
rect 7387 18717 7421 18751
rect 9413 18717 9447 18751
rect 11253 18717 11287 18751
rect 11527 18717 11561 18751
rect 14289 18717 14323 18751
rect 15301 18717 15335 18751
rect 16295 18687 16329 18721
rect 17601 18717 17635 18751
rect 17859 18687 17893 18721
rect 19625 18717 19659 18751
rect 20177 18717 20211 18751
rect 22753 18717 22787 18751
rect 22937 18717 22971 18751
rect 23213 18717 23247 18751
rect 23397 18717 23431 18751
rect 23857 18717 23891 18751
rect 24225 18717 24259 18751
rect 3065 18649 3099 18683
rect 9137 18649 9171 18683
rect 9505 18649 9539 18683
rect 9873 18649 9907 18683
rect 10241 18649 10275 18683
rect 2605 18581 2639 18615
rect 12265 18581 12299 18615
rect 15945 18581 15979 18615
rect 18613 18581 18647 18615
rect 23029 18581 23063 18615
rect 1869 18377 1903 18411
rect 5549 18377 5583 18411
rect 9229 18377 9263 18411
rect 15209 18377 15243 18411
rect 3525 18309 3559 18343
rect 11713 18309 11747 18343
rect 12081 18309 12115 18343
rect 12817 18309 12851 18343
rect 22814 18309 22848 18343
rect 24133 18309 24167 18343
rect 1777 18241 1811 18275
rect 2327 18241 2361 18275
rect 4259 18241 4293 18275
rect 5457 18241 5491 18275
rect 8217 18241 8251 18275
rect 8491 18241 8525 18275
rect 9855 18271 9889 18305
rect 11345 18241 11379 18275
rect 11989 18241 12023 18275
rect 12449 18241 12483 18275
rect 14197 18241 14231 18275
rect 14471 18241 14505 18275
rect 17141 18241 17175 18275
rect 17325 18241 17359 18275
rect 18337 18241 18371 18275
rect 2053 18173 2087 18207
rect 3985 18173 4019 18207
rect 9597 18173 9631 18207
rect 18061 18173 18095 18207
rect 18199 18173 18233 18207
rect 22569 18173 22603 18207
rect 13001 18105 13035 18139
rect 17785 18105 17819 18139
rect 3065 18037 3099 18071
rect 3617 18037 3651 18071
rect 4997 18037 5031 18071
rect 10609 18037 10643 18071
rect 18981 18037 19015 18071
rect 23949 18037 23983 18071
rect 24409 18037 24443 18071
rect 18153 17833 18187 17867
rect 23765 17833 23799 17867
rect 2421 17765 2455 17799
rect 4445 17765 4479 17799
rect 6009 17765 6043 17799
rect 10425 17765 10459 17799
rect 18705 17765 18739 17799
rect 22109 17765 22143 17799
rect 1961 17697 1995 17731
rect 3801 17697 3835 17731
rect 4721 17697 4755 17731
rect 6101 17697 6135 17731
rect 9781 17697 9815 17731
rect 10818 17697 10852 17731
rect 12265 17697 12299 17731
rect 12725 17697 12759 17731
rect 13001 17697 13035 17731
rect 14289 17697 14323 17731
rect 22753 17697 22787 17731
rect 1409 17629 1443 17663
rect 1777 17629 1811 17663
rect 2697 17629 2731 17663
rect 2814 17629 2848 17663
rect 2973 17629 3007 17663
rect 3985 17629 4019 17663
rect 4859 17629 4893 17663
rect 4997 17629 5031 17663
rect 6375 17629 6409 17663
rect 9965 17629 9999 17663
rect 10701 17629 10735 17663
rect 10977 17629 11011 17663
rect 11621 17629 11655 17663
rect 11713 17629 11747 17663
rect 12081 17629 12115 17663
rect 13118 17629 13152 17663
rect 13277 17629 13311 17663
rect 17141 17629 17175 17663
rect 17383 17629 17417 17663
rect 19257 17629 19291 17663
rect 19524 17629 19558 17663
rect 20729 17629 20763 17663
rect 22201 17629 22235 17663
rect 22661 17629 22695 17663
rect 23011 17599 23045 17633
rect 20985 17561 21019 17595
rect 1593 17493 1627 17527
rect 3617 17493 3651 17527
rect 5641 17493 5675 17527
rect 7113 17493 7147 17527
rect 11897 17493 11931 17527
rect 13921 17493 13955 17527
rect 20637 17493 20671 17527
rect 22293 17493 22327 17527
rect 22477 17493 22511 17527
rect 7665 17289 7699 17323
rect 11069 17289 11103 17323
rect 13645 17289 13679 17323
rect 19533 17289 19567 17323
rect 21005 17289 21039 17323
rect 23581 17289 23615 17323
rect 6561 17221 6595 17255
rect 6929 17221 6963 17255
rect 1593 17153 1627 17187
rect 1685 17153 1719 17187
rect 2881 17153 2915 17187
rect 3801 17153 3835 17187
rect 5147 17153 5181 17187
rect 6837 17153 6871 17187
rect 7297 17153 7331 17187
rect 10057 17153 10091 17187
rect 10331 17153 10365 17187
rect 12265 17153 12299 17187
rect 12633 17153 12667 17187
rect 12907 17153 12941 17187
rect 15451 17153 15485 17187
rect 16923 17153 16957 17187
rect 19717 17153 19751 17187
rect 20085 17153 20119 17187
rect 20729 17153 20763 17187
rect 21189 17153 21223 17187
rect 21465 17153 21499 17187
rect 21649 17153 21683 17187
rect 22075 17153 22109 17187
rect 23397 17153 23431 17187
rect 23857 17153 23891 17187
rect 24317 17153 24351 17187
rect 1869 17085 1903 17119
rect 2329 17085 2363 17119
rect 2605 17085 2639 17119
rect 2743 17085 2777 17119
rect 4905 17085 4939 17119
rect 15209 17085 15243 17119
rect 16681 17085 16715 17119
rect 21833 17085 21867 17119
rect 5917 17017 5951 17051
rect 7849 17017 7883 17051
rect 1409 16949 1443 16983
rect 3525 16949 3559 16983
rect 3617 16949 3651 16983
rect 12449 16949 12483 16983
rect 14473 16949 14507 16983
rect 16221 16949 16255 16983
rect 17693 16949 17727 16983
rect 20177 16949 20211 16983
rect 20545 16949 20579 16983
rect 21557 16949 21591 16983
rect 22845 16949 22879 16983
rect 24133 16949 24167 16983
rect 24409 16949 24443 16983
rect 1961 16745 1995 16779
rect 3985 16745 4019 16779
rect 8769 16745 8803 16779
rect 15577 16745 15611 16779
rect 21281 16745 21315 16779
rect 13645 16677 13679 16711
rect 16405 16677 16439 16711
rect 22017 16677 22051 16711
rect 6929 16609 6963 16643
rect 7573 16609 7607 16643
rect 7966 16609 8000 16643
rect 8125 16609 8159 16643
rect 12633 16609 12667 16643
rect 15761 16609 15795 16643
rect 15945 16609 15979 16643
rect 16798 16609 16832 16643
rect 16957 16609 16991 16643
rect 19809 16609 19843 16643
rect 21465 16609 21499 16643
rect 22201 16609 22235 16643
rect 23949 16609 23983 16643
rect 1409 16541 1443 16575
rect 2421 16541 2455 16575
rect 3617 16541 3651 16575
rect 7113 16541 7147 16575
rect 7849 16541 7883 16575
rect 12875 16541 12909 16575
rect 14565 16541 14599 16575
rect 15025 16541 15059 16575
rect 16681 16541 16715 16575
rect 17601 16541 17635 16575
rect 17693 16541 17727 16575
rect 20051 16531 20085 16565
rect 21189 16541 21223 16575
rect 21925 16541 21959 16575
rect 23489 16541 23523 16575
rect 23673 16541 23707 16575
rect 1869 16473 1903 16507
rect 2973 16473 3007 16507
rect 3893 16473 3927 16507
rect 14657 16473 14691 16507
rect 22201 16473 22235 16507
rect 1593 16405 1627 16439
rect 2697 16405 2731 16439
rect 3065 16405 3099 16439
rect 3433 16405 3467 16439
rect 14289 16405 14323 16439
rect 15393 16405 15427 16439
rect 17877 16405 17911 16439
rect 20821 16405 20855 16439
rect 21465 16405 21499 16439
rect 23305 16405 23339 16439
rect 1777 16201 1811 16235
rect 5365 16201 5399 16235
rect 8493 16201 8527 16235
rect 13093 16201 13127 16235
rect 15393 16201 15427 16235
rect 19257 16201 19291 16235
rect 20821 16201 20855 16235
rect 24317 16201 24351 16235
rect 1685 16133 1719 16167
rect 18122 16133 18156 16167
rect 2145 16065 2179 16099
rect 2403 16095 2437 16129
rect 3525 16065 3559 16099
rect 4445 16065 4479 16099
rect 4562 16065 4596 16099
rect 7739 16065 7773 16099
rect 8861 16065 8895 16099
rect 9135 16065 9169 16099
rect 10609 16065 10643 16099
rect 12081 16065 12115 16099
rect 12339 16095 12373 16129
rect 14623 16065 14657 16099
rect 19349 16065 19383 16099
rect 19809 16065 19843 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 22903 16065 22937 16099
rect 24041 16065 24075 16099
rect 24133 16065 24167 16099
rect 3709 15997 3743 16031
rect 4721 15997 4755 16031
rect 7481 15997 7515 16031
rect 14381 15997 14415 16031
rect 17877 15997 17911 16031
rect 22661 15997 22695 16031
rect 24317 15997 24351 16031
rect 3157 15929 3191 15963
rect 4169 15929 4203 15963
rect 10425 15929 10459 15963
rect 9873 15861 9907 15895
rect 19441 15861 19475 15895
rect 19625 15861 19659 15895
rect 23673 15861 23707 15895
rect 2881 15657 2915 15691
rect 4813 15657 4847 15691
rect 7849 15657 7883 15691
rect 10793 15657 10827 15691
rect 18337 15657 18371 15691
rect 24133 15657 24167 15691
rect 9597 15589 9631 15623
rect 3801 15521 3835 15555
rect 5457 15521 5491 15555
rect 6837 15521 6871 15555
rect 8953 15521 8987 15555
rect 9990 15521 10024 15555
rect 22385 15521 22419 15555
rect 3433 15453 3467 15487
rect 4043 15453 4077 15487
rect 5699 15453 5733 15487
rect 7111 15453 7145 15487
rect 9137 15453 9171 15487
rect 9873 15453 9907 15487
rect 10149 15453 10183 15487
rect 10885 15453 10919 15487
rect 11159 15453 11193 15487
rect 18521 15453 18555 15487
rect 19257 15453 19291 15487
rect 19499 15443 19533 15477
rect 22293 15453 22327 15487
rect 23949 15453 23983 15487
rect 1869 15385 1903 15419
rect 2237 15385 2271 15419
rect 2789 15385 2823 15419
rect 22630 15385 22664 15419
rect 2329 15317 2363 15351
rect 3249 15317 3283 15351
rect 6469 15317 6503 15351
rect 11897 15317 11931 15351
rect 20269 15317 20303 15351
rect 22109 15317 22143 15351
rect 23765 15317 23799 15351
rect 1593 15113 1627 15147
rect 10241 15113 10275 15147
rect 12817 15113 12851 15147
rect 13001 15113 13035 15147
rect 19717 15113 19751 15147
rect 3341 15045 3375 15079
rect 11713 15045 11747 15079
rect 11989 15045 12023 15079
rect 17408 15045 17442 15079
rect 23765 15045 23799 15079
rect 1777 14977 1811 15011
rect 1869 14977 1903 15011
rect 2143 14977 2177 15011
rect 3893 14977 3927 15011
rect 4353 14977 4387 15011
rect 4611 15007 4645 15041
rect 6561 14977 6595 15011
rect 7435 14977 7469 15011
rect 9503 14977 9537 15011
rect 12081 14977 12115 15011
rect 12449 14977 12483 15011
rect 14195 14987 14229 15021
rect 17141 14977 17175 15011
rect 19441 14977 19475 15011
rect 19533 14977 19567 15011
rect 19809 14977 19843 15011
rect 19993 14977 20027 15011
rect 20269 14977 20303 15011
rect 20525 14977 20559 15011
rect 22075 14977 22109 15011
rect 23397 14977 23431 15011
rect 24225 14977 24259 15011
rect 6377 14909 6411 14943
rect 7021 14909 7055 14943
rect 7297 14909 7331 14943
rect 7573 14909 7607 14943
rect 9229 14909 9263 14943
rect 13921 14909 13955 14943
rect 19717 14909 19751 14943
rect 19901 14909 19935 14943
rect 21833 14909 21867 14943
rect 24501 14909 24535 14943
rect 23489 14841 23523 14875
rect 24317 14841 24351 14875
rect 2881 14773 2915 14807
rect 3433 14773 3467 14807
rect 3985 14773 4019 14807
rect 5365 14773 5399 14807
rect 8217 14773 8251 14807
rect 14933 14773 14967 14807
rect 18521 14773 18555 14807
rect 21649 14773 21683 14807
rect 22845 14773 22879 14807
rect 24041 14773 24075 14807
rect 24409 14773 24443 14807
rect 7849 14569 7883 14603
rect 12265 14569 12299 14603
rect 21557 14569 21591 14603
rect 21925 14569 21959 14603
rect 2421 14501 2455 14535
rect 4077 14501 4111 14535
rect 5549 14501 5583 14535
rect 6745 14501 6779 14535
rect 18153 14501 18187 14535
rect 23581 14501 23615 14535
rect 2835 14433 2869 14467
rect 4537 14433 4571 14467
rect 5963 14433 5997 14467
rect 11253 14433 11287 14467
rect 14473 14433 14507 14467
rect 14933 14433 14967 14467
rect 15209 14433 15243 14467
rect 15347 14433 15381 14467
rect 16865 14433 16899 14467
rect 17258 14433 17292 14467
rect 18061 14433 18095 14467
rect 22109 14433 22143 14467
rect 22569 14433 22603 14467
rect 24133 14433 24167 14467
rect 1777 14365 1811 14399
rect 1961 14365 1995 14399
rect 2697 14365 2731 14399
rect 2973 14365 3007 14399
rect 3985 14365 4019 14399
rect 4261 14365 4295 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 5825 14365 5859 14399
rect 6101 14365 6135 14399
rect 6837 14365 6871 14399
rect 7111 14365 7145 14399
rect 11527 14365 11561 14399
rect 12633 14365 12667 14399
rect 12875 14365 12909 14399
rect 14289 14365 14323 14399
rect 15485 14365 15519 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 17141 14365 17175 14399
rect 17417 14365 17451 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 18889 14365 18923 14399
rect 21097 14365 21131 14399
rect 21465 14365 21499 14399
rect 21833 14365 21867 14399
rect 22385 14365 22419 14399
rect 22477 14365 22511 14399
rect 22661 14365 22695 14399
rect 23305 14365 23339 14399
rect 23397 14365 23431 14399
rect 23857 14365 23891 14399
rect 16129 14297 16163 14331
rect 3617 14229 3651 14263
rect 3801 14229 3835 14263
rect 13645 14229 13679 14263
rect 18521 14229 18555 14263
rect 18705 14229 18739 14263
rect 20913 14229 20947 14263
rect 22109 14229 22143 14263
rect 22201 14229 22235 14263
rect 23121 14229 23155 14263
rect 1593 14025 1627 14059
rect 3249 14025 3283 14059
rect 5917 14025 5951 14059
rect 14289 14025 14323 14059
rect 15669 14025 15703 14059
rect 17693 14025 17727 14059
rect 23213 14025 23247 14059
rect 1501 13957 1535 13991
rect 22845 13957 22879 13991
rect 23857 13957 23891 13991
rect 2145 13889 2179 13923
rect 2511 13889 2545 13923
rect 3709 13889 3743 13923
rect 4353 13889 4387 13923
rect 5179 13889 5213 13923
rect 6837 13889 6871 13923
rect 7111 13889 7145 13923
rect 8491 13889 8525 13923
rect 9839 13889 9873 13923
rect 12449 13889 12483 13923
rect 13369 13889 13403 13923
rect 13507 13889 13541 13923
rect 14915 13919 14949 13953
rect 16681 13889 16715 13923
rect 16939 13919 16973 13953
rect 18303 13889 18337 13923
rect 19441 13889 19475 13923
rect 19625 13889 19659 13923
rect 22753 13889 22787 13923
rect 22937 13889 22971 13923
rect 23029 13889 23063 13923
rect 23213 13889 23247 13923
rect 23489 13889 23523 13923
rect 24133 13889 24167 13923
rect 2237 13821 2271 13855
rect 4905 13821 4939 13855
rect 8217 13821 8251 13855
rect 9597 13821 9631 13855
rect 12633 13821 12667 13855
rect 13093 13821 13127 13855
rect 13645 13821 13679 13855
rect 14657 13821 14691 13855
rect 18061 13821 18095 13855
rect 19533 13821 19567 13855
rect 23397 13821 23431 13855
rect 4169 13753 4203 13787
rect 19073 13753 19107 13787
rect 23489 13753 23523 13787
rect 1961 13685 1995 13719
rect 3801 13685 3835 13719
rect 7849 13685 7883 13719
rect 9229 13685 9263 13719
rect 10609 13685 10643 13719
rect 24409 13685 24443 13719
rect 2329 13481 2363 13515
rect 2881 13481 2915 13515
rect 13645 13481 13679 13515
rect 16497 13481 16531 13515
rect 18613 13481 18647 13515
rect 18705 13481 18739 13515
rect 22661 13481 22695 13515
rect 1685 13413 1719 13447
rect 9321 13413 9355 13447
rect 22293 13413 22327 13447
rect 3801 13345 3835 13379
rect 9965 13345 9999 13379
rect 10425 13345 10459 13379
rect 10839 13345 10873 13379
rect 15485 13345 15519 13379
rect 18797 13345 18831 13379
rect 20453 13345 20487 13379
rect 22845 13345 22879 13379
rect 1501 13277 1535 13311
rect 3433 13277 3467 13311
rect 4059 13277 4093 13311
rect 9505 13293 9539 13327
rect 9781 13277 9815 13311
rect 10701 13277 10735 13311
rect 10977 13277 11011 13311
rect 12633 13277 12667 13311
rect 12907 13277 12941 13311
rect 15727 13277 15761 13311
rect 18521 13277 18555 13311
rect 19717 13277 19751 13311
rect 19901 13277 19935 13311
rect 20361 13277 20395 13311
rect 20637 13277 20671 13311
rect 20821 13277 20855 13311
rect 22477 13277 22511 13311
rect 22593 13279 22627 13313
rect 2237 13209 2271 13243
rect 2789 13209 2823 13243
rect 20177 13209 20211 13243
rect 20269 13209 20303 13243
rect 20729 13209 20763 13243
rect 23112 13209 23146 13243
rect 3249 13141 3283 13175
rect 4813 13141 4847 13175
rect 11621 13141 11655 13175
rect 24225 13141 24259 13175
rect 9873 12937 9907 12971
rect 11069 12937 11103 12971
rect 21373 12937 21407 12971
rect 22201 12937 22235 12971
rect 23397 12937 23431 12971
rect 1501 12869 1535 12903
rect 1869 12869 1903 12903
rect 23949 12869 23983 12903
rect 2329 12801 2363 12835
rect 2603 12801 2637 12835
rect 3709 12801 3743 12835
rect 4746 12801 4780 12835
rect 4905 12801 4939 12835
rect 6619 12801 6653 12835
rect 8033 12801 8067 12835
rect 8217 12801 8251 12835
rect 9070 12801 9104 12835
rect 9229 12801 9263 12835
rect 10331 12801 10365 12835
rect 11987 12801 12021 12835
rect 14179 12831 14213 12865
rect 17031 12831 17065 12865
rect 18245 12801 18279 12835
rect 18519 12801 18553 12835
rect 19625 12801 19659 12835
rect 19892 12801 19926 12835
rect 21281 12801 21315 12835
rect 21557 12801 21591 12835
rect 22109 12801 22143 12835
rect 22643 12831 22677 12865
rect 3893 12733 3927 12767
rect 4353 12733 4387 12767
rect 4629 12733 4663 12767
rect 6377 12733 6411 12767
rect 8953 12733 8987 12767
rect 10057 12733 10091 12767
rect 11713 12733 11747 12767
rect 13921 12733 13955 12767
rect 16773 12733 16807 12767
rect 22385 12733 22419 12767
rect 7389 12665 7423 12699
rect 8677 12665 8711 12699
rect 19257 12665 19291 12699
rect 21005 12665 21039 12699
rect 3341 12597 3375 12631
rect 5549 12597 5583 12631
rect 12725 12597 12759 12631
rect 14933 12597 14967 12631
rect 17785 12597 17819 12631
rect 21097 12597 21131 12631
rect 24225 12597 24259 12631
rect 3985 12393 4019 12427
rect 22661 12393 22695 12427
rect 24133 12393 24167 12427
rect 5549 12325 5583 12359
rect 7481 12325 7515 12359
rect 15577 12325 15611 12359
rect 23305 12325 23339 12359
rect 23765 12325 23799 12359
rect 1777 12257 1811 12291
rect 1961 12257 1995 12291
rect 2421 12257 2455 12291
rect 2697 12257 2731 12291
rect 2835 12257 2869 12291
rect 2973 12257 3007 12291
rect 5825 12257 5859 12291
rect 6101 12257 6135 12291
rect 6837 12257 6871 12291
rect 7874 12257 7908 12291
rect 17049 12257 17083 12291
rect 17442 12257 17476 12291
rect 17601 12257 17635 12291
rect 3893 12189 3927 12223
rect 4445 12189 4479 12223
rect 4905 12189 4939 12223
rect 5089 12189 5123 12223
rect 5963 12189 5997 12223
rect 7021 12189 7055 12223
rect 7757 12189 7791 12223
rect 8033 12189 8067 12223
rect 11897 12189 11931 12223
rect 14657 12189 14691 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 17325 12189 17359 12223
rect 19901 12189 19935 12223
rect 20143 12189 20177 12223
rect 21281 12189 21315 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 23949 12189 23983 12223
rect 11805 12121 11839 12155
rect 12265 12121 12299 12155
rect 14565 12121 14599 12155
rect 15025 12121 15059 12155
rect 21548 12121 21582 12155
rect 3617 12053 3651 12087
rect 4537 12053 4571 12087
rect 6745 12053 6779 12087
rect 8677 12053 8711 12087
rect 11529 12053 11563 12087
rect 12633 12053 12667 12087
rect 12817 12053 12851 12087
rect 14289 12053 14323 12087
rect 15393 12053 15427 12087
rect 18245 12053 18279 12087
rect 20913 12053 20947 12087
rect 22845 12053 22879 12087
rect 23121 12053 23155 12087
rect 2881 11849 2915 11883
rect 4537 11849 4571 11883
rect 5917 11849 5951 11883
rect 7941 11849 7975 11883
rect 12541 11849 12575 11883
rect 13921 11849 13955 11883
rect 17693 11849 17727 11883
rect 21465 11849 21499 11883
rect 23397 11849 23431 11883
rect 2143 11713 2177 11747
rect 3433 11737 3467 11771
rect 3525 11713 3559 11747
rect 3799 11713 3833 11747
rect 5179 11713 5213 11747
rect 6929 11713 6963 11747
rect 7187 11743 7221 11777
rect 8309 11713 8343 11747
rect 8583 11713 8617 11747
rect 11529 11713 11563 11747
rect 11803 11713 11837 11747
rect 12909 11713 12943 11747
rect 13183 11713 13217 11747
rect 14933 11713 14967 11747
rect 15207 11713 15241 11747
rect 16923 11713 16957 11747
rect 18303 11713 18337 11747
rect 21649 11713 21683 11747
rect 22385 11713 22419 11747
rect 22753 11713 22787 11747
rect 23305 11713 23339 11747
rect 23581 11713 23615 11747
rect 23673 11713 23707 11747
rect 24133 11713 24167 11747
rect 1869 11645 1903 11679
rect 4905 11645 4939 11679
rect 16681 11645 16715 11679
rect 18061 11645 18095 11679
rect 21925 11645 21959 11679
rect 22661 11577 22695 11611
rect 23121 11577 23155 11611
rect 3249 11509 3283 11543
rect 9321 11509 9355 11543
rect 15945 11509 15979 11543
rect 19073 11509 19107 11543
rect 23857 11509 23891 11543
rect 24409 11509 24443 11543
rect 1777 11305 1811 11339
rect 2329 11305 2363 11339
rect 4537 11305 4571 11339
rect 5089 11305 5123 11339
rect 7665 11305 7699 11339
rect 18153 11305 18187 11339
rect 23765 11305 23799 11339
rect 5457 11237 5491 11271
rect 15853 11237 15887 11271
rect 17049 11237 17083 11271
rect 18705 11237 18739 11271
rect 8953 11169 8987 11203
rect 9590 11169 9624 11203
rect 9873 11169 9907 11203
rect 16129 11169 16163 11203
rect 16246 11169 16280 11203
rect 16405 11169 16439 11203
rect 18889 11169 18923 11203
rect 3617 11101 3651 11135
rect 4997 11101 5031 11135
rect 5641 11101 5675 11135
rect 6653 11101 6687 11135
rect 6927 11101 6961 11135
rect 9137 11101 9171 11135
rect 9990 11101 10024 11135
rect 10149 11101 10183 11135
rect 15209 11101 15243 11135
rect 15393 11101 15427 11135
rect 17141 11101 17175 11135
rect 17415 11101 17449 11135
rect 18705 11101 18739 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 20085 11101 20119 11135
rect 20269 11101 20303 11135
rect 20729 11101 20763 11135
rect 22753 11101 22787 11135
rect 23027 11101 23061 11135
rect 1685 11033 1719 11067
rect 2237 11033 2271 11067
rect 2973 11033 3007 11067
rect 3893 11033 3927 11067
rect 4445 11033 4479 11067
rect 10793 11033 10827 11067
rect 19073 11033 19107 11067
rect 19349 11033 19383 11067
rect 21005 11033 21039 11067
rect 3065 10965 3099 10999
rect 3433 10965 3467 10999
rect 3985 10965 4019 10999
rect 1593 10761 1627 10795
rect 3801 10761 3835 10795
rect 10241 10761 10275 10795
rect 10977 10761 11011 10795
rect 14933 10761 14967 10795
rect 20269 10761 20303 10795
rect 20729 10761 20763 10795
rect 20913 10761 20947 10795
rect 1501 10693 1535 10727
rect 13645 10693 13679 10727
rect 14749 10693 14783 10727
rect 2145 10625 2179 10659
rect 2511 10635 2545 10669
rect 3985 10625 4019 10659
rect 4351 10625 4385 10659
rect 6377 10625 6411 10659
rect 6651 10625 6685 10659
rect 9229 10625 9263 10659
rect 9503 10625 9537 10659
rect 10793 10625 10827 10659
rect 12323 10625 12357 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 14381 10625 14415 10659
rect 17693 10625 17727 10659
rect 17785 10625 17819 10659
rect 18052 10625 18086 10659
rect 19257 10625 19291 10659
rect 19531 10625 19565 10659
rect 20637 10625 20671 10659
rect 20821 10625 20855 10659
rect 21097 10625 21131 10659
rect 22661 10625 22695 10659
rect 22995 10625 23029 10659
rect 2237 10557 2271 10591
rect 4077 10557 4111 10591
rect 12081 10557 12115 10591
rect 22753 10557 22787 10591
rect 3249 10489 3283 10523
rect 13093 10489 13127 10523
rect 1961 10421 1995 10455
rect 5089 10421 5123 10455
rect 7389 10421 7423 10455
rect 17509 10421 17543 10455
rect 19165 10421 19199 10455
rect 22477 10421 22511 10455
rect 23765 10421 23799 10455
rect 7573 10217 7607 10251
rect 15117 10217 15151 10251
rect 18429 10217 18463 10251
rect 20177 10217 20211 10251
rect 10977 10149 11011 10183
rect 20361 10149 20395 10183
rect 1777 10081 1811 10115
rect 1961 10081 1995 10115
rect 2421 10081 2455 10115
rect 2697 10081 2731 10115
rect 2973 10081 3007 10115
rect 4445 10081 4479 10115
rect 4721 10081 4755 10115
rect 4859 10081 4893 10115
rect 4997 10081 5031 10115
rect 5917 10081 5951 10115
rect 6377 10081 6411 10115
rect 6653 10081 6687 10115
rect 6770 10081 6804 10115
rect 6929 10081 6963 10115
rect 9965 10081 9999 10115
rect 20821 10081 20855 10115
rect 1685 10013 1719 10047
rect 2835 10013 2869 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 5733 10013 5767 10047
rect 10223 9983 10257 10017
rect 11897 10013 11931 10047
rect 14105 10013 14139 10047
rect 14379 10013 14413 10047
rect 18337 10013 18371 10047
rect 19073 10013 19107 10047
rect 20085 10013 20119 10047
rect 20545 10013 20579 10047
rect 21095 10013 21129 10047
rect 22477 10013 22511 10047
rect 22753 10013 22787 10047
rect 22995 10013 23029 10047
rect 11805 9945 11839 9979
rect 12265 9945 12299 9979
rect 1501 9877 1535 9911
rect 3617 9877 3651 9911
rect 5641 9877 5675 9911
rect 11529 9877 11563 9911
rect 12633 9877 12667 9911
rect 12817 9877 12851 9911
rect 18889 9877 18923 9911
rect 21833 9877 21867 9911
rect 22293 9877 22327 9911
rect 23765 9877 23799 9911
rect 2697 9673 2731 9707
rect 4537 9673 4571 9707
rect 5917 9673 5951 9707
rect 11253 9673 11287 9707
rect 12817 9673 12851 9707
rect 21097 9673 21131 9707
rect 19984 9605 20018 9639
rect 1593 9561 1627 9595
rect 1685 9537 1719 9571
rect 1959 9537 1993 9571
rect 3249 9537 3283 9571
rect 3767 9537 3801 9571
rect 5147 9537 5181 9571
rect 7481 9537 7515 9571
rect 8401 9537 8435 9571
rect 8677 9537 8711 9571
rect 9597 9537 9631 9571
rect 10450 9537 10484 9571
rect 10609 9537 10643 9571
rect 12079 9537 12113 9571
rect 18337 9537 18371 9571
rect 18595 9567 18629 9601
rect 21833 9537 21867 9571
rect 22109 9537 22143 9571
rect 22293 9537 22327 9571
rect 22569 9537 22603 9571
rect 22995 9537 23029 9571
rect 24317 9537 24351 9571
rect 3525 9469 3559 9503
rect 4905 9469 4939 9503
rect 7665 9469 7699 9503
rect 8125 9469 8159 9503
rect 8539 9469 8573 9503
rect 9413 9469 9447 9503
rect 10333 9469 10367 9503
rect 11805 9469 11839 9503
rect 19717 9469 19751 9503
rect 22753 9469 22787 9503
rect 9321 9401 9355 9435
rect 10057 9401 10091 9435
rect 22385 9401 22419 9435
rect 23765 9401 23799 9435
rect 1409 9333 1443 9367
rect 3065 9333 3099 9367
rect 19349 9333 19383 9367
rect 21925 9333 21959 9367
rect 22201 9333 22235 9367
rect 24133 9333 24167 9367
rect 2697 9129 2731 9163
rect 4077 9129 4111 9163
rect 8493 9129 8527 9163
rect 10793 9129 10827 9163
rect 22661 9129 22695 9163
rect 23397 9129 23431 9163
rect 23949 9129 23983 9163
rect 2237 9061 2271 9095
rect 9781 8993 9815 9027
rect 14105 8993 14139 9027
rect 15485 8993 15519 9027
rect 16865 8993 16899 9027
rect 1501 8925 1535 8959
rect 2053 8925 2087 8959
rect 3157 8925 3191 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 7481 8925 7515 8959
rect 7755 8925 7789 8959
rect 10055 8925 10089 8959
rect 14347 8925 14381 8959
rect 15759 8925 15793 8959
rect 17107 8925 17141 8959
rect 21281 8925 21315 8959
rect 22937 8925 22971 8959
rect 23673 8925 23707 8959
rect 2605 8857 2639 8891
rect 21548 8857 21582 8891
rect 23121 8857 23155 8891
rect 1593 8789 1627 8823
rect 3249 8789 3283 8823
rect 3801 8789 3835 8823
rect 15117 8789 15151 8823
rect 16497 8789 16531 8823
rect 17877 8789 17911 8823
rect 22753 8789 22787 8823
rect 1593 8585 1627 8619
rect 7113 8585 7147 8619
rect 8401 8585 8435 8619
rect 10149 8585 10183 8619
rect 13001 8585 13035 8619
rect 17141 8585 17175 8619
rect 19625 8585 19659 8619
rect 1501 8517 1535 8551
rect 2605 8517 2639 8551
rect 11713 8517 11747 8551
rect 11989 8517 12023 8551
rect 12449 8517 12483 8551
rect 12817 8517 12851 8551
rect 13829 8517 13863 8551
rect 14197 8517 14231 8551
rect 14933 8517 14967 8551
rect 17417 8517 17451 8551
rect 17509 8517 17543 8551
rect 22937 8517 22971 8551
rect 2053 8449 2087 8483
rect 2421 8449 2455 8483
rect 3157 8449 3191 8483
rect 3709 8449 3743 8483
rect 7297 8449 7331 8483
rect 7663 8449 7697 8483
rect 9379 8449 9413 8483
rect 12081 8449 12115 8483
rect 14105 8449 14139 8483
rect 14565 8449 14599 8483
rect 17877 8449 17911 8483
rect 18259 8449 18293 8483
rect 18613 8449 18647 8483
rect 18887 8449 18921 8483
rect 19993 8449 20027 8483
rect 20177 8449 20211 8483
rect 21833 8449 21867 8483
rect 22201 8449 22235 8483
rect 22661 8449 22695 8483
rect 23489 8449 23523 8483
rect 24041 8449 24075 8483
rect 24501 8449 24535 8483
rect 7389 8381 7423 8415
rect 9137 8381 9171 8415
rect 23305 8381 23339 8415
rect 2789 8313 2823 8347
rect 3341 8313 3375 8347
rect 3893 8313 3927 8347
rect 15117 8313 15151 8347
rect 23949 8313 23983 8347
rect 18429 8245 18463 8279
rect 20085 8245 20119 8279
rect 24317 8245 24351 8279
rect 1777 8041 1811 8075
rect 3341 8041 3375 8075
rect 8125 8041 8159 8075
rect 10885 8041 10919 8075
rect 12265 8041 12299 8075
rect 13645 8041 13679 8075
rect 19901 8041 19935 8075
rect 22661 8041 22695 8075
rect 5917 7973 5951 8007
rect 6929 7973 6963 8007
rect 15945 7973 15979 8007
rect 19441 7973 19475 8007
rect 6285 7905 6319 7939
rect 6469 7905 6503 7939
rect 7205 7905 7239 7939
rect 7343 7905 7377 7939
rect 9873 7905 9907 7939
rect 11253 7905 11287 7939
rect 12633 7905 12667 7939
rect 15485 7905 15519 7939
rect 16338 7905 16372 7939
rect 16497 7905 16531 7939
rect 18889 7905 18923 7939
rect 21189 7905 21223 7939
rect 22845 7905 22879 7939
rect 1501 7837 1535 7871
rect 1961 7837 1995 7871
rect 2235 7837 2269 7871
rect 3525 7837 3559 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 4905 7837 4939 7871
rect 5179 7837 5213 7871
rect 7481 7837 7515 7871
rect 10147 7837 10181 7871
rect 11527 7837 11561 7871
rect 12891 7807 12925 7841
rect 15301 7837 15335 7871
rect 16221 7837 16255 7871
rect 17233 7837 17267 7871
rect 17507 7837 17541 7871
rect 18797 7837 18831 7871
rect 19441 7837 19475 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 20361 7837 20395 7871
rect 20637 7837 20671 7871
rect 21097 7837 21131 7871
rect 22477 7837 22511 7871
rect 22569 7837 22603 7871
rect 19809 7769 19843 7803
rect 23112 7769 23146 7803
rect 2973 7701 3007 7735
rect 3801 7701 3835 7735
rect 4077 7701 4111 7735
rect 17141 7701 17175 7735
rect 18245 7701 18279 7735
rect 22293 7701 22327 7735
rect 24225 7701 24259 7735
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 4261 7497 4295 7531
rect 7481 7497 7515 7531
rect 14381 7497 14415 7531
rect 14565 7497 14599 7531
rect 19533 7497 19567 7531
rect 19993 7497 20027 7531
rect 21557 7497 21591 7531
rect 23305 7497 23339 7531
rect 13277 7429 13311 7463
rect 13553 7429 13587 7463
rect 23857 7429 23891 7463
rect 1501 7361 1535 7395
rect 2329 7361 2363 7395
rect 3458 7361 3492 7395
rect 3617 7361 3651 7395
rect 5273 7361 5307 7395
rect 6469 7361 6503 7395
rect 6727 7391 6761 7425
rect 8291 7391 8325 7425
rect 9687 7371 9721 7405
rect 13645 7361 13679 7395
rect 14013 7361 14047 7395
rect 18153 7361 18187 7395
rect 18420 7361 18454 7395
rect 19901 7361 19935 7395
rect 20444 7361 20478 7395
rect 22017 7361 22051 7395
rect 22551 7391 22585 7425
rect 24501 7361 24535 7395
rect 2421 7293 2455 7327
rect 2605 7293 2639 7327
rect 3065 7293 3099 7327
rect 3341 7293 3375 7327
rect 4353 7293 4387 7327
rect 4537 7293 4571 7327
rect 5390 7293 5424 7327
rect 5549 7293 5583 7327
rect 8033 7293 8067 7327
rect 9413 7293 9447 7327
rect 20177 7293 20211 7327
rect 22293 7293 22327 7327
rect 24133 7293 24167 7327
rect 4997 7225 5031 7259
rect 6193 7225 6227 7259
rect 24317 7225 24351 7259
rect 9045 7157 9079 7191
rect 10425 7157 10459 7191
rect 21833 7157 21867 7191
rect 3341 6953 3375 6987
rect 5549 6953 5583 6987
rect 13553 6953 13587 6987
rect 18613 6953 18647 6987
rect 20361 6953 20395 6987
rect 20729 6953 20763 6987
rect 21097 6953 21131 6987
rect 21281 6953 21315 6987
rect 9597 6885 9631 6919
rect 22661 6885 22695 6919
rect 1961 6817 1995 6851
rect 2329 6817 2363 6851
rect 4537 6817 4571 6851
rect 8953 6817 8987 6851
rect 9137 6817 9171 6851
rect 9873 6817 9907 6851
rect 10149 6817 10183 6851
rect 12541 6817 12575 6851
rect 22017 6817 22051 6851
rect 24041 6817 24075 6851
rect 1685 6749 1719 6783
rect 2587 6719 2621 6753
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 4811 6749 4845 6783
rect 10011 6749 10045 6783
rect 12815 6749 12849 6783
rect 18797 6749 18831 6783
rect 19349 6749 19383 6783
rect 19623 6749 19657 6783
rect 20913 6749 20947 6783
rect 21005 6749 21039 6783
rect 21189 6749 21223 6783
rect 21465 6749 21499 6783
rect 21557 6749 21591 6783
rect 22201 6749 22235 6783
rect 22753 6749 22787 6783
rect 23397 6749 23431 6783
rect 23489 6749 23523 6783
rect 23949 6749 23983 6783
rect 24133 6749 24167 6783
rect 3801 6613 3835 6647
rect 4077 6613 4111 6647
rect 10793 6613 10827 6647
rect 21741 6613 21775 6647
rect 23213 6613 23247 6647
rect 23581 6613 23615 6647
rect 3433 6409 3467 6443
rect 4997 6409 5031 6443
rect 8309 6409 8343 6443
rect 14473 6409 14507 6443
rect 17969 6409 18003 6443
rect 20637 6409 20671 6443
rect 23305 6409 23339 6443
rect 23949 6409 23983 6443
rect 24317 6409 24351 6443
rect 2605 6341 2639 6375
rect 3341 6341 3375 6375
rect 21281 6341 21315 6375
rect 1501 6273 1535 6307
rect 2237 6273 2271 6307
rect 2789 6273 2823 6307
rect 3985 6273 4019 6307
rect 4259 6273 4293 6307
rect 5549 6273 5583 6307
rect 5825 6273 5859 6307
rect 6101 6273 6135 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7297 6273 7331 6307
rect 7414 6273 7448 6307
rect 7573 6273 7607 6307
rect 8217 6273 8251 6307
rect 8493 6273 8527 6307
rect 9045 6273 9079 6307
rect 9781 6273 9815 6307
rect 9898 6273 9932 6307
rect 11529 6273 11563 6307
rect 12587 6273 12621 6307
rect 12725 6273 12759 6307
rect 13703 6273 13737 6307
rect 15207 6273 15241 6307
rect 17693 6273 17727 6307
rect 20545 6273 20579 6307
rect 20821 6273 20855 6307
rect 21097 6273 21131 6307
rect 21189 6273 21223 6307
rect 21649 6273 21683 6307
rect 22107 6273 22141 6307
rect 23213 6273 23247 6307
rect 23397 6273 23431 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 24041 6273 24075 6307
rect 24501 6273 24535 6307
rect 8861 6205 8895 6239
rect 10057 6205 10091 6239
rect 11713 6205 11747 6239
rect 12449 6205 12483 6239
rect 13461 6205 13495 6239
rect 14933 6205 14967 6239
rect 17969 6205 18003 6239
rect 21833 6205 21867 6239
rect 5641 6137 5675 6171
rect 7021 6137 7055 6171
rect 9505 6137 9539 6171
rect 12173 6137 12207 6171
rect 17785 6137 17819 6171
rect 20361 6137 20395 6171
rect 21465 6137 21499 6171
rect 22845 6137 22879 6171
rect 24225 6137 24259 6171
rect 1593 6069 1627 6103
rect 2881 6069 2915 6103
rect 5365 6069 5399 6103
rect 5917 6069 5951 6103
rect 10701 6069 10735 6103
rect 13369 6069 13403 6103
rect 15945 6069 15979 6103
rect 20913 6069 20947 6103
rect 23581 6069 23615 6103
rect 1777 5865 1811 5899
rect 2145 5865 2179 5899
rect 3249 5865 3283 5899
rect 5549 5865 5583 5899
rect 7113 5865 7147 5899
rect 8493 5865 8527 5899
rect 10885 5865 10919 5899
rect 12265 5865 12299 5899
rect 18245 5865 18279 5899
rect 21189 5865 21223 5899
rect 21465 5865 21499 5899
rect 22937 5865 22971 5899
rect 15945 5797 15979 5831
rect 6101 5729 6135 5763
rect 7481 5729 7515 5763
rect 16338 5729 16372 5763
rect 16497 5729 16531 5763
rect 19257 5729 19291 5763
rect 1685 5661 1719 5695
rect 2329 5661 2363 5695
rect 3157 5661 3191 5695
rect 3985 5661 4019 5695
rect 4259 5661 4293 5695
rect 6359 5631 6393 5665
rect 7755 5661 7789 5695
rect 9873 5661 9907 5695
rect 10147 5661 10181 5695
rect 11253 5661 11287 5695
rect 11527 5661 11561 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 16221 5661 16255 5695
rect 17233 5661 17267 5695
rect 17507 5661 17541 5695
rect 19499 5661 19533 5695
rect 20913 5661 20947 5695
rect 21005 5661 21039 5695
rect 21281 5661 21315 5695
rect 21557 5661 21591 5695
rect 23305 5661 23339 5695
rect 23581 5661 23615 5695
rect 23949 5661 23983 5695
rect 2605 5593 2639 5627
rect 5457 5593 5491 5627
rect 21824 5593 21858 5627
rect 24225 5593 24259 5627
rect 2881 5525 2915 5559
rect 4997 5525 5031 5559
rect 17141 5525 17175 5559
rect 20269 5525 20303 5559
rect 20729 5525 20763 5559
rect 6193 5321 6227 5355
rect 7389 5321 7423 5355
rect 10241 5321 10275 5355
rect 16497 5321 16531 5355
rect 17693 5321 17727 5355
rect 18153 5321 18187 5355
rect 18429 5321 18463 5355
rect 22017 5321 22051 5355
rect 24501 5321 24535 5355
rect 1409 5185 1443 5219
rect 1683 5185 1717 5219
rect 2789 5185 2823 5219
rect 3063 5185 3097 5219
rect 4353 5185 4387 5219
rect 5273 5185 5307 5219
rect 5549 5185 5583 5219
rect 6377 5185 6411 5219
rect 6651 5185 6685 5219
rect 9487 5215 9521 5249
rect 12725 5185 12759 5219
rect 14657 5185 14691 5219
rect 16681 5185 16715 5219
rect 16955 5185 16989 5219
rect 18061 5185 18095 5219
rect 18337 5185 18371 5219
rect 18521 5185 18555 5219
rect 18797 5185 18831 5219
rect 19165 5185 19199 5219
rect 19349 5185 19383 5219
rect 19515 5185 19549 5219
rect 19867 5185 19901 5219
rect 21189 5185 21223 5219
rect 21557 5185 21591 5219
rect 21833 5185 21867 5219
rect 22109 5185 22143 5219
rect 22569 5185 22603 5219
rect 22661 5185 22695 5219
rect 23377 5185 23411 5219
rect 4537 5117 4571 5151
rect 4997 5117 5031 5151
rect 5390 5117 5424 5151
rect 9229 5117 9263 5151
rect 12909 5117 12943 5151
rect 13645 5117 13679 5151
rect 13783 5117 13817 5151
rect 13921 5117 13955 5151
rect 14841 5117 14875 5151
rect 15577 5117 15611 5151
rect 15715 5117 15749 5151
rect 15853 5117 15887 5151
rect 19625 5117 19659 5151
rect 21005 5117 21039 5151
rect 23121 5117 23155 5151
rect 13369 5049 13403 5083
rect 15301 5049 15335 5083
rect 18613 5049 18647 5083
rect 19165 5049 19199 5083
rect 20637 5049 20671 5083
rect 21189 5049 21223 5083
rect 22293 5049 22327 5083
rect 2421 4981 2455 5015
rect 3801 4981 3835 5015
rect 14565 4981 14599 5015
rect 22385 4981 22419 5015
rect 22753 4981 22787 5015
rect 1501 4777 1535 4811
rect 5549 4777 5583 4811
rect 13645 4777 13679 4811
rect 16405 4777 16439 4811
rect 18797 4777 18831 4811
rect 19349 4777 19383 4811
rect 19625 4777 19659 4811
rect 20361 4777 20395 4811
rect 21005 4777 21039 4811
rect 21281 4777 21315 4811
rect 22201 4777 22235 4811
rect 24041 4777 24075 4811
rect 3801 4709 3835 4743
rect 18889 4709 18923 4743
rect 1961 4641 1995 4675
rect 2421 4641 2455 4675
rect 2697 4641 2731 4675
rect 2835 4641 2869 4675
rect 22477 4641 22511 4675
rect 1685 4573 1719 4607
rect 1777 4573 1811 4607
rect 2973 4573 3007 4607
rect 3985 4573 4019 4607
rect 4261 4573 4295 4607
rect 4537 4573 4571 4607
rect 4811 4573 4845 4607
rect 12633 4573 12667 4607
rect 12907 4573 12941 4607
rect 15393 4573 15427 4607
rect 15667 4573 15701 4607
rect 17417 4573 17451 4607
rect 19073 4573 19107 4607
rect 19257 4573 19291 4607
rect 19533 4573 19567 4607
rect 19717 4573 19751 4607
rect 19993 4573 20027 4607
rect 20085 4573 20119 4607
rect 20269 4573 20303 4607
rect 20545 4573 20579 4607
rect 20821 4573 20855 4607
rect 20913 4573 20947 4607
rect 21189 4573 21223 4607
rect 21373 4573 21407 4607
rect 21649 4573 21683 4607
rect 21925 4573 21959 4607
rect 22017 4573 22051 4607
rect 22719 4573 22753 4607
rect 17684 4505 17718 4539
rect 23949 4505 23983 4539
rect 3617 4437 3651 4471
rect 4077 4437 4111 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 20637 4437 20671 4471
rect 21465 4437 21499 4471
rect 21741 4437 21775 4471
rect 23489 4437 23523 4471
rect 4353 4233 4387 4267
rect 15577 4233 15611 4267
rect 17693 4233 17727 4267
rect 18337 4233 18371 4267
rect 19165 4233 19199 4267
rect 21465 4233 21499 4267
rect 1501 4165 1535 4199
rect 19625 4165 19659 4199
rect 24317 4165 24351 4199
rect 2305 4097 2339 4131
rect 2421 4097 2455 4131
rect 2605 4097 2639 4131
rect 3341 4097 3375 4131
rect 3479 4097 3513 4131
rect 3617 4097 3651 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 6745 4097 6779 4131
rect 7019 4097 7053 4131
rect 9321 4097 9355 4131
rect 10331 4097 10365 4131
rect 11529 4097 11563 4131
rect 11803 4097 11837 4131
rect 14565 4097 14599 4131
rect 14839 4097 14873 4131
rect 17877 4097 17911 4131
rect 18521 4097 18555 4131
rect 18797 4097 18831 4131
rect 19073 4097 19107 4131
rect 19349 4097 19383 4131
rect 20352 4097 20386 4131
rect 22385 4097 22419 4131
rect 22661 4097 22695 4131
rect 23029 4097 23063 4131
rect 24501 4097 24535 4131
rect 8125 4029 8159 4063
rect 8309 4029 8343 4063
rect 9045 4029 9079 4063
rect 9183 4029 9217 4063
rect 10057 4029 10091 4063
rect 20085 4029 20119 4063
rect 22017 4029 22051 4063
rect 23857 4029 23891 4063
rect 1685 3961 1719 3995
rect 3065 3961 3099 3995
rect 7757 3961 7791 3995
rect 8769 3961 8803 3995
rect 22661 3961 22695 3995
rect 2145 3893 2179 3927
rect 9965 3893 9999 3927
rect 11069 3893 11103 3927
rect 12541 3893 12575 3927
rect 18613 3893 18647 3927
rect 18889 3893 18923 3927
rect 19717 3893 19751 3927
rect 1777 3689 1811 3723
rect 13369 3689 13403 3723
rect 15117 3689 15151 3723
rect 20637 3689 20671 3723
rect 23949 3689 23983 3723
rect 2421 3621 2455 3655
rect 2881 3621 2915 3655
rect 7205 3621 7239 3655
rect 8493 3621 8527 3655
rect 18521 3621 18555 3655
rect 7481 3553 7515 3587
rect 9597 3553 9631 3587
rect 9873 3553 9907 3587
rect 9990 3553 10024 3587
rect 19257 3553 19291 3587
rect 21281 3553 21315 3587
rect 23213 3553 23247 3587
rect 1685 3485 1719 3519
rect 2697 3485 2731 3519
rect 4813 3485 4847 3519
rect 5089 3485 5123 3519
rect 5363 3485 5397 3519
rect 7389 3485 7423 3519
rect 7755 3485 7789 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 10149 3485 10183 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 14379 3485 14413 3519
rect 17969 3461 18003 3495
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 18797 3485 18831 3519
rect 19073 3485 19107 3519
rect 20821 3485 20855 3519
rect 21555 3485 21589 3519
rect 22661 3485 22695 3519
rect 23765 3485 23799 3519
rect 2237 3417 2271 3451
rect 6929 3417 6963 3451
rect 12081 3417 12115 3451
rect 12357 3417 12391 3451
rect 12449 3417 12483 3451
rect 12817 3417 12851 3451
rect 19524 3417 19558 3451
rect 4905 3349 4939 3383
rect 6101 3349 6135 3383
rect 10793 3349 10827 3383
rect 13185 3349 13219 3383
rect 13553 3349 13587 3383
rect 17785 3349 17819 3383
rect 18245 3349 18279 3383
rect 18613 3349 18647 3383
rect 18889 3349 18923 3383
rect 20913 3349 20947 3383
rect 22293 3349 22327 3383
rect 1593 3145 1627 3179
rect 2605 3145 2639 3179
rect 3341 3145 3375 3179
rect 4537 3145 4571 3179
rect 7849 3145 7883 3179
rect 9137 3145 9171 3179
rect 9965 3145 9999 3179
rect 13185 3145 13219 3179
rect 17141 3145 17175 3179
rect 18061 3145 18095 3179
rect 18797 3145 18831 3179
rect 23397 3145 23431 3179
rect 6561 3077 6595 3111
rect 7665 3077 7699 3111
rect 10241 3077 10275 3111
rect 10333 3077 10367 3111
rect 11069 3077 11103 3111
rect 24317 3077 24351 3111
rect 1501 3009 1535 3043
rect 2053 3009 2087 3043
rect 2237 3009 2271 3043
rect 2513 3009 2547 3043
rect 2789 3009 2823 3043
rect 3249 3009 3283 3043
rect 4445 3009 4479 3043
rect 6837 3009 6871 3043
rect 6929 3009 6963 3043
rect 7297 3009 7331 3043
rect 8125 3009 8159 3043
rect 8399 3009 8433 3043
rect 9689 3009 9723 3043
rect 10701 3009 10735 3043
rect 11713 3009 11747 3043
rect 12081 3009 12115 3043
rect 12447 3009 12481 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17509 3009 17543 3043
rect 17969 3009 18003 3043
rect 18245 3009 18279 3043
rect 18521 3033 18555 3067
rect 18705 3009 18739 3043
rect 19257 3009 19291 3043
rect 19717 3009 19751 3043
rect 20821 3009 20855 3043
rect 21925 3009 21959 3043
rect 22385 3009 22419 3043
rect 22659 3009 22693 3043
rect 23765 3009 23799 3043
rect 23949 3009 23983 3043
rect 12173 2941 12207 2975
rect 19993 2941 20027 2975
rect 21465 2941 21499 2975
rect 11253 2873 11287 2907
rect 17693 2873 17727 2907
rect 17785 2873 17819 2907
rect 23949 2873 23983 2907
rect 2329 2805 2363 2839
rect 9505 2805 9539 2839
rect 11529 2805 11563 2839
rect 11897 2805 11931 2839
rect 17417 2805 17451 2839
rect 18337 2805 18371 2839
rect 19349 2805 19383 2839
rect 22017 2805 22051 2839
rect 1961 2601 1995 2635
rect 3249 2601 3283 2635
rect 4629 2601 4663 2635
rect 6837 2601 6871 2635
rect 9505 2601 9539 2635
rect 10885 2601 10919 2635
rect 17693 2601 17727 2635
rect 24225 2601 24259 2635
rect 1685 2533 1719 2567
rect 3985 2533 4019 2567
rect 11897 2533 11931 2567
rect 16773 2533 16807 2567
rect 2237 2465 2271 2499
rect 19809 2465 19843 2499
rect 1777 2397 1811 2431
rect 2511 2397 2545 2431
rect 3801 2397 3835 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 5733 2397 5767 2431
rect 5825 2397 5859 2431
rect 6099 2397 6133 2431
rect 7389 2397 7423 2431
rect 7665 2397 7699 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 8769 2397 8803 2431
rect 9137 2397 9171 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 10115 2397 10149 2431
rect 11529 2397 11563 2431
rect 11805 2397 11839 2431
rect 12081 2397 12115 2431
rect 12357 2397 12391 2431
rect 12633 2397 12667 2431
rect 12909 2397 12943 2431
rect 13277 2397 13311 2431
rect 14841 2397 14875 2431
rect 15117 2397 15151 2431
rect 15393 2397 15427 2431
rect 15669 2397 15703 2431
rect 16405 2397 16439 2431
rect 16681 2397 16715 2431
rect 16957 2397 16991 2431
rect 17233 2397 17267 2431
rect 18153 2397 18187 2431
rect 18705 2397 18739 2431
rect 19441 2397 19475 2431
rect 19533 2397 19567 2431
rect 20637 2397 20671 2431
rect 21281 2397 21315 2431
rect 21557 2397 21591 2431
rect 22845 2397 22879 2431
rect 23101 2397 23135 2431
rect 1501 2329 1535 2363
rect 17601 2329 17635 2363
rect 22385 2329 22419 2363
rect 4721 2261 4755 2295
rect 5549 2261 5583 2295
rect 7205 2261 7239 2295
rect 7481 2261 7515 2295
rect 7757 2261 7791 2295
rect 8033 2261 8067 2295
rect 8309 2261 8343 2295
rect 8585 2261 8619 2295
rect 8953 2261 8987 2295
rect 11345 2261 11379 2295
rect 11621 2261 11655 2295
rect 12173 2261 12207 2295
rect 12449 2261 12483 2295
rect 12725 2261 12759 2295
rect 13093 2261 13127 2295
rect 14657 2261 14691 2295
rect 14933 2261 14967 2295
rect 15209 2261 15243 2295
rect 15485 2261 15519 2295
rect 16221 2261 16255 2295
rect 16497 2261 16531 2295
rect 17049 2261 17083 2295
rect 18245 2261 18279 2295
rect 18797 2261 18831 2295
rect 19257 2261 19291 2295
rect 2697 2057 2731 2091
rect 3525 2057 3559 2091
rect 4537 2057 4571 2091
rect 5089 2057 5123 2091
rect 6561 2057 6595 2091
rect 7665 2057 7699 2091
rect 8033 2057 8067 2091
rect 8401 2057 8435 2091
rect 8769 2057 8803 2091
rect 9965 2057 9999 2091
rect 15209 2057 15243 2091
rect 18337 2057 18371 2091
rect 23213 2057 23247 2091
rect 3893 1989 3927 2023
rect 6009 1989 6043 2023
rect 6193 1989 6227 2023
rect 6469 1989 6503 2023
rect 7941 1989 7975 2023
rect 8677 1989 8711 2023
rect 10425 1989 10459 2023
rect 10977 1989 11011 2023
rect 11989 1989 12023 2023
rect 12817 1989 12851 2023
rect 16773 1989 16807 2023
rect 17877 1989 17911 2023
rect 21465 1989 21499 2023
rect 22078 1989 22112 2023
rect 1409 1921 1443 1955
rect 1943 1951 1977 1985
rect 3249 1921 3283 1955
rect 3709 1921 3743 1955
rect 4445 1921 4479 1955
rect 4813 1921 4847 1955
rect 5273 1921 5307 1955
rect 5457 1921 5491 1955
rect 6745 1921 6779 1955
rect 7113 1921 7147 1955
rect 7573 1921 7607 1955
rect 8217 1921 8251 1955
rect 8953 1921 8987 1955
rect 9211 1951 9245 1985
rect 11805 1921 11839 1955
rect 12633 1921 12667 1955
rect 13553 1921 13587 1955
rect 13829 1921 13863 1955
rect 14289 1921 14323 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 15669 1921 15703 1955
rect 16129 1921 16163 1955
rect 17325 1921 17359 1955
rect 18521 1921 18555 1955
rect 19717 1921 19751 1955
rect 20821 1921 20855 1955
rect 23305 1921 23339 1955
rect 1685 1853 1719 1887
rect 4169 1853 4203 1887
rect 18613 1853 18647 1887
rect 18889 1853 18923 1887
rect 19993 1853 20027 1887
rect 21833 1853 21867 1887
rect 23765 1853 23799 1887
rect 3433 1785 3467 1819
rect 4997 1785 5031 1819
rect 6929 1785 6963 1819
rect 7297 1785 7331 1819
rect 13369 1785 13403 1819
rect 1593 1717 1627 1751
rect 5733 1717 5767 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11621 1717 11655 1751
rect 12081 1717 12115 1751
rect 12449 1717 12483 1751
rect 12909 1717 12943 1751
rect 13645 1717 13679 1751
rect 14105 1717 14139 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15761 1717 15795 1751
rect 16313 1717 16347 1751
rect 16865 1717 16899 1751
rect 17417 1717 17451 1751
rect 17969 1717 18003 1751
rect 1593 1513 1627 1547
rect 8677 1513 8711 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 17969 1513 18003 1547
rect 18521 1513 18555 1547
rect 20545 1513 20579 1547
rect 2513 1445 2547 1479
rect 11529 1445 11563 1479
rect 16957 1445 16991 1479
rect 17509 1445 17543 1479
rect 9597 1377 9631 1411
rect 10885 1377 10919 1411
rect 1409 1309 1443 1343
rect 1961 1309 1995 1343
rect 3065 1309 3099 1343
rect 3617 1309 3651 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 5273 1309 5307 1343
rect 5549 1309 5583 1343
rect 6377 1309 6411 1343
rect 7021 1309 7055 1343
rect 7941 1309 7975 1343
rect 8401 1309 8435 1343
rect 8493 1309 8527 1343
rect 9137 1309 9171 1343
rect 9781 1309 9815 1343
rect 10149 1309 10183 1343
rect 10609 1309 10643 1343
rect 11069 1309 11103 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12265 1309 12299 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 13829 1309 13863 1343
rect 14657 1309 14691 1343
rect 15301 1309 15335 1343
rect 16497 1309 16531 1343
rect 17325 1309 17359 1343
rect 17877 1309 17911 1343
rect 18429 1309 18463 1343
rect 18889 1309 18923 1343
rect 21465 1309 21499 1343
rect 21649 1309 21683 1343
rect 22201 1309 22235 1343
rect 22376 1309 22410 1343
rect 22477 1309 22511 1343
rect 24225 1309 24259 1343
rect 1777 1241 1811 1275
rect 2329 1241 2363 1275
rect 2697 1241 2731 1275
rect 4997 1241 5031 1275
rect 7389 1241 7423 1275
rect 7757 1241 7791 1275
rect 9321 1241 9355 1275
rect 14197 1241 14231 1275
rect 15853 1241 15887 1275
rect 16773 1241 16807 1275
rect 19257 1241 19291 1275
rect 21189 1241 21223 1275
rect 21925 1241 21959 1275
rect 22109 1241 22143 1275
rect 2789 1173 2823 1207
rect 3249 1173 3283 1207
rect 3433 1173 3467 1207
rect 5089 1173 5123 1207
rect 6561 1173 6595 1207
rect 7113 1173 7147 1207
rect 7481 1173 7515 1207
rect 8217 1173 8251 1207
rect 8953 1173 8987 1207
rect 9965 1173 9999 1207
rect 10333 1173 10367 1207
rect 11253 1173 11287 1207
rect 11989 1173 12023 1207
rect 12357 1173 12391 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 13645 1173 13679 1207
rect 14841 1173 14875 1207
rect 19073 1173 19107 1207
rect 21281 1173 21315 1207
rect 21649 1173 21683 1207
rect 22385 1173 22419 1207
<< metal1 >>
rect 18598 43800 18604 43852
rect 18656 43840 18662 43852
rect 20714 43840 20720 43852
rect 18656 43812 20720 43840
rect 18656 43800 18662 43812
rect 20714 43800 20720 43812
rect 20772 43800 20778 43852
rect 19426 43732 19432 43784
rect 19484 43772 19490 43784
rect 19794 43772 19800 43784
rect 19484 43744 19800 43772
rect 19484 43732 19490 43744
rect 19794 43732 19800 43744
rect 19852 43732 19858 43784
rect 15286 43664 15292 43716
rect 15344 43704 15350 43716
rect 15344 43676 22094 43704
rect 15344 43664 15350 43676
rect 5350 43596 5356 43648
rect 5408 43636 5414 43648
rect 10502 43636 10508 43648
rect 5408 43608 10508 43636
rect 5408 43596 5414 43608
rect 10502 43596 10508 43608
rect 10560 43596 10566 43648
rect 17494 43596 17500 43648
rect 17552 43636 17558 43648
rect 21266 43636 21272 43648
rect 17552 43608 21272 43636
rect 17552 43596 17558 43608
rect 21266 43596 21272 43608
rect 21324 43596 21330 43648
rect 22066 43636 22094 43676
rect 24394 43636 24400 43648
rect 22066 43608 24400 43636
rect 24394 43596 24400 43608
rect 24452 43596 24458 43648
rect 1104 43546 25000 43568
rect 1104 43494 6884 43546
rect 6936 43494 6948 43546
rect 7000 43494 7012 43546
rect 7064 43494 7076 43546
rect 7128 43494 7140 43546
rect 7192 43494 12818 43546
rect 12870 43494 12882 43546
rect 12934 43494 12946 43546
rect 12998 43494 13010 43546
rect 13062 43494 13074 43546
rect 13126 43494 18752 43546
rect 18804 43494 18816 43546
rect 18868 43494 18880 43546
rect 18932 43494 18944 43546
rect 18996 43494 19008 43546
rect 19060 43494 24686 43546
rect 24738 43494 24750 43546
rect 24802 43494 24814 43546
rect 24866 43494 24878 43546
rect 24930 43494 24942 43546
rect 24994 43494 25000 43546
rect 1104 43472 25000 43494
rect 1854 43392 1860 43444
rect 1912 43392 1918 43444
rect 2777 43435 2835 43441
rect 2777 43401 2789 43435
rect 2823 43432 2835 43435
rect 2958 43432 2964 43444
rect 2823 43404 2964 43432
rect 2823 43401 2835 43404
rect 2777 43395 2835 43401
rect 2958 43392 2964 43404
rect 3016 43392 3022 43444
rect 3145 43435 3203 43441
rect 3145 43401 3157 43435
rect 3191 43401 3203 43435
rect 3145 43395 3203 43401
rect 382 43324 388 43376
rect 440 43364 446 43376
rect 3160 43364 3188 43395
rect 4338 43392 4344 43444
rect 4396 43432 4402 43444
rect 4617 43435 4675 43441
rect 4617 43432 4629 43435
rect 4396 43404 4629 43432
rect 4396 43392 4402 43404
rect 4617 43401 4629 43404
rect 4663 43401 4675 43435
rect 4617 43395 4675 43401
rect 5534 43392 5540 43444
rect 5592 43392 5598 43444
rect 6089 43435 6147 43441
rect 6089 43401 6101 43435
rect 6135 43432 6147 43435
rect 6270 43432 6276 43444
rect 6135 43404 6276 43432
rect 6135 43401 6147 43404
rect 6089 43395 6147 43401
rect 6270 43392 6276 43404
rect 6328 43392 6334 43444
rect 6365 43435 6423 43441
rect 6365 43401 6377 43435
rect 6411 43432 6423 43435
rect 6411 43404 6776 43432
rect 6411 43401 6423 43404
rect 6365 43395 6423 43401
rect 440 43336 3188 43364
rect 440 43324 446 43336
rect 3418 43324 3424 43376
rect 3476 43364 3482 43376
rect 6748 43373 6776 43404
rect 6822 43392 6828 43444
rect 6880 43392 6886 43444
rect 7377 43435 7435 43441
rect 7377 43401 7389 43435
rect 7423 43432 7435 43435
rect 7650 43432 7656 43444
rect 7423 43404 7656 43432
rect 7423 43401 7435 43404
rect 7377 43395 7435 43401
rect 7650 43392 7656 43404
rect 7708 43392 7714 43444
rect 7745 43435 7803 43441
rect 7745 43401 7757 43435
rect 7791 43432 7803 43435
rect 7926 43432 7932 43444
rect 7791 43404 7932 43432
rect 7791 43401 7803 43404
rect 7745 43395 7803 43401
rect 7926 43392 7932 43404
rect 7984 43392 7990 43444
rect 8297 43435 8355 43441
rect 8297 43401 8309 43435
rect 8343 43432 8355 43435
rect 8478 43432 8484 43444
rect 8343 43404 8484 43432
rect 8343 43401 8355 43404
rect 8297 43395 8355 43401
rect 8478 43392 8484 43404
rect 8536 43392 8542 43444
rect 8665 43435 8723 43441
rect 8665 43401 8677 43435
rect 8711 43432 8723 43435
rect 9030 43432 9036 43444
rect 8711 43404 9036 43432
rect 8711 43401 8723 43404
rect 8665 43395 8723 43401
rect 9030 43392 9036 43404
rect 9088 43392 9094 43444
rect 9217 43435 9275 43441
rect 9217 43401 9229 43435
rect 9263 43432 9275 43435
rect 9582 43432 9588 43444
rect 9263 43404 9588 43432
rect 9263 43401 9275 43404
rect 9217 43395 9275 43401
rect 9582 43392 9588 43404
rect 9640 43392 9646 43444
rect 9769 43435 9827 43441
rect 9769 43401 9781 43435
rect 9815 43432 9827 43435
rect 9858 43432 9864 43444
rect 9815 43404 9864 43432
rect 9815 43401 9827 43404
rect 9769 43395 9827 43401
rect 9858 43392 9864 43404
rect 9916 43392 9922 43444
rect 10502 43392 10508 43444
rect 10560 43392 10566 43444
rect 13354 43392 13360 43444
rect 13412 43432 13418 43444
rect 15197 43435 15255 43441
rect 13412 43404 14228 43432
rect 13412 43392 13418 43404
rect 4525 43367 4583 43373
rect 4525 43364 4537 43367
rect 3476 43336 4537 43364
rect 3476 43324 3482 43336
rect 4525 43333 4537 43336
rect 4571 43333 4583 43367
rect 4525 43327 4583 43333
rect 6733 43367 6791 43373
rect 6733 43333 6745 43367
rect 6779 43333 6791 43367
rect 6733 43327 6791 43333
rect 8021 43367 8079 43373
rect 8021 43333 8033 43367
rect 8067 43364 8079 43367
rect 8570 43364 8576 43376
rect 8067 43336 8576 43364
rect 8067 43333 8079 43336
rect 8021 43327 8079 43333
rect 8570 43324 8576 43336
rect 8628 43324 8634 43376
rect 9398 43364 9404 43376
rect 8956 43336 9404 43364
rect 1210 43256 1216 43308
rect 1268 43296 1274 43308
rect 1581 43299 1639 43305
rect 1581 43296 1593 43299
rect 1268 43268 1593 43296
rect 1268 43256 1274 43268
rect 1581 43265 1593 43268
rect 1627 43265 1639 43299
rect 1581 43259 1639 43265
rect 1762 43256 1768 43308
rect 1820 43256 1826 43308
rect 2498 43256 2504 43308
rect 2556 43256 2562 43308
rect 3050 43256 3056 43308
rect 3108 43256 3114 43308
rect 3973 43300 4031 43305
rect 3973 43299 4106 43300
rect 3973 43265 3985 43299
rect 4019 43272 4106 43299
rect 4019 43265 4031 43272
rect 3973 43259 4031 43265
rect 4078 43228 4106 43272
rect 5258 43256 5264 43308
rect 5316 43256 5322 43308
rect 5905 43299 5963 43305
rect 5905 43265 5917 43299
rect 5951 43296 5963 43299
rect 5994 43296 6000 43308
rect 5951 43268 6000 43296
rect 5951 43265 5963 43268
rect 5905 43259 5963 43265
rect 5994 43256 6000 43268
rect 6052 43256 6058 43308
rect 6270 43256 6276 43308
rect 6328 43296 6334 43308
rect 6549 43299 6607 43305
rect 6549 43296 6561 43299
rect 6328 43268 6561 43296
rect 6328 43256 6334 43268
rect 6549 43265 6561 43268
rect 6595 43265 6607 43299
rect 6549 43259 6607 43265
rect 7193 43299 7251 43305
rect 7193 43265 7205 43299
rect 7239 43296 7251 43299
rect 7282 43296 7288 43308
rect 7239 43268 7288 43296
rect 7239 43265 7251 43268
rect 7193 43259 7251 43265
rect 7282 43256 7288 43268
rect 7340 43256 7346 43308
rect 7561 43299 7619 43305
rect 7561 43265 7573 43299
rect 7607 43296 7619 43299
rect 8110 43296 8116 43308
rect 7607 43268 8116 43296
rect 7607 43265 7619 43268
rect 7561 43259 7619 43265
rect 8110 43256 8116 43268
rect 8168 43256 8174 43308
rect 8481 43299 8539 43305
rect 8481 43265 8493 43299
rect 8527 43296 8539 43299
rect 8956 43296 8984 43336
rect 9398 43324 9404 43336
rect 9456 43324 9462 43376
rect 9508 43336 12204 43364
rect 9508 43305 9536 43336
rect 8527 43268 8984 43296
rect 9033 43299 9091 43305
rect 8527 43265 8539 43268
rect 8481 43259 8539 43265
rect 9033 43265 9045 43299
rect 9079 43265 9091 43299
rect 9033 43259 9091 43265
rect 9493 43299 9551 43305
rect 9493 43265 9505 43299
rect 9539 43265 9551 43299
rect 9493 43259 9551 43265
rect 4798 43228 4804 43240
rect 4078 43200 4804 43228
rect 4798 43188 4804 43200
rect 4856 43188 4862 43240
rect 9048 43228 9076 43259
rect 9950 43256 9956 43308
rect 10008 43256 10014 43308
rect 10318 43256 10324 43308
rect 10376 43256 10382 43308
rect 10686 43256 10692 43308
rect 10744 43256 10750 43308
rect 11054 43256 11060 43308
rect 11112 43256 11118 43308
rect 11238 43256 11244 43308
rect 11296 43296 11302 43308
rect 11517 43299 11575 43305
rect 11517 43296 11529 43299
rect 11296 43268 11529 43296
rect 11296 43256 11302 43268
rect 11517 43265 11529 43268
rect 11563 43265 11575 43299
rect 11517 43259 11575 43265
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 12176 43296 12204 43336
rect 12434 43324 12440 43376
rect 12492 43324 12498 43376
rect 12802 43324 12808 43376
rect 12860 43324 12866 43376
rect 13446 43324 13452 43376
rect 13504 43364 13510 43376
rect 14200 43373 14228 43404
rect 15197 43401 15209 43435
rect 15243 43432 15255 43435
rect 15286 43432 15292 43444
rect 15243 43404 15292 43432
rect 15243 43401 15255 43404
rect 15197 43395 15255 43401
rect 15286 43392 15292 43404
rect 15344 43392 15350 43444
rect 17034 43392 17040 43444
rect 17092 43432 17098 43444
rect 17092 43404 18000 43432
rect 17092 43392 17098 43404
rect 13725 43367 13783 43373
rect 13725 43364 13737 43367
rect 13504 43336 13737 43364
rect 13504 43324 13510 43336
rect 13725 43333 13737 43336
rect 13771 43333 13783 43367
rect 13725 43327 13783 43333
rect 14185 43367 14243 43373
rect 14185 43333 14197 43367
rect 14231 43333 14243 43367
rect 14185 43327 14243 43333
rect 14734 43324 14740 43376
rect 14792 43324 14798 43376
rect 14826 43324 14832 43376
rect 14884 43364 14890 43376
rect 15105 43367 15163 43373
rect 15105 43364 15117 43367
rect 14884 43336 15117 43364
rect 14884 43324 14890 43336
rect 15105 43333 15117 43336
rect 15151 43333 15163 43367
rect 15105 43327 15163 43333
rect 15562 43324 15568 43376
rect 15620 43324 15626 43376
rect 15930 43324 15936 43376
rect 15988 43364 15994 43376
rect 16301 43367 16359 43373
rect 16301 43364 16313 43367
rect 15988 43336 16313 43364
rect 15988 43324 15994 43336
rect 16301 43333 16313 43336
rect 16347 43333 16359 43367
rect 16301 43327 16359 43333
rect 16390 43324 16396 43376
rect 16448 43364 16454 43376
rect 16761 43367 16819 43373
rect 16761 43364 16773 43367
rect 16448 43336 16773 43364
rect 16448 43324 16454 43336
rect 16761 43333 16773 43336
rect 16807 43333 16819 43367
rect 16761 43327 16819 43333
rect 16850 43324 16856 43376
rect 16908 43364 16914 43376
rect 16908 43336 17816 43364
rect 16908 43324 16914 43336
rect 13630 43296 13636 43308
rect 12176 43268 13636 43296
rect 13630 43256 13636 43268
rect 13688 43256 13694 43308
rect 15838 43256 15844 43308
rect 15896 43256 15902 43308
rect 17788 43305 17816 43336
rect 17497 43299 17555 43305
rect 17497 43296 17509 43299
rect 16684 43268 17509 43296
rect 9674 43228 9680 43240
rect 9048 43200 9680 43228
rect 9674 43188 9680 43200
rect 9732 43188 9738 43240
rect 16485 43231 16543 43237
rect 16485 43228 16497 43231
rect 9784 43200 16497 43228
rect 3789 43163 3847 43169
rect 3789 43129 3801 43163
rect 3835 43160 3847 43163
rect 4706 43160 4712 43172
rect 3835 43132 4712 43160
rect 3835 43129 3847 43132
rect 3789 43123 3847 43129
rect 4706 43120 4712 43132
rect 4764 43120 4770 43172
rect 9122 43120 9128 43172
rect 9180 43160 9186 43172
rect 9784 43160 9812 43200
rect 16485 43197 16497 43200
rect 16531 43197 16543 43231
rect 16485 43191 16543 43197
rect 9180 43132 9812 43160
rect 10137 43163 10195 43169
rect 9180 43120 9186 43132
rect 10137 43129 10149 43163
rect 10183 43160 10195 43163
rect 10183 43132 14780 43160
rect 10183 43129 10195 43132
rect 10137 43123 10195 43129
rect 14752 43104 14780 43132
rect 14918 43120 14924 43172
rect 14976 43120 14982 43172
rect 15562 43120 15568 43172
rect 15620 43160 15626 43172
rect 15620 43132 16068 43160
rect 15620 43120 15626 43132
rect 1397 43095 1455 43101
rect 1397 43061 1409 43095
rect 1443 43092 1455 43095
rect 1670 43092 1676 43104
rect 1443 43064 1676 43092
rect 1443 43061 1455 43064
rect 1397 43055 1455 43061
rect 1670 43052 1676 43064
rect 1728 43052 1734 43104
rect 3602 43052 3608 43104
rect 3660 43092 3666 43104
rect 4249 43095 4307 43101
rect 4249 43092 4261 43095
rect 3660 43064 4261 43092
rect 3660 43052 3666 43064
rect 4249 43061 4261 43064
rect 4295 43092 4307 43095
rect 4430 43092 4436 43104
rect 4295 43064 4436 43092
rect 4295 43061 4307 43064
rect 4249 43055 4307 43061
rect 4430 43052 4436 43064
rect 4488 43052 4494 43104
rect 9398 43052 9404 43104
rect 9456 43092 9462 43104
rect 10594 43092 10600 43104
rect 9456 43064 10600 43092
rect 9456 43052 9462 43064
rect 10594 43052 10600 43064
rect 10652 43052 10658 43104
rect 10870 43052 10876 43104
rect 10928 43052 10934 43104
rect 11238 43052 11244 43104
rect 11296 43052 11302 43104
rect 11698 43052 11704 43104
rect 11756 43052 11762 43104
rect 12250 43052 12256 43104
rect 12308 43052 12314 43104
rect 12526 43052 12532 43104
rect 12584 43052 12590 43104
rect 12618 43052 12624 43104
rect 12676 43092 12682 43104
rect 12897 43095 12955 43101
rect 12897 43092 12909 43095
rect 12676 43064 12909 43092
rect 12676 43052 12682 43064
rect 12897 43061 12909 43064
rect 12943 43061 12955 43095
rect 12897 43055 12955 43061
rect 13814 43052 13820 43104
rect 13872 43052 13878 43104
rect 14274 43052 14280 43104
rect 14332 43052 14338 43104
rect 14734 43052 14740 43104
rect 14792 43052 14798 43104
rect 15654 43052 15660 43104
rect 15712 43052 15718 43104
rect 16040 43101 16068 43132
rect 16298 43120 16304 43172
rect 16356 43160 16362 43172
rect 16684 43160 16712 43268
rect 17497 43265 17509 43268
rect 17543 43265 17555 43299
rect 17497 43259 17555 43265
rect 17773 43299 17831 43305
rect 17773 43265 17785 43299
rect 17819 43265 17831 43299
rect 17972 43296 18000 43404
rect 18138 43392 18144 43444
rect 18196 43432 18202 43444
rect 20073 43435 20131 43441
rect 18196 43404 19472 43432
rect 18196 43392 18202 43404
rect 18230 43324 18236 43376
rect 18288 43364 18294 43376
rect 18288 43336 18644 43364
rect 18288 43324 18294 43336
rect 18616 43305 18644 43336
rect 18049 43299 18107 43305
rect 18049 43296 18061 43299
rect 17972 43268 18061 43296
rect 17773 43259 17831 43265
rect 18049 43265 18061 43268
rect 18095 43265 18107 43299
rect 18049 43259 18107 43265
rect 18325 43299 18383 43305
rect 18325 43265 18337 43299
rect 18371 43265 18383 43299
rect 18325 43259 18383 43265
rect 18601 43299 18659 43305
rect 18601 43265 18613 43299
rect 18647 43265 18659 43299
rect 18601 43259 18659 43265
rect 18877 43299 18935 43305
rect 18877 43265 18889 43299
rect 18923 43296 18935 43299
rect 19334 43296 19340 43308
rect 18923 43268 19340 43296
rect 18923 43265 18935 43268
rect 18877 43259 18935 43265
rect 17402 43188 17408 43240
rect 17460 43228 17466 43240
rect 18340 43228 18368 43259
rect 19334 43256 19340 43268
rect 19392 43256 19398 43308
rect 19444 43305 19472 43404
rect 20073 43401 20085 43435
rect 20119 43432 20131 43435
rect 20346 43432 20352 43444
rect 20119 43404 20352 43432
rect 20119 43401 20131 43404
rect 20073 43395 20131 43401
rect 20346 43392 20352 43404
rect 20404 43392 20410 43444
rect 20622 43392 20628 43444
rect 20680 43432 20686 43444
rect 20993 43435 21051 43441
rect 20993 43432 21005 43435
rect 20680 43404 21005 43432
rect 20680 43392 20686 43404
rect 20993 43401 21005 43404
rect 21039 43401 21051 43435
rect 20993 43395 21051 43401
rect 21174 43392 21180 43444
rect 21232 43432 21238 43444
rect 22005 43435 22063 43441
rect 22005 43432 22017 43435
rect 21232 43404 22017 43432
rect 21232 43392 21238 43404
rect 22005 43401 22017 43404
rect 22051 43401 22063 43435
rect 22005 43395 22063 43401
rect 22373 43435 22431 43441
rect 22373 43401 22385 43435
rect 22419 43401 22431 43435
rect 22373 43395 22431 43401
rect 19978 43324 19984 43376
rect 20036 43364 20042 43376
rect 20036 43336 21404 43364
rect 20036 43324 20042 43336
rect 19429 43299 19487 43305
rect 19429 43265 19441 43299
rect 19475 43265 19487 43299
rect 19429 43259 19487 43265
rect 19702 43256 19708 43308
rect 19760 43256 19766 43308
rect 19886 43256 19892 43308
rect 19944 43256 19950 43308
rect 20349 43299 20407 43305
rect 20349 43265 20361 43299
rect 20395 43265 20407 43299
rect 20349 43259 20407 43265
rect 17460 43200 18368 43228
rect 17460 43188 17466 43200
rect 16356 43132 16712 43160
rect 16356 43120 16362 43132
rect 17770 43120 17776 43172
rect 17828 43160 17834 43172
rect 18141 43163 18199 43169
rect 18141 43160 18153 43163
rect 17828 43132 18153 43160
rect 17828 43120 17834 43132
rect 18141 43129 18153 43132
rect 18187 43129 18199 43163
rect 18141 43123 18199 43129
rect 18230 43120 18236 43172
rect 18288 43160 18294 43172
rect 18693 43163 18751 43169
rect 18693 43160 18705 43163
rect 18288 43132 18705 43160
rect 18288 43120 18294 43132
rect 18693 43129 18705 43132
rect 18739 43129 18751 43163
rect 18693 43123 18751 43129
rect 19150 43120 19156 43172
rect 19208 43160 19214 43172
rect 19702 43160 19708 43172
rect 19208 43132 19708 43160
rect 19208 43120 19214 43132
rect 19702 43120 19708 43132
rect 19760 43120 19766 43172
rect 16025 43095 16083 43101
rect 16025 43061 16037 43095
rect 16071 43061 16083 43095
rect 16025 43055 16083 43061
rect 16850 43052 16856 43104
rect 16908 43052 16914 43104
rect 17313 43095 17371 43101
rect 17313 43061 17325 43095
rect 17359 43092 17371 43095
rect 17494 43092 17500 43104
rect 17359 43064 17500 43092
rect 17359 43061 17371 43064
rect 17313 43055 17371 43061
rect 17494 43052 17500 43064
rect 17552 43052 17558 43104
rect 17586 43052 17592 43104
rect 17644 43052 17650 43104
rect 17862 43052 17868 43104
rect 17920 43052 17926 43104
rect 18046 43052 18052 43104
rect 18104 43092 18110 43104
rect 18417 43095 18475 43101
rect 18417 43092 18429 43095
rect 18104 43064 18429 43092
rect 18104 43052 18110 43064
rect 18417 43061 18429 43064
rect 18463 43061 18475 43095
rect 18417 43055 18475 43061
rect 18598 43052 18604 43104
rect 18656 43092 18662 43104
rect 19245 43095 19303 43101
rect 19245 43092 19257 43095
rect 18656 43064 19257 43092
rect 18656 43052 18662 43064
rect 19245 43061 19257 43064
rect 19291 43061 19303 43095
rect 19245 43055 19303 43061
rect 19518 43052 19524 43104
rect 19576 43052 19582 43104
rect 20364 43092 20392 43259
rect 20438 43256 20444 43308
rect 20496 43296 20502 43308
rect 21376 43305 21404 43336
rect 21542 43324 21548 43376
rect 21600 43364 21606 43376
rect 22388 43364 22416 43395
rect 23106 43392 23112 43444
rect 23164 43432 23170 43444
rect 23477 43435 23535 43441
rect 23477 43432 23489 43435
rect 23164 43404 23489 43432
rect 23164 43392 23170 43404
rect 23477 43401 23489 43404
rect 23523 43401 23535 43435
rect 23477 43395 23535 43401
rect 21600 43336 22416 43364
rect 21600 43324 21606 43336
rect 20901 43299 20959 43305
rect 20901 43296 20913 43299
rect 20496 43268 20913 43296
rect 20496 43256 20502 43268
rect 20901 43265 20913 43268
rect 20947 43265 20959 43299
rect 20901 43259 20959 43265
rect 21361 43299 21419 43305
rect 21361 43265 21373 43299
rect 21407 43265 21419 43299
rect 21361 43259 21419 43265
rect 21634 43256 21640 43308
rect 21692 43296 21698 43308
rect 21821 43299 21879 43305
rect 21821 43296 21833 43299
rect 21692 43268 21833 43296
rect 21692 43256 21698 43268
rect 21821 43265 21833 43268
rect 21867 43265 21879 43299
rect 21821 43259 21879 43265
rect 22281 43299 22339 43305
rect 22281 43265 22293 43299
rect 22327 43296 22339 43299
rect 22370 43296 22376 43308
rect 22327 43268 22376 43296
rect 22327 43265 22339 43268
rect 22281 43259 22339 43265
rect 22370 43256 22376 43268
rect 22428 43256 22434 43308
rect 22646 43256 22652 43308
rect 22704 43296 22710 43308
rect 22833 43299 22891 43305
rect 22833 43296 22845 43299
rect 22704 43268 22845 43296
rect 22704 43256 22710 43268
rect 22833 43265 22845 43268
rect 22879 43265 22891 43299
rect 22833 43259 22891 43265
rect 23385 43299 23443 43305
rect 23385 43265 23397 43299
rect 23431 43265 23443 43299
rect 23385 43259 23443 43265
rect 20625 43231 20683 43237
rect 20625 43197 20637 43231
rect 20671 43228 20683 43231
rect 22554 43228 22560 43240
rect 20671 43200 22560 43228
rect 20671 43197 20683 43200
rect 20625 43191 20683 43197
rect 22554 43188 22560 43200
rect 22612 43188 22618 43240
rect 20898 43120 20904 43172
rect 20956 43160 20962 43172
rect 21545 43163 21603 43169
rect 21545 43160 21557 43163
rect 20956 43132 21557 43160
rect 20956 43120 20962 43132
rect 21545 43129 21557 43132
rect 21591 43129 21603 43163
rect 21545 43123 21603 43129
rect 22186 43120 22192 43172
rect 22244 43160 22250 43172
rect 23400 43160 23428 43259
rect 23474 43256 23480 43308
rect 23532 43296 23538 43308
rect 23937 43299 23995 43305
rect 23937 43296 23949 43299
rect 23532 43268 23949 43296
rect 23532 43256 23538 43268
rect 23937 43265 23949 43268
rect 23983 43265 23995 43299
rect 23937 43259 23995 43265
rect 22244 43132 23428 43160
rect 22244 43120 22250 43132
rect 21358 43092 21364 43104
rect 20364 43064 21364 43092
rect 21358 43052 21364 43064
rect 21416 43052 21422 43104
rect 21910 43052 21916 43104
rect 21968 43092 21974 43104
rect 22925 43095 22983 43101
rect 22925 43092 22937 43095
rect 21968 43064 22937 43092
rect 21968 43052 21974 43064
rect 22925 43061 22937 43064
rect 22971 43061 22983 43095
rect 22925 43055 22983 43061
rect 24118 43052 24124 43104
rect 24176 43052 24182 43104
rect 1104 43002 24840 43024
rect 1104 42950 3917 43002
rect 3969 42950 3981 43002
rect 4033 42950 4045 43002
rect 4097 42950 4109 43002
rect 4161 42950 4173 43002
rect 4225 42950 9851 43002
rect 9903 42950 9915 43002
rect 9967 42950 9979 43002
rect 10031 42950 10043 43002
rect 10095 42950 10107 43002
rect 10159 42950 15785 43002
rect 15837 42950 15849 43002
rect 15901 42950 15913 43002
rect 15965 42950 15977 43002
rect 16029 42950 16041 43002
rect 16093 42950 21719 43002
rect 21771 42950 21783 43002
rect 21835 42950 21847 43002
rect 21899 42950 21911 43002
rect 21963 42950 21975 43002
rect 22027 42950 24840 43002
rect 1104 42928 24840 42950
rect 2222 42848 2228 42900
rect 2280 42848 2286 42900
rect 3326 42848 3332 42900
rect 3384 42848 3390 42900
rect 6086 42848 6092 42900
rect 6144 42848 6150 42900
rect 6822 42848 6828 42900
rect 6880 42848 6886 42900
rect 7374 42848 7380 42900
rect 7432 42848 7438 42900
rect 9122 42888 9128 42900
rect 7484 42860 9128 42888
rect 4264 42792 5488 42820
rect 1394 42712 1400 42764
rect 1452 42752 1458 42764
rect 1765 42755 1823 42761
rect 1765 42752 1777 42755
rect 1452 42724 1777 42752
rect 1452 42712 1458 42724
rect 1765 42721 1777 42724
rect 1811 42721 1823 42755
rect 3694 42752 3700 42764
rect 1765 42715 1823 42721
rect 1872 42724 3700 42752
rect 14 42644 20 42696
rect 72 42684 78 42696
rect 1872 42684 1900 42724
rect 3694 42712 3700 42724
rect 3752 42712 3758 42764
rect 4264 42752 4292 42792
rect 4172 42724 4292 42752
rect 72 42656 1900 42684
rect 2133 42687 2191 42693
rect 72 42644 78 42656
rect 2133 42653 2145 42687
rect 2179 42684 2191 42687
rect 4172 42684 4200 42724
rect 4338 42712 4344 42764
rect 4396 42712 4402 42764
rect 4890 42712 4896 42764
rect 4948 42752 4954 42764
rect 5353 42755 5411 42761
rect 5353 42752 5365 42755
rect 4948 42724 5365 42752
rect 4948 42712 4954 42724
rect 5353 42721 5365 42724
rect 5399 42721 5411 42755
rect 5460 42752 5488 42792
rect 5534 42780 5540 42832
rect 5592 42820 5598 42832
rect 7484 42820 7512 42860
rect 9122 42848 9128 42860
rect 9180 42848 9186 42900
rect 9674 42848 9680 42900
rect 9732 42888 9738 42900
rect 10321 42891 10379 42897
rect 10321 42888 10333 42891
rect 9732 42860 10333 42888
rect 9732 42848 9738 42860
rect 10321 42857 10333 42860
rect 10367 42857 10379 42891
rect 10321 42851 10379 42857
rect 10594 42848 10600 42900
rect 10652 42848 10658 42900
rect 16850 42888 16856 42900
rect 12406 42860 16856 42888
rect 5592 42792 7512 42820
rect 5592 42780 5598 42792
rect 9214 42780 9220 42832
rect 9272 42820 9278 42832
rect 12406 42820 12434 42860
rect 16850 42848 16856 42860
rect 16908 42848 16914 42900
rect 17862 42848 17868 42900
rect 17920 42848 17926 42900
rect 18138 42848 18144 42900
rect 18196 42888 18202 42900
rect 18877 42891 18935 42897
rect 18877 42888 18889 42891
rect 18196 42860 18889 42888
rect 18196 42848 18202 42860
rect 18877 42857 18889 42860
rect 18923 42857 18935 42891
rect 18877 42851 18935 42857
rect 19306 42860 21220 42888
rect 9272 42792 12434 42820
rect 13173 42823 13231 42829
rect 9272 42780 9278 42792
rect 13173 42789 13185 42823
rect 13219 42789 13231 42823
rect 13173 42783 13231 42789
rect 8478 42752 8484 42764
rect 5460 42724 8484 42752
rect 5353 42715 5411 42721
rect 8478 42712 8484 42724
rect 8536 42712 8542 42764
rect 8665 42755 8723 42761
rect 8665 42721 8677 42755
rect 8711 42752 8723 42755
rect 8754 42752 8760 42764
rect 8711 42724 8760 42752
rect 8711 42721 8723 42724
rect 8665 42715 8723 42721
rect 8754 42712 8760 42724
rect 8812 42712 8818 42764
rect 9306 42712 9312 42764
rect 9364 42752 9370 42764
rect 9769 42755 9827 42761
rect 9769 42752 9781 42755
rect 9364 42724 9781 42752
rect 9364 42712 9370 42724
rect 9769 42721 9781 42724
rect 9815 42721 9827 42755
rect 12250 42752 12256 42764
rect 9769 42715 9827 42721
rect 10060 42724 12256 42752
rect 2179 42656 4200 42684
rect 2179 42653 2191 42656
rect 2133 42647 2191 42653
rect 4246 42644 4252 42696
rect 4304 42684 4310 42696
rect 4525 42687 4583 42693
rect 4525 42684 4537 42687
rect 4304 42656 4537 42684
rect 4304 42644 4310 42656
rect 4525 42653 4537 42656
rect 4571 42653 4583 42687
rect 4525 42647 4583 42653
rect 4706 42644 4712 42696
rect 4764 42684 4770 42696
rect 5077 42687 5135 42693
rect 5077 42684 5089 42687
rect 4764 42656 5089 42684
rect 4764 42644 4770 42656
rect 5077 42653 5089 42656
rect 5123 42653 5135 42687
rect 5077 42647 5135 42653
rect 5534 42644 5540 42696
rect 5592 42644 5598 42696
rect 7558 42644 7564 42696
rect 7616 42684 7622 42696
rect 7745 42687 7803 42693
rect 7745 42684 7757 42687
rect 7616 42656 7757 42684
rect 7616 42644 7622 42656
rect 7745 42653 7757 42656
rect 7791 42653 7803 42687
rect 7745 42647 7803 42653
rect 8386 42644 8392 42696
rect 8444 42644 8450 42696
rect 9030 42644 9036 42696
rect 9088 42680 9094 42696
rect 9125 42687 9183 42693
rect 9125 42680 9137 42687
rect 9088 42653 9137 42680
rect 9171 42653 9183 42687
rect 9088 42652 9183 42653
rect 9088 42644 9094 42652
rect 9125 42647 9183 42652
rect 9398 42644 9404 42696
rect 9456 42684 9462 42696
rect 9950 42684 9956 42696
rect 9456 42656 9956 42684
rect 9456 42644 9462 42656
rect 9950 42644 9956 42656
rect 10008 42644 10014 42696
rect 10060 42693 10088 42724
rect 12250 42712 12256 42724
rect 12308 42712 12314 42764
rect 12434 42712 12440 42764
rect 12492 42752 12498 42764
rect 13188 42752 13216 42783
rect 14734 42780 14740 42832
rect 14792 42820 14798 42832
rect 17126 42820 17132 42832
rect 14792 42792 17132 42820
rect 14792 42780 14798 42792
rect 17126 42780 17132 42792
rect 17184 42780 17190 42832
rect 12492 42724 13216 42752
rect 12492 42712 12498 42724
rect 13814 42712 13820 42764
rect 13872 42752 13878 42764
rect 13872 42724 14688 42752
rect 13872 42712 13878 42724
rect 10045 42687 10103 42693
rect 10045 42653 10057 42687
rect 10091 42653 10103 42687
rect 10505 42687 10563 42693
rect 10505 42684 10517 42687
rect 10045 42647 10103 42653
rect 10152 42656 10517 42684
rect 1489 42619 1547 42625
rect 1489 42585 1501 42619
rect 1535 42616 1547 42619
rect 2314 42616 2320 42628
rect 1535 42588 2320 42616
rect 1535 42585 1547 42588
rect 1489 42579 1547 42585
rect 2314 42576 2320 42588
rect 2372 42576 2378 42628
rect 2685 42619 2743 42625
rect 2685 42585 2697 42619
rect 2731 42616 2743 42619
rect 2866 42616 2872 42628
rect 2731 42588 2872 42616
rect 2731 42585 2743 42588
rect 2685 42579 2743 42585
rect 2866 42576 2872 42588
rect 2924 42576 2930 42628
rect 3234 42576 3240 42628
rect 3292 42576 3298 42628
rect 4065 42619 4123 42625
rect 4065 42585 4077 42619
rect 4111 42616 4123 42619
rect 4430 42616 4436 42628
rect 4111 42588 4436 42616
rect 4111 42585 4123 42588
rect 4065 42579 4123 42585
rect 4430 42576 4436 42588
rect 4488 42576 4494 42628
rect 5994 42576 6000 42628
rect 6052 42576 6058 42628
rect 6733 42619 6791 42625
rect 6733 42585 6745 42619
rect 6779 42585 6791 42619
rect 6733 42579 6791 42585
rect 2774 42508 2780 42560
rect 2832 42508 2838 42560
rect 4614 42508 4620 42560
rect 4672 42548 4678 42560
rect 4709 42551 4767 42557
rect 4709 42548 4721 42551
rect 4672 42520 4721 42548
rect 4672 42508 4678 42520
rect 4709 42517 4721 42520
rect 4755 42517 4767 42551
rect 4709 42511 4767 42517
rect 5718 42508 5724 42560
rect 5776 42508 5782 42560
rect 5902 42508 5908 42560
rect 5960 42548 5966 42560
rect 6748 42548 6776 42579
rect 7282 42576 7288 42628
rect 7340 42576 7346 42628
rect 9493 42619 9551 42625
rect 9493 42616 9505 42619
rect 8956 42588 9505 42616
rect 5960 42520 6776 42548
rect 5960 42508 5966 42520
rect 7466 42508 7472 42560
rect 7524 42548 7530 42560
rect 8956 42557 8984 42588
rect 9493 42585 9505 42588
rect 9539 42585 9551 42619
rect 9493 42579 9551 42585
rect 9582 42576 9588 42628
rect 9640 42616 9646 42628
rect 10152 42616 10180 42656
rect 10505 42653 10517 42656
rect 10551 42653 10563 42687
rect 10505 42647 10563 42653
rect 10781 42687 10839 42693
rect 10781 42653 10793 42687
rect 10827 42653 10839 42687
rect 10781 42647 10839 42653
rect 9640 42588 10180 42616
rect 9640 42576 9646 42588
rect 10410 42576 10416 42628
rect 10468 42616 10474 42628
rect 10796 42616 10824 42647
rect 11606 42644 11612 42696
rect 11664 42644 11670 42696
rect 11882 42644 11888 42696
rect 11940 42644 11946 42696
rect 12713 42687 12771 42693
rect 12713 42653 12725 42687
rect 12759 42653 12771 42687
rect 12713 42647 12771 42653
rect 10468 42588 10824 42616
rect 10468 42576 10474 42588
rect 11330 42576 11336 42628
rect 11388 42616 11394 42628
rect 12728 42616 12756 42647
rect 12986 42644 12992 42696
rect 13044 42644 13050 42696
rect 14090 42644 14096 42696
rect 14148 42644 14154 42696
rect 14366 42644 14372 42696
rect 14424 42644 14430 42696
rect 14660 42693 14688 42724
rect 15194 42712 15200 42764
rect 15252 42752 15258 42764
rect 17880 42752 17908 42848
rect 18322 42780 18328 42832
rect 18380 42820 18386 42832
rect 19306 42820 19334 42860
rect 18380 42792 19334 42820
rect 21085 42823 21143 42829
rect 18380 42780 18386 42792
rect 21085 42789 21097 42823
rect 21131 42789 21143 42823
rect 21085 42783 21143 42789
rect 18598 42752 18604 42764
rect 15252 42724 15608 42752
rect 15252 42712 15258 42724
rect 14645 42687 14703 42693
rect 14645 42653 14657 42687
rect 14691 42653 14703 42687
rect 14645 42647 14703 42653
rect 15286 42644 15292 42696
rect 15344 42644 15350 42696
rect 15580 42693 15608 42724
rect 17420 42724 17908 42752
rect 18432 42724 18604 42752
rect 15565 42687 15623 42693
rect 15565 42653 15577 42687
rect 15611 42653 15623 42687
rect 15565 42647 15623 42653
rect 16482 42644 16488 42696
rect 16540 42644 16546 42696
rect 16574 42644 16580 42696
rect 16632 42644 16638 42696
rect 17420 42693 17448 42724
rect 17129 42687 17187 42693
rect 17129 42653 17141 42687
rect 17175 42653 17187 42687
rect 17129 42647 17187 42653
rect 17405 42687 17463 42693
rect 17405 42653 17417 42687
rect 17451 42653 17463 42687
rect 17405 42647 17463 42653
rect 13262 42616 13268 42628
rect 11388 42588 12112 42616
rect 12728 42588 13268 42616
rect 11388 42576 11394 42588
rect 7929 42551 7987 42557
rect 7929 42548 7941 42551
rect 7524 42520 7941 42548
rect 7524 42508 7530 42520
rect 7929 42517 7941 42520
rect 7975 42517 7987 42551
rect 7929 42511 7987 42517
rect 8941 42551 8999 42557
rect 8941 42517 8953 42551
rect 8987 42517 8999 42551
rect 8941 42511 8999 42517
rect 9122 42508 9128 42560
rect 9180 42548 9186 42560
rect 10229 42551 10287 42557
rect 10229 42548 10241 42551
rect 9180 42520 10241 42548
rect 9180 42508 9186 42520
rect 10229 42517 10241 42520
rect 10275 42517 10287 42551
rect 10229 42511 10287 42517
rect 11790 42508 11796 42560
rect 11848 42508 11854 42560
rect 12084 42557 12112 42588
rect 13262 42576 13268 42588
rect 13320 42576 13326 42628
rect 14734 42576 14740 42628
rect 14792 42616 14798 42628
rect 17144 42616 17172 42647
rect 17586 42644 17592 42696
rect 17644 42644 17650 42696
rect 17681 42687 17739 42693
rect 17681 42653 17693 42687
rect 17727 42684 17739 42687
rect 17770 42684 17776 42696
rect 17727 42656 17776 42684
rect 17727 42653 17739 42656
rect 17681 42647 17739 42653
rect 17770 42644 17776 42656
rect 17828 42644 17834 42696
rect 17957 42687 18015 42693
rect 17957 42653 17969 42687
rect 18003 42684 18015 42687
rect 18046 42684 18052 42696
rect 18003 42656 18052 42684
rect 18003 42653 18015 42656
rect 17957 42647 18015 42653
rect 18046 42644 18052 42656
rect 18104 42644 18110 42696
rect 18233 42687 18291 42693
rect 18233 42653 18245 42687
rect 18279 42684 18291 42687
rect 18432 42684 18460 42724
rect 18598 42712 18604 42724
rect 18656 42712 18662 42764
rect 21100 42752 21128 42783
rect 18708 42724 21128 42752
rect 18279 42656 18460 42684
rect 18509 42687 18567 42693
rect 18279 42653 18291 42656
rect 18233 42647 18291 42653
rect 18509 42653 18521 42687
rect 18555 42684 18567 42687
rect 18708 42684 18736 42724
rect 18555 42656 18736 42684
rect 18555 42653 18567 42656
rect 18509 42647 18567 42653
rect 18782 42644 18788 42696
rect 18840 42644 18846 42696
rect 19058 42644 19064 42696
rect 19116 42644 19122 42696
rect 21192 42684 21220 42860
rect 21266 42780 21272 42832
rect 21324 42820 21330 42832
rect 21324 42792 22094 42820
rect 21324 42780 21330 42792
rect 21269 42687 21327 42693
rect 21269 42684 21281 42687
rect 21192 42656 21281 42684
rect 21269 42653 21281 42656
rect 21315 42653 21327 42687
rect 21269 42647 21327 42653
rect 21376 42656 21680 42684
rect 17604 42616 17632 42644
rect 18785 42643 18843 42644
rect 14792 42588 15792 42616
rect 17144 42588 17632 42616
rect 14792 42576 14798 42588
rect 12069 42551 12127 42557
rect 12069 42517 12081 42551
rect 12115 42517 12127 42551
rect 12069 42511 12127 42517
rect 12158 42508 12164 42560
rect 12216 42548 12222 42560
rect 12897 42551 12955 42557
rect 12897 42548 12909 42551
rect 12216 42520 12909 42548
rect 12216 42508 12222 42520
rect 12897 42517 12909 42520
rect 12943 42517 12955 42551
rect 12897 42511 12955 42517
rect 13446 42508 13452 42560
rect 13504 42548 13510 42560
rect 14277 42551 14335 42557
rect 14277 42548 14289 42551
rect 13504 42520 14289 42548
rect 13504 42508 13510 42520
rect 14277 42517 14289 42520
rect 14323 42517 14335 42551
rect 14277 42511 14335 42517
rect 14550 42508 14556 42560
rect 14608 42508 14614 42560
rect 14826 42508 14832 42560
rect 14884 42508 14890 42560
rect 15470 42508 15476 42560
rect 15528 42508 15534 42560
rect 15764 42557 15792 42588
rect 19242 42576 19248 42628
rect 19300 42576 19306 42628
rect 20806 42616 20812 42628
rect 20456 42588 20812 42616
rect 15749 42551 15807 42557
rect 15749 42517 15761 42551
rect 15795 42517 15807 42551
rect 15749 42511 15807 42517
rect 15838 42508 15844 42560
rect 15896 42548 15902 42560
rect 16301 42551 16359 42557
rect 16301 42548 16313 42551
rect 15896 42520 16313 42548
rect 15896 42508 15902 42520
rect 16301 42517 16313 42520
rect 16347 42517 16359 42551
rect 16301 42511 16359 42517
rect 16758 42508 16764 42560
rect 16816 42508 16822 42560
rect 16942 42508 16948 42560
rect 17000 42508 17006 42560
rect 17218 42508 17224 42560
rect 17276 42508 17282 42560
rect 17310 42508 17316 42560
rect 17368 42548 17374 42560
rect 17497 42551 17555 42557
rect 17497 42548 17509 42551
rect 17368 42520 17509 42548
rect 17368 42508 17374 42520
rect 17497 42517 17509 42520
rect 17543 42517 17555 42551
rect 17497 42511 17555 42517
rect 17770 42508 17776 42560
rect 17828 42508 17834 42560
rect 18046 42508 18052 42560
rect 18104 42508 18110 42560
rect 18322 42508 18328 42560
rect 18380 42508 18386 42560
rect 18598 42508 18604 42560
rect 18656 42508 18662 42560
rect 18966 42508 18972 42560
rect 19024 42548 19030 42560
rect 20456 42548 20484 42588
rect 20806 42576 20812 42588
rect 20864 42576 20870 42628
rect 21082 42576 21088 42628
rect 21140 42616 21146 42628
rect 21376 42616 21404 42656
rect 21140 42588 21404 42616
rect 21140 42576 21146 42588
rect 21542 42576 21548 42628
rect 21600 42576 21606 42628
rect 21652 42616 21680 42656
rect 21910 42644 21916 42696
rect 21968 42644 21974 42696
rect 22066 42684 22094 42792
rect 22370 42780 22376 42832
rect 22428 42820 22434 42832
rect 23014 42820 23020 42832
rect 22428 42792 23020 42820
rect 22428 42780 22434 42792
rect 23014 42780 23020 42792
rect 23072 42780 23078 42832
rect 22278 42712 22284 42764
rect 22336 42752 22342 42764
rect 22925 42755 22983 42761
rect 22925 42752 22937 42755
rect 22336 42724 22937 42752
rect 22336 42712 22342 42724
rect 22925 42721 22937 42724
rect 22971 42721 22983 42755
rect 22925 42715 22983 42721
rect 23477 42755 23535 42761
rect 23477 42721 23489 42755
rect 23523 42752 23535 42755
rect 25130 42752 25136 42764
rect 23523 42724 25136 42752
rect 23523 42721 23535 42724
rect 23477 42715 23535 42721
rect 25130 42712 25136 42724
rect 25188 42712 25194 42764
rect 22465 42687 22523 42693
rect 22066 42656 22232 42684
rect 22097 42619 22155 42625
rect 21652 42588 22048 42616
rect 19024 42520 20484 42548
rect 19024 42508 19030 42520
rect 20530 42508 20536 42560
rect 20588 42508 20594 42560
rect 20990 42508 20996 42560
rect 21048 42548 21054 42560
rect 21910 42548 21916 42560
rect 21048 42520 21916 42548
rect 21048 42508 21054 42520
rect 21910 42508 21916 42520
rect 21968 42508 21974 42560
rect 22020 42548 22048 42588
rect 22097 42585 22109 42619
rect 22143 42585 22155 42619
rect 22204 42616 22232 42656
rect 22465 42653 22477 42687
rect 22511 42684 22523 42687
rect 24121 42687 24179 42693
rect 22511 42656 23888 42684
rect 22511 42653 22523 42656
rect 22465 42647 22523 42653
rect 22649 42619 22707 42625
rect 22649 42616 22661 42619
rect 22204 42588 22661 42616
rect 22097 42579 22155 42585
rect 22649 42585 22661 42588
rect 22695 42585 22707 42619
rect 22649 42579 22707 42585
rect 23201 42619 23259 42625
rect 23201 42585 23213 42619
rect 23247 42585 23259 42619
rect 23201 42579 23259 42585
rect 22112 42548 22140 42579
rect 22020 42520 22140 42548
rect 22186 42508 22192 42560
rect 22244 42548 22250 42560
rect 23216 42548 23244 42579
rect 23750 42576 23756 42628
rect 23808 42576 23814 42628
rect 23860 42616 23888 42656
rect 24121 42653 24133 42687
rect 24167 42684 24179 42687
rect 24210 42684 24216 42696
rect 24167 42656 24216 42684
rect 24167 42653 24179 42656
rect 24121 42647 24179 42653
rect 24210 42644 24216 42656
rect 24268 42644 24274 42696
rect 24578 42644 24584 42696
rect 24636 42644 24642 42696
rect 24596 42616 24624 42644
rect 23860 42588 24624 42616
rect 22244 42520 23244 42548
rect 22244 42508 22250 42520
rect 1104 42458 25000 42480
rect 1104 42406 6884 42458
rect 6936 42406 6948 42458
rect 7000 42406 7012 42458
rect 7064 42406 7076 42458
rect 7128 42406 7140 42458
rect 7192 42406 12818 42458
rect 12870 42406 12882 42458
rect 12934 42406 12946 42458
rect 12998 42406 13010 42458
rect 13062 42406 13074 42458
rect 13126 42406 18752 42458
rect 18804 42406 18816 42458
rect 18868 42406 18880 42458
rect 18932 42406 18944 42458
rect 18996 42406 19008 42458
rect 19060 42406 24686 42458
rect 24738 42406 24750 42458
rect 24802 42406 24814 42458
rect 24866 42406 24878 42458
rect 24930 42406 24942 42458
rect 24994 42406 25000 42458
rect 1104 42384 25000 42406
rect 474 42304 480 42356
rect 532 42344 538 42356
rect 1581 42347 1639 42353
rect 1581 42344 1593 42347
rect 532 42316 1593 42344
rect 532 42304 538 42316
rect 1581 42313 1593 42316
rect 1627 42313 1639 42347
rect 1581 42307 1639 42313
rect 1762 42304 1768 42356
rect 1820 42344 1826 42356
rect 2501 42347 2559 42353
rect 2501 42344 2513 42347
rect 1820 42316 2513 42344
rect 1820 42304 1826 42316
rect 2501 42313 2513 42316
rect 2547 42313 2559 42347
rect 2501 42307 2559 42313
rect 3234 42304 3240 42356
rect 3292 42344 3298 42356
rect 3421 42347 3479 42353
rect 3421 42344 3433 42347
rect 3292 42316 3433 42344
rect 3292 42304 3298 42316
rect 3421 42313 3433 42316
rect 3467 42313 3479 42347
rect 3421 42307 3479 42313
rect 3602 42304 3608 42356
rect 3660 42304 3666 42356
rect 3697 42347 3755 42353
rect 3697 42313 3709 42347
rect 3743 42313 3755 42347
rect 3697 42307 3755 42313
rect 1489 42279 1547 42285
rect 1489 42245 1501 42279
rect 1535 42276 1547 42279
rect 1535 42248 3188 42276
rect 1535 42245 1547 42248
rect 1489 42239 1547 42245
rect 2041 42211 2099 42217
rect 2041 42177 2053 42211
rect 2087 42177 2099 42211
rect 2041 42171 2099 42177
rect 2056 42140 2084 42171
rect 2406 42168 2412 42220
rect 2464 42208 2470 42220
rect 2685 42211 2743 42217
rect 2685 42208 2697 42211
rect 2464 42180 2697 42208
rect 2464 42168 2470 42180
rect 2685 42177 2697 42180
rect 2731 42177 2743 42211
rect 2685 42171 2743 42177
rect 2774 42168 2780 42220
rect 2832 42168 2838 42220
rect 3160 42152 3188 42248
rect 3620 42217 3648 42304
rect 3712 42276 3740 42307
rect 3786 42304 3792 42356
rect 3844 42344 3850 42356
rect 4157 42347 4215 42353
rect 4157 42344 4169 42347
rect 3844 42316 4169 42344
rect 3844 42304 3850 42316
rect 4157 42313 4169 42316
rect 4203 42313 4215 42347
rect 4985 42347 5043 42353
rect 4157 42307 4215 42313
rect 4356 42316 4844 42344
rect 4356 42276 4384 42316
rect 3712 42248 4384 42276
rect 3605 42211 3663 42217
rect 3605 42177 3617 42211
rect 3651 42177 3663 42211
rect 3605 42171 3663 42177
rect 3878 42168 3884 42220
rect 3936 42168 3942 42220
rect 3973 42211 4031 42217
rect 3973 42177 3985 42211
rect 4019 42177 4031 42211
rect 3973 42171 4031 42177
rect 2056 42112 2912 42140
rect 1210 41964 1216 42016
rect 1268 42004 1274 42016
rect 2133 42007 2191 42013
rect 2133 42004 2145 42007
rect 1268 41976 2145 42004
rect 1268 41964 1274 41976
rect 2133 41973 2145 41976
rect 2179 41973 2191 42007
rect 2884 42004 2912 42112
rect 3142 42100 3148 42152
rect 3200 42100 3206 42152
rect 2961 42075 3019 42081
rect 2961 42041 2973 42075
rect 3007 42072 3019 42075
rect 3510 42072 3516 42084
rect 3007 42044 3516 42072
rect 3007 42041 3019 42044
rect 2961 42035 3019 42041
rect 3510 42032 3516 42044
rect 3568 42032 3574 42084
rect 3602 42032 3608 42084
rect 3660 42072 3666 42084
rect 3994 42072 4022 42171
rect 4706 42168 4712 42220
rect 4764 42168 4770 42220
rect 4816 42217 4844 42316
rect 4985 42313 4997 42347
rect 5031 42344 5043 42347
rect 5166 42344 5172 42356
rect 5031 42316 5172 42344
rect 5031 42313 5043 42316
rect 4985 42307 5043 42313
rect 5166 42304 5172 42316
rect 5224 42304 5230 42356
rect 5997 42347 6055 42353
rect 5997 42313 6009 42347
rect 6043 42344 6055 42347
rect 6270 42344 6276 42356
rect 6043 42316 6276 42344
rect 6043 42313 6055 42316
rect 5997 42307 6055 42313
rect 6270 42304 6276 42316
rect 6328 42304 6334 42356
rect 7006 42304 7012 42356
rect 7064 42344 7070 42356
rect 7374 42344 7380 42356
rect 7064 42316 7380 42344
rect 7064 42304 7070 42316
rect 7374 42304 7380 42316
rect 7432 42304 7438 42356
rect 8202 42304 8208 42356
rect 8260 42344 8266 42356
rect 8481 42347 8539 42353
rect 8481 42344 8493 42347
rect 8260 42316 8493 42344
rect 8260 42304 8266 42316
rect 8481 42313 8493 42316
rect 8527 42313 8539 42347
rect 8481 42307 8539 42313
rect 8570 42304 8576 42356
rect 8628 42344 8634 42356
rect 8941 42347 8999 42353
rect 8941 42344 8953 42347
rect 8628 42316 8953 42344
rect 8628 42304 8634 42316
rect 8941 42313 8953 42316
rect 8987 42313 8999 42347
rect 8941 42307 8999 42313
rect 9122 42304 9128 42356
rect 9180 42344 9186 42356
rect 9217 42347 9275 42353
rect 9217 42344 9229 42347
rect 9180 42316 9229 42344
rect 9180 42304 9186 42316
rect 9217 42313 9229 42316
rect 9263 42313 9275 42347
rect 9217 42307 9275 42313
rect 9490 42304 9496 42356
rect 9548 42344 9554 42356
rect 9677 42347 9735 42353
rect 9677 42344 9689 42347
rect 9548 42316 9689 42344
rect 9548 42304 9554 42316
rect 9677 42313 9689 42316
rect 9723 42313 9735 42347
rect 9677 42307 9735 42313
rect 9950 42304 9956 42356
rect 10008 42304 10014 42356
rect 15470 42344 15476 42356
rect 12406 42316 15476 42344
rect 12406 42276 12434 42316
rect 15470 42304 15476 42316
rect 15528 42304 15534 42356
rect 17218 42344 17224 42356
rect 16776 42316 17224 42344
rect 5368 42248 9536 42276
rect 4801 42211 4859 42217
rect 4801 42177 4813 42211
rect 4847 42177 4859 42211
rect 4801 42171 4859 42177
rect 3660 42044 4022 42072
rect 4525 42075 4583 42081
rect 3660 42032 3666 42044
rect 4525 42041 4537 42075
rect 4571 42072 4583 42075
rect 5074 42072 5080 42084
rect 4571 42044 5080 42072
rect 4571 42041 4583 42044
rect 4525 42035 4583 42041
rect 5074 42032 5080 42044
rect 5132 42032 5138 42084
rect 5368 42004 5396 42248
rect 5445 42211 5503 42217
rect 5445 42177 5457 42211
rect 5491 42208 5503 42211
rect 5718 42208 5724 42220
rect 5491 42180 5724 42208
rect 5491 42177 5503 42180
rect 5445 42171 5503 42177
rect 5718 42168 5724 42180
rect 5776 42208 5782 42220
rect 5905 42211 5963 42217
rect 5905 42208 5917 42211
rect 5776 42180 5917 42208
rect 5776 42168 5782 42180
rect 5905 42177 5917 42180
rect 5951 42177 5963 42211
rect 5905 42171 5963 42177
rect 6178 42168 6184 42220
rect 6236 42168 6242 42220
rect 6546 42168 6552 42220
rect 6604 42168 6610 42220
rect 7101 42211 7159 42217
rect 7101 42177 7113 42211
rect 7147 42208 7159 42211
rect 7147 42180 7236 42208
rect 7147 42177 7159 42180
rect 7101 42171 7159 42177
rect 7208 42152 7236 42180
rect 7374 42168 7380 42220
rect 7432 42168 7438 42220
rect 7650 42168 7656 42220
rect 7708 42168 7714 42220
rect 7926 42168 7932 42220
rect 7984 42168 7990 42220
rect 8202 42168 8208 42220
rect 8260 42168 8266 42220
rect 8389 42211 8447 42217
rect 8389 42177 8401 42211
rect 8435 42177 8447 42211
rect 8389 42171 8447 42177
rect 7190 42100 7196 42152
rect 7248 42100 7254 42152
rect 7834 42100 7840 42152
rect 7892 42140 7898 42152
rect 8404 42140 8432 42171
rect 9122 42168 9128 42220
rect 9180 42168 9186 42220
rect 9398 42168 9404 42220
rect 9456 42168 9462 42220
rect 9508 42208 9536 42248
rect 9646 42248 12434 42276
rect 9646 42208 9674 42248
rect 13630 42236 13636 42288
rect 13688 42276 13694 42288
rect 15838 42276 15844 42288
rect 13688 42248 15844 42276
rect 13688 42236 13694 42248
rect 15838 42236 15844 42248
rect 15896 42236 15902 42288
rect 16776 42285 16804 42316
rect 17218 42304 17224 42316
rect 17276 42304 17282 42356
rect 17310 42304 17316 42356
rect 17368 42304 17374 42356
rect 17770 42304 17776 42356
rect 17828 42304 17834 42356
rect 18046 42304 18052 42356
rect 18104 42304 18110 42356
rect 18322 42344 18328 42356
rect 18248 42316 18328 42344
rect 16761 42279 16819 42285
rect 16761 42245 16773 42279
rect 16807 42245 16819 42279
rect 16761 42239 16819 42245
rect 16942 42236 16948 42288
rect 17000 42236 17006 42288
rect 17129 42279 17187 42285
rect 17129 42245 17141 42279
rect 17175 42276 17187 42279
rect 17328 42276 17356 42304
rect 17175 42248 17356 42276
rect 17497 42279 17555 42285
rect 17175 42245 17187 42248
rect 17129 42239 17187 42245
rect 17497 42245 17509 42279
rect 17543 42276 17555 42279
rect 17788 42276 17816 42304
rect 17543 42248 17816 42276
rect 17865 42279 17923 42285
rect 17543 42245 17555 42248
rect 17497 42239 17555 42245
rect 17865 42245 17877 42279
rect 17911 42276 17923 42279
rect 18064 42276 18092 42304
rect 17911 42248 18092 42276
rect 17911 42245 17923 42248
rect 17865 42239 17923 42245
rect 18138 42236 18144 42288
rect 18196 42236 18202 42288
rect 18248 42285 18276 42316
rect 18322 42304 18328 42316
rect 18380 42304 18386 42356
rect 19058 42304 19064 42356
rect 19116 42344 19122 42356
rect 19426 42344 19432 42356
rect 19116 42316 19432 42344
rect 19116 42304 19122 42316
rect 19426 42304 19432 42316
rect 19484 42304 19490 42356
rect 19705 42347 19763 42353
rect 19705 42313 19717 42347
rect 19751 42313 19763 42347
rect 19705 42307 19763 42313
rect 19981 42347 20039 42353
rect 19981 42313 19993 42347
rect 20027 42344 20039 42347
rect 20027 42316 20484 42344
rect 20027 42313 20039 42316
rect 19981 42307 20039 42313
rect 18233 42279 18291 42285
rect 18233 42245 18245 42279
rect 18279 42245 18291 42279
rect 18233 42239 18291 42245
rect 18598 42236 18604 42288
rect 18656 42236 18662 42288
rect 18969 42279 19027 42285
rect 18969 42276 18981 42279
rect 18800 42248 18981 42276
rect 9508 42180 9674 42208
rect 9858 42168 9864 42220
rect 9916 42168 9922 42220
rect 10137 42211 10195 42217
rect 10137 42177 10149 42211
rect 10183 42177 10195 42211
rect 12158 42208 12164 42220
rect 10137 42171 10195 42177
rect 10244 42180 12164 42208
rect 7892 42112 8432 42140
rect 7892 42100 7898 42112
rect 9490 42100 9496 42152
rect 9548 42140 9554 42152
rect 10152 42140 10180 42171
rect 9548 42112 10180 42140
rect 9548 42100 9554 42112
rect 5626 42032 5632 42084
rect 5684 42072 5690 42084
rect 6365 42075 6423 42081
rect 6365 42072 6377 42075
rect 5684 42044 6377 42072
rect 5684 42032 5690 42044
rect 6365 42041 6377 42044
rect 6411 42041 6423 42075
rect 6365 42035 6423 42041
rect 6454 42032 6460 42084
rect 6512 42072 6518 42084
rect 6512 42044 8156 42072
rect 6512 42032 6518 42044
rect 2884 41976 5396 42004
rect 2133 41967 2191 41973
rect 5718 41964 5724 42016
rect 5776 41964 5782 42016
rect 6914 41964 6920 42016
rect 6972 41964 6978 42016
rect 7193 42007 7251 42013
rect 7193 41973 7205 42007
rect 7239 42004 7251 42007
rect 7374 42004 7380 42016
rect 7239 41976 7380 42004
rect 7239 41973 7251 41976
rect 7193 41967 7251 41973
rect 7374 41964 7380 41976
rect 7432 41964 7438 42016
rect 7466 41964 7472 42016
rect 7524 41964 7530 42016
rect 7742 41964 7748 42016
rect 7800 41964 7806 42016
rect 8018 41964 8024 42016
rect 8076 41964 8082 42016
rect 8128 42004 8156 42044
rect 8294 42032 8300 42084
rect 8352 42072 8358 42084
rect 10244 42072 10272 42180
rect 12158 42168 12164 42180
rect 12216 42168 12222 42220
rect 16209 42211 16267 42217
rect 16209 42177 16221 42211
rect 16255 42208 16267 42211
rect 16960 42208 16988 42236
rect 16255 42180 16988 42208
rect 18156 42208 18184 42236
rect 18800 42208 18828 42248
rect 18969 42245 18981 42248
rect 19015 42245 19027 42279
rect 18969 42239 19027 42245
rect 19337 42279 19395 42285
rect 19337 42245 19349 42279
rect 19383 42276 19395 42279
rect 19518 42276 19524 42288
rect 19383 42248 19524 42276
rect 19383 42245 19395 42248
rect 19337 42239 19395 42245
rect 19518 42236 19524 42248
rect 19576 42236 19582 42288
rect 19720 42276 19748 42307
rect 19720 42248 20208 42276
rect 18156 42180 18828 42208
rect 16255 42177 16267 42180
rect 16209 42171 16267 42177
rect 18874 42168 18880 42220
rect 18932 42208 18938 42220
rect 20180 42217 20208 42248
rect 20456 42217 20484 42316
rect 20806 42304 20812 42356
rect 20864 42304 20870 42356
rect 21634 42304 21640 42356
rect 21692 42344 21698 42356
rect 21821 42347 21879 42353
rect 21821 42344 21833 42347
rect 21692 42316 21833 42344
rect 21692 42304 21698 42316
rect 21821 42313 21833 42316
rect 21867 42313 21879 42347
rect 21821 42307 21879 42313
rect 22830 42304 22836 42356
rect 22888 42304 22894 42356
rect 23109 42347 23167 42353
rect 23109 42313 23121 42347
rect 23155 42344 23167 42347
rect 23198 42344 23204 42356
rect 23155 42316 23204 42344
rect 23155 42313 23167 42316
rect 23109 42307 23167 42313
rect 23198 42304 23204 42316
rect 23256 42304 23262 42356
rect 23661 42347 23719 42353
rect 23661 42313 23673 42347
rect 23707 42344 23719 42347
rect 24486 42344 24492 42356
rect 23707 42316 24492 42344
rect 23707 42313 23719 42316
rect 23661 42307 23719 42313
rect 24486 42304 24492 42316
rect 24544 42304 24550 42356
rect 22848 42276 22876 42304
rect 24578 42276 24584 42288
rect 21652 42248 22876 42276
rect 23400 42248 24584 42276
rect 19889 42211 19947 42217
rect 19889 42208 19901 42211
rect 18932 42180 19901 42208
rect 18932 42168 18938 42180
rect 19889 42177 19901 42180
rect 19935 42177 19947 42211
rect 19889 42171 19947 42177
rect 20165 42211 20223 42217
rect 20165 42177 20177 42211
rect 20211 42177 20223 42211
rect 20165 42171 20223 42177
rect 20441 42211 20499 42217
rect 20441 42177 20453 42211
rect 20487 42177 20499 42211
rect 20441 42171 20499 42177
rect 20717 42211 20775 42217
rect 20717 42177 20729 42211
rect 20763 42177 20775 42211
rect 20717 42171 20775 42177
rect 18064 42112 20208 42140
rect 8352 42044 10272 42072
rect 8352 42032 8358 42044
rect 15286 42032 15292 42084
rect 15344 42072 15350 42084
rect 16114 42072 16120 42084
rect 15344 42044 16120 42072
rect 15344 42032 15350 42044
rect 16114 42032 16120 42044
rect 16172 42032 16178 42084
rect 16390 42032 16396 42084
rect 16448 42032 16454 42084
rect 17310 42032 17316 42084
rect 17368 42032 17374 42084
rect 18064 42081 18092 42112
rect 18049 42075 18107 42081
rect 18049 42041 18061 42075
rect 18095 42041 18107 42075
rect 18049 42035 18107 42041
rect 18414 42032 18420 42084
rect 18472 42032 18478 42084
rect 18966 42072 18972 42084
rect 18616 42044 18972 42072
rect 15194 42004 15200 42016
rect 8128 41976 15200 42004
rect 15194 41964 15200 41976
rect 15252 41964 15258 42016
rect 15378 41964 15384 42016
rect 15436 42004 15442 42016
rect 16482 42004 16488 42016
rect 15436 41976 16488 42004
rect 15436 41964 15442 41976
rect 16482 41964 16488 41976
rect 16540 41964 16546 42016
rect 16850 41964 16856 42016
rect 16908 41964 16914 42016
rect 17586 41964 17592 42016
rect 17644 41964 17650 42016
rect 18138 41964 18144 42016
rect 18196 42004 18202 42016
rect 18616 42004 18644 42044
rect 18966 42032 18972 42044
rect 19024 42032 19030 42084
rect 19886 42032 19892 42084
rect 19944 42032 19950 42084
rect 20180 42072 20208 42112
rect 20254 42100 20260 42152
rect 20312 42140 20318 42152
rect 20732 42140 20760 42171
rect 20806 42168 20812 42220
rect 20864 42208 20870 42220
rect 20993 42211 21051 42217
rect 20993 42208 21005 42211
rect 20864 42180 21005 42208
rect 20864 42168 20870 42180
rect 20993 42177 21005 42180
rect 21039 42177 21051 42211
rect 20993 42171 21051 42177
rect 21266 42168 21272 42220
rect 21324 42168 21330 42220
rect 21652 42217 21680 42248
rect 21637 42211 21695 42217
rect 21637 42177 21649 42211
rect 21683 42177 21695 42211
rect 21637 42171 21695 42177
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 20312 42112 20760 42140
rect 20312 42100 20318 42112
rect 20898 42100 20904 42152
rect 20956 42140 20962 42152
rect 22020 42140 22048 42171
rect 22186 42168 22192 42220
rect 22244 42168 22250 42220
rect 22281 42211 22339 42217
rect 22281 42177 22293 42211
rect 22327 42177 22339 42211
rect 22281 42171 22339 42177
rect 20956 42112 22048 42140
rect 20956 42100 20962 42112
rect 20180 42044 20392 42072
rect 18196 41976 18644 42004
rect 18196 41964 18202 41976
rect 18690 41964 18696 42016
rect 18748 41964 18754 42016
rect 18782 41964 18788 42016
rect 18840 42004 18846 42016
rect 19061 42007 19119 42013
rect 19061 42004 19073 42007
rect 18840 41976 19073 42004
rect 18840 41964 18846 41976
rect 19061 41973 19073 41976
rect 19107 41973 19119 42007
rect 19061 41967 19119 41973
rect 19426 41964 19432 42016
rect 19484 41964 19490 42016
rect 19904 42004 19932 42032
rect 20257 42007 20315 42013
rect 20257 42004 20269 42007
rect 19904 41976 20269 42004
rect 20257 41973 20269 41976
rect 20303 41973 20315 42007
rect 20364 42004 20392 42044
rect 20438 42032 20444 42084
rect 20496 42072 20502 42084
rect 20533 42075 20591 42081
rect 20533 42072 20545 42075
rect 20496 42044 20545 42072
rect 20496 42032 20502 42044
rect 20533 42041 20545 42044
rect 20579 42041 20591 42075
rect 21910 42072 21916 42084
rect 20533 42035 20591 42041
rect 20732 42044 21916 42072
rect 20732 42004 20760 42044
rect 21910 42032 21916 42044
rect 21968 42032 21974 42084
rect 22002 42032 22008 42084
rect 22060 42072 22066 42084
rect 22204 42072 22232 42168
rect 22060 42044 22232 42072
rect 22296 42072 22324 42171
rect 22830 42168 22836 42220
rect 22888 42168 22894 42220
rect 23400 42217 23428 42248
rect 24578 42236 24584 42248
rect 24636 42236 24642 42288
rect 23385 42211 23443 42217
rect 23385 42177 23397 42211
rect 23431 42177 23443 42211
rect 23385 42171 23443 42177
rect 24026 42168 24032 42220
rect 24084 42168 24090 42220
rect 22557 42143 22615 42149
rect 22557 42109 22569 42143
rect 22603 42140 22615 42143
rect 25590 42140 25596 42152
rect 22603 42112 25596 42140
rect 22603 42109 22615 42112
rect 22557 42103 22615 42109
rect 25590 42100 25596 42112
rect 25648 42100 25654 42152
rect 24210 42072 24216 42084
rect 22296 42044 24216 42072
rect 22060 42032 22066 42044
rect 24210 42032 24216 42044
rect 24268 42032 24274 42084
rect 20364 41976 20760 42004
rect 20257 41967 20315 41973
rect 21174 41964 21180 42016
rect 21232 42004 21238 42016
rect 23474 42004 23480 42016
rect 21232 41976 23480 42004
rect 21232 41964 21238 41976
rect 23474 41964 23480 41976
rect 23532 41964 23538 42016
rect 24305 42007 24363 42013
rect 24305 41973 24317 42007
rect 24351 42004 24363 42007
rect 25222 42004 25228 42016
rect 24351 41976 25228 42004
rect 24351 41973 24363 41976
rect 24305 41967 24363 41973
rect 25222 41964 25228 41976
rect 25280 41964 25286 42016
rect 1104 41914 24840 41936
rect 1104 41862 3917 41914
rect 3969 41862 3981 41914
rect 4033 41862 4045 41914
rect 4097 41862 4109 41914
rect 4161 41862 4173 41914
rect 4225 41862 9851 41914
rect 9903 41862 9915 41914
rect 9967 41862 9979 41914
rect 10031 41862 10043 41914
rect 10095 41862 10107 41914
rect 10159 41862 15785 41914
rect 15837 41862 15849 41914
rect 15901 41862 15913 41914
rect 15965 41862 15977 41914
rect 16029 41862 16041 41914
rect 16093 41862 21719 41914
rect 21771 41862 21783 41914
rect 21835 41862 21847 41914
rect 21899 41862 21911 41914
rect 21963 41862 21975 41914
rect 22027 41862 24840 41914
rect 1104 41840 24840 41862
rect 934 41760 940 41812
rect 992 41800 998 41812
rect 1581 41803 1639 41809
rect 1581 41800 1593 41803
rect 992 41772 1593 41800
rect 992 41760 998 41772
rect 1581 41769 1593 41772
rect 1627 41769 1639 41803
rect 1581 41763 1639 41769
rect 2590 41760 2596 41812
rect 2648 41800 2654 41812
rect 2685 41803 2743 41809
rect 2685 41800 2697 41803
rect 2648 41772 2697 41800
rect 2648 41760 2654 41772
rect 2685 41769 2697 41772
rect 2731 41769 2743 41803
rect 2685 41763 2743 41769
rect 2774 41760 2780 41812
rect 2832 41800 2838 41812
rect 2869 41803 2927 41809
rect 2869 41800 2881 41803
rect 2832 41772 2881 41800
rect 2832 41760 2838 41772
rect 2869 41769 2881 41772
rect 2915 41769 2927 41803
rect 2869 41763 2927 41769
rect 3145 41803 3203 41809
rect 3145 41769 3157 41803
rect 3191 41800 3203 41803
rect 3326 41800 3332 41812
rect 3191 41772 3332 41800
rect 3191 41769 3203 41772
rect 3145 41763 3203 41769
rect 3326 41760 3332 41772
rect 3384 41760 3390 41812
rect 3421 41803 3479 41809
rect 3421 41769 3433 41803
rect 3467 41800 3479 41803
rect 3602 41800 3608 41812
rect 3467 41772 3608 41800
rect 3467 41769 3479 41772
rect 3421 41763 3479 41769
rect 3602 41760 3608 41772
rect 3660 41760 3666 41812
rect 3789 41803 3847 41809
rect 3789 41769 3801 41803
rect 3835 41800 3847 41803
rect 4246 41800 4252 41812
rect 3835 41772 4252 41800
rect 3835 41769 3847 41772
rect 3789 41763 3847 41769
rect 4246 41760 4252 41772
rect 4304 41760 4310 41812
rect 4430 41760 4436 41812
rect 4488 41760 4494 41812
rect 4709 41803 4767 41809
rect 4709 41769 4721 41803
rect 4755 41800 4767 41803
rect 5258 41800 5264 41812
rect 4755 41772 5264 41800
rect 4755 41769 4767 41772
rect 4709 41763 4767 41769
rect 5258 41760 5264 41772
rect 5316 41760 5322 41812
rect 5445 41803 5503 41809
rect 5445 41769 5457 41803
rect 5491 41800 5503 41803
rect 5534 41800 5540 41812
rect 5491 41772 5540 41800
rect 5491 41769 5503 41772
rect 5445 41763 5503 41769
rect 5534 41760 5540 41772
rect 5592 41760 5598 41812
rect 5813 41803 5871 41809
rect 5813 41769 5825 41803
rect 5859 41800 5871 41803
rect 5902 41800 5908 41812
rect 5859 41772 5908 41800
rect 5859 41769 5871 41772
rect 5813 41763 5871 41769
rect 5902 41760 5908 41772
rect 5960 41760 5966 41812
rect 5994 41760 6000 41812
rect 6052 41800 6058 41812
rect 6181 41803 6239 41809
rect 6181 41800 6193 41803
rect 6052 41772 6193 41800
rect 6052 41760 6058 41772
rect 6181 41769 6193 41772
rect 6227 41769 6239 41803
rect 6181 41763 6239 41769
rect 6914 41760 6920 41812
rect 6972 41760 6978 41812
rect 7193 41803 7251 41809
rect 7193 41769 7205 41803
rect 7239 41800 7251 41803
rect 7282 41800 7288 41812
rect 7239 41772 7288 41800
rect 7239 41769 7251 41772
rect 7193 41763 7251 41769
rect 7282 41760 7288 41772
rect 7340 41760 7346 41812
rect 7374 41760 7380 41812
rect 7432 41760 7438 41812
rect 7466 41760 7472 41812
rect 7524 41760 7530 41812
rect 7558 41760 7564 41812
rect 7616 41760 7622 41812
rect 7742 41760 7748 41812
rect 7800 41800 7806 41812
rect 8389 41803 8447 41809
rect 7800 41772 8340 41800
rect 7800 41760 7806 41772
rect 3786 41624 3792 41676
rect 3844 41664 3850 41676
rect 4982 41664 4988 41676
rect 3844 41636 4988 41664
rect 3844 41624 3850 41636
rect 4982 41624 4988 41636
rect 5040 41624 5046 41676
rect 5074 41624 5080 41676
rect 5132 41664 5138 41676
rect 5132 41636 6408 41664
rect 5132 41624 5138 41636
rect 1486 41556 1492 41608
rect 1544 41556 1550 41608
rect 2501 41599 2559 41605
rect 2501 41565 2513 41599
rect 2547 41565 2559 41599
rect 2501 41559 2559 41565
rect 3053 41599 3111 41605
rect 3053 41565 3065 41599
rect 3099 41565 3111 41599
rect 3053 41559 3111 41565
rect 1670 41488 1676 41540
rect 1728 41528 1734 41540
rect 2041 41531 2099 41537
rect 2041 41528 2053 41531
rect 1728 41500 2053 41528
rect 1728 41488 1734 41500
rect 2041 41497 2053 41500
rect 2087 41497 2099 41531
rect 2041 41491 2099 41497
rect 2314 41488 2320 41540
rect 2372 41488 2378 41540
rect 2516 41528 2544 41559
rect 2958 41528 2964 41540
rect 2516 41500 2964 41528
rect 2958 41488 2964 41500
rect 3016 41488 3022 41540
rect 3068 41528 3096 41559
rect 3326 41556 3332 41608
rect 3384 41556 3390 41608
rect 3602 41556 3608 41608
rect 3660 41556 3666 41608
rect 3694 41556 3700 41608
rect 3752 41596 3758 41608
rect 3973 41599 4031 41605
rect 3973 41596 3985 41599
rect 3752 41568 3985 41596
rect 3752 41556 3758 41568
rect 3973 41565 3985 41568
rect 4019 41565 4031 41599
rect 3973 41559 4031 41565
rect 4246 41556 4252 41608
rect 4304 41556 4310 41608
rect 4614 41556 4620 41608
rect 4672 41556 4678 41608
rect 4893 41599 4951 41605
rect 4893 41565 4905 41599
rect 4939 41565 4951 41599
rect 4893 41559 4951 41565
rect 5353 41599 5411 41605
rect 5353 41565 5365 41599
rect 5399 41565 5411 41599
rect 5353 41559 5411 41565
rect 3418 41528 3424 41540
rect 3068 41500 3424 41528
rect 3418 41488 3424 41500
rect 3476 41488 3482 41540
rect 4154 41488 4160 41540
rect 4212 41528 4218 41540
rect 4908 41528 4936 41559
rect 4212 41500 4936 41528
rect 5368 41528 5396 41559
rect 5626 41556 5632 41608
rect 5684 41556 5690 41608
rect 5718 41556 5724 41608
rect 5776 41596 5782 41608
rect 6380 41605 6408 41636
rect 5997 41599 6055 41605
rect 5997 41596 6009 41599
rect 5776 41568 6009 41596
rect 5776 41556 5782 41568
rect 5997 41565 6009 41568
rect 6043 41565 6055 41599
rect 5997 41559 6055 41565
rect 6365 41599 6423 41605
rect 6365 41565 6377 41599
rect 6411 41565 6423 41599
rect 6365 41559 6423 41565
rect 6730 41556 6736 41608
rect 6788 41556 6794 41608
rect 6932 41596 6960 41760
rect 7392 41664 7420 41760
rect 7484 41732 7512 41760
rect 7484 41704 8064 41732
rect 7392 41636 7788 41664
rect 7760 41605 7788 41636
rect 8036 41605 8064 41704
rect 8110 41692 8116 41744
rect 8168 41692 8174 41744
rect 8312 41605 8340 41772
rect 8389 41769 8401 41803
rect 8435 41800 8447 41803
rect 8478 41800 8484 41812
rect 8435 41772 8484 41800
rect 8435 41769 8447 41772
rect 8389 41763 8447 41769
rect 8478 41760 8484 41772
rect 8536 41760 8542 41812
rect 10042 41800 10048 41812
rect 9692 41772 10048 41800
rect 9692 41673 9720 41772
rect 10042 41760 10048 41772
rect 10100 41800 10106 41812
rect 10100 41772 16160 41800
rect 10100 41760 10106 41772
rect 16132 41732 16160 41772
rect 17954 41760 17960 41812
rect 18012 41760 18018 41812
rect 18046 41760 18052 41812
rect 18104 41800 18110 41812
rect 18417 41803 18475 41809
rect 18417 41800 18429 41803
rect 18104 41772 18429 41800
rect 18104 41760 18110 41772
rect 18417 41769 18429 41772
rect 18463 41769 18475 41803
rect 18417 41763 18475 41769
rect 18506 41760 18512 41812
rect 18564 41800 18570 41812
rect 18785 41803 18843 41809
rect 18785 41800 18797 41803
rect 18564 41772 18797 41800
rect 18564 41760 18570 41772
rect 18785 41769 18797 41772
rect 18831 41769 18843 41803
rect 18785 41763 18843 41769
rect 18874 41760 18880 41812
rect 18932 41760 18938 41812
rect 19518 41760 19524 41812
rect 19576 41800 19582 41812
rect 19613 41803 19671 41809
rect 19613 41800 19625 41803
rect 19576 41772 19625 41800
rect 19576 41760 19582 41772
rect 19613 41769 19625 41772
rect 19659 41769 19671 41803
rect 19613 41763 19671 41769
rect 20254 41760 20260 41812
rect 20312 41760 20318 41812
rect 20530 41760 20536 41812
rect 20588 41800 20594 41812
rect 20588 41772 20668 41800
rect 20588 41760 20594 41772
rect 18892 41732 18920 41760
rect 16132 41704 18920 41732
rect 19337 41735 19395 41741
rect 19337 41701 19349 41735
rect 19383 41701 19395 41735
rect 19337 41695 19395 41701
rect 19981 41735 20039 41741
rect 19981 41701 19993 41735
rect 20027 41732 20039 41735
rect 20346 41732 20352 41744
rect 20027 41704 20352 41732
rect 20027 41701 20039 41704
rect 19981 41695 20039 41701
rect 9677 41667 9735 41673
rect 9677 41633 9689 41667
rect 9723 41633 9735 41667
rect 19352 41664 19380 41695
rect 20346 41692 20352 41704
rect 20404 41692 20410 41744
rect 20640 41664 20668 41772
rect 20714 41760 20720 41812
rect 20772 41760 20778 41812
rect 21174 41760 21180 41812
rect 21232 41760 21238 41812
rect 21358 41760 21364 41812
rect 21416 41800 21422 41812
rect 22278 41800 22284 41812
rect 21416 41772 22284 41800
rect 21416 41760 21422 41772
rect 22278 41760 22284 41772
rect 22336 41760 22342 41812
rect 23017 41803 23075 41809
rect 23017 41769 23029 41803
rect 23063 41800 23075 41803
rect 23934 41800 23940 41812
rect 23063 41772 23940 41800
rect 23063 41769 23075 41772
rect 23017 41763 23075 41769
rect 23934 41760 23940 41772
rect 23992 41760 23998 41812
rect 24121 41803 24179 41809
rect 24121 41769 24133 41803
rect 24167 41800 24179 41803
rect 25314 41800 25320 41812
rect 24167 41772 25320 41800
rect 24167 41769 24179 41772
rect 24121 41763 24179 41769
rect 25314 41760 25320 41772
rect 25372 41760 25378 41812
rect 25406 41760 25412 41812
rect 25464 41760 25470 41812
rect 23569 41735 23627 41741
rect 9677 41627 9735 41633
rect 12406 41636 19104 41664
rect 19352 41636 20208 41664
rect 7377 41599 7435 41605
rect 7377 41596 7389 41599
rect 6932 41568 7389 41596
rect 7377 41565 7389 41568
rect 7423 41565 7435 41599
rect 7377 41559 7435 41565
rect 7745 41599 7803 41605
rect 7745 41565 7757 41599
rect 7791 41565 7803 41599
rect 7745 41559 7803 41565
rect 8021 41599 8079 41605
rect 8021 41565 8033 41599
rect 8067 41565 8079 41599
rect 8021 41559 8079 41565
rect 8297 41599 8355 41605
rect 8297 41565 8309 41599
rect 8343 41565 8355 41599
rect 8297 41559 8355 41565
rect 8573 41599 8631 41605
rect 8573 41565 8585 41599
rect 8619 41596 8631 41599
rect 8846 41596 8852 41608
rect 8619 41568 8852 41596
rect 8619 41565 8631 41568
rect 8573 41559 8631 41565
rect 8846 41556 8852 41568
rect 8904 41556 8910 41608
rect 9951 41599 10009 41605
rect 9951 41565 9963 41599
rect 9997 41596 10009 41599
rect 10318 41596 10324 41608
rect 9997 41568 10324 41596
rect 9997 41565 10009 41568
rect 9951 41559 10009 41565
rect 10318 41556 10324 41568
rect 10376 41596 10382 41608
rect 12406 41596 12434 41636
rect 10376 41568 12434 41596
rect 10376 41556 10382 41568
rect 17954 41556 17960 41608
rect 18012 41596 18018 41608
rect 18012 41568 18092 41596
rect 18012 41556 18018 41568
rect 5368 41500 6592 41528
rect 4212 41488 4218 41500
rect 1578 41420 1584 41472
rect 1636 41460 1642 41472
rect 2133 41463 2191 41469
rect 2133 41460 2145 41463
rect 1636 41432 2145 41460
rect 1636 41420 1642 41432
rect 2133 41429 2145 41432
rect 2179 41429 2191 41463
rect 2332 41460 2360 41488
rect 4065 41463 4123 41469
rect 4065 41460 4077 41463
rect 2332 41432 4077 41460
rect 2133 41423 2191 41429
rect 4065 41429 4077 41432
rect 4111 41429 4123 41463
rect 4065 41423 4123 41429
rect 5169 41463 5227 41469
rect 5169 41429 5181 41463
rect 5215 41460 5227 41463
rect 6086 41460 6092 41472
rect 5215 41432 6092 41460
rect 5215 41429 5227 41432
rect 5169 41423 5227 41429
rect 6086 41420 6092 41432
rect 6144 41420 6150 41472
rect 6564 41469 6592 41500
rect 7006 41488 7012 41540
rect 7064 41528 7070 41540
rect 7064 41500 7880 41528
rect 7064 41488 7070 41500
rect 6549 41463 6607 41469
rect 6549 41429 6561 41463
rect 6595 41429 6607 41463
rect 6549 41423 6607 41429
rect 7101 41463 7159 41469
rect 7101 41429 7113 41463
rect 7147 41460 7159 41463
rect 7282 41460 7288 41472
rect 7147 41432 7288 41460
rect 7147 41429 7159 41432
rect 7101 41423 7159 41429
rect 7282 41420 7288 41432
rect 7340 41420 7346 41472
rect 7852 41469 7880 41500
rect 15470 41488 15476 41540
rect 15528 41528 15534 41540
rect 17770 41528 17776 41540
rect 15528 41500 17776 41528
rect 15528 41488 15534 41500
rect 17770 41488 17776 41500
rect 17828 41488 17834 41540
rect 18064 41528 18092 41568
rect 18138 41556 18144 41608
rect 18196 41556 18202 41608
rect 18230 41556 18236 41608
rect 18288 41596 18294 41608
rect 18325 41599 18383 41605
rect 18325 41596 18337 41599
rect 18288 41568 18337 41596
rect 18288 41556 18294 41568
rect 18325 41565 18337 41568
rect 18371 41565 18383 41599
rect 18325 41559 18383 41565
rect 18414 41556 18420 41608
rect 18472 41596 18478 41608
rect 18969 41599 19027 41605
rect 18969 41596 18981 41599
rect 18472 41568 18981 41596
rect 18472 41556 18478 41568
rect 18969 41565 18981 41568
rect 19015 41565 19027 41599
rect 19076 41596 19104 41636
rect 19521 41599 19579 41605
rect 19521 41596 19533 41599
rect 19076 41568 19533 41596
rect 18969 41559 19027 41565
rect 19521 41565 19533 41568
rect 19567 41565 19579 41599
rect 19521 41559 19579 41565
rect 19702 41556 19708 41608
rect 19760 41596 19766 41608
rect 20180 41605 20208 41636
rect 20548 41636 20668 41664
rect 21192 41704 23336 41732
rect 19797 41599 19855 41605
rect 19797 41596 19809 41599
rect 19760 41568 19809 41596
rect 19760 41556 19766 41568
rect 19797 41565 19809 41568
rect 19843 41565 19855 41599
rect 19797 41559 19855 41565
rect 20165 41599 20223 41605
rect 20165 41565 20177 41599
rect 20211 41565 20223 41599
rect 20165 41559 20223 41565
rect 20254 41556 20260 41608
rect 20312 41596 20318 41608
rect 20441 41599 20499 41605
rect 20548 41601 20576 41636
rect 21192 41608 21220 41704
rect 20441 41596 20453 41599
rect 20312 41568 20453 41596
rect 20312 41556 20318 41568
rect 20441 41565 20453 41568
rect 20487 41565 20499 41599
rect 20441 41559 20499 41565
rect 20533 41595 20591 41601
rect 21085 41599 21143 41605
rect 21085 41596 21097 41599
rect 20533 41561 20545 41595
rect 20579 41561 20591 41595
rect 20533 41555 20591 41561
rect 20640 41568 21097 41596
rect 19334 41528 19340 41540
rect 18064 41500 19340 41528
rect 19334 41488 19340 41500
rect 19392 41488 19398 41540
rect 7837 41463 7895 41469
rect 7837 41429 7849 41463
rect 7883 41429 7895 41463
rect 7837 41423 7895 41429
rect 10686 41420 10692 41472
rect 10744 41420 10750 41472
rect 15194 41420 15200 41472
rect 15252 41460 15258 41472
rect 20640 41460 20668 41568
rect 21085 41565 21097 41568
rect 21131 41565 21143 41599
rect 21085 41559 21143 41565
rect 21174 41556 21180 41608
rect 21232 41556 21238 41608
rect 21358 41556 21364 41608
rect 21416 41556 21422 41608
rect 21634 41556 21640 41608
rect 21692 41556 21698 41608
rect 23308 41605 23336 41704
rect 23569 41701 23581 41735
rect 23615 41732 23627 41735
rect 25424 41732 25452 41760
rect 23615 41704 25452 41732
rect 23615 41701 23627 41704
rect 23569 41695 23627 41701
rect 21913 41599 21971 41605
rect 21913 41596 21925 41599
rect 21744 41568 21925 41596
rect 21744 41528 21772 41568
rect 21913 41565 21925 41568
rect 21959 41565 21971 41599
rect 22741 41599 22799 41605
rect 22741 41596 22753 41599
rect 21913 41559 21971 41565
rect 22066 41568 22753 41596
rect 20916 41500 21772 41528
rect 20916 41469 20944 41500
rect 21818 41488 21824 41540
rect 21876 41528 21882 41540
rect 22066 41528 22094 41568
rect 22741 41565 22753 41568
rect 22787 41565 22799 41599
rect 22741 41559 22799 41565
rect 23293 41599 23351 41605
rect 23293 41565 23305 41599
rect 23339 41565 23351 41599
rect 23293 41559 23351 41565
rect 23566 41556 23572 41608
rect 23624 41596 23630 41608
rect 25774 41596 25780 41608
rect 23624 41568 25780 41596
rect 23624 41556 23630 41568
rect 25774 41556 25780 41568
rect 25832 41556 25838 41608
rect 21876 41500 22094 41528
rect 22189 41531 22247 41537
rect 21876 41488 21882 41500
rect 22189 41497 22201 41531
rect 22235 41528 22247 41531
rect 22235 41500 23796 41528
rect 22235 41497 22247 41500
rect 22189 41491 22247 41497
rect 15252 41432 20668 41460
rect 20901 41463 20959 41469
rect 15252 41420 15258 41432
rect 20901 41429 20913 41463
rect 20947 41429 20959 41463
rect 20901 41423 20959 41429
rect 21450 41420 21456 41472
rect 21508 41420 21514 41472
rect 21729 41463 21787 41469
rect 21729 41429 21741 41463
rect 21775 41460 21787 41463
rect 22370 41460 22376 41472
rect 21775 41432 22376 41460
rect 21775 41429 21787 41432
rect 21729 41423 21787 41429
rect 22370 41420 22376 41432
rect 22428 41420 22434 41472
rect 22465 41463 22523 41469
rect 22465 41429 22477 41463
rect 22511 41460 22523 41463
rect 23658 41460 23664 41472
rect 22511 41432 23664 41460
rect 22511 41429 22523 41432
rect 22465 41423 22523 41429
rect 23658 41420 23664 41432
rect 23716 41420 23722 41472
rect 23768 41460 23796 41500
rect 23842 41488 23848 41540
rect 23900 41488 23906 41540
rect 23934 41460 23940 41472
rect 23768 41432 23940 41460
rect 23934 41420 23940 41432
rect 23992 41420 23998 41472
rect 1104 41370 25000 41392
rect 1104 41318 6884 41370
rect 6936 41318 6948 41370
rect 7000 41318 7012 41370
rect 7064 41318 7076 41370
rect 7128 41318 7140 41370
rect 7192 41318 12818 41370
rect 12870 41318 12882 41370
rect 12934 41318 12946 41370
rect 12998 41318 13010 41370
rect 13062 41318 13074 41370
rect 13126 41318 18752 41370
rect 18804 41318 18816 41370
rect 18868 41318 18880 41370
rect 18932 41318 18944 41370
rect 18996 41318 19008 41370
rect 19060 41318 24686 41370
rect 24738 41318 24750 41370
rect 24802 41318 24814 41370
rect 24866 41318 24878 41370
rect 24930 41318 24942 41370
rect 24994 41318 25000 41370
rect 1104 41296 25000 41318
rect 2498 41216 2504 41268
rect 2556 41216 2562 41268
rect 2774 41216 2780 41268
rect 2832 41216 2838 41268
rect 2958 41216 2964 41268
rect 3016 41256 3022 41268
rect 3053 41259 3111 41265
rect 3053 41256 3065 41259
rect 3016 41228 3065 41256
rect 3016 41216 3022 41228
rect 3053 41225 3065 41228
rect 3099 41225 3111 41259
rect 3053 41219 3111 41225
rect 7745 41259 7803 41265
rect 7745 41225 7757 41259
rect 7791 41256 7803 41259
rect 7834 41256 7840 41268
rect 7791 41228 7840 41256
rect 7791 41225 7803 41228
rect 7745 41219 7803 41225
rect 7834 41216 7840 41228
rect 7892 41216 7898 41268
rect 15102 41256 15108 41268
rect 7944 41228 15108 41256
rect 2225 41191 2283 41197
rect 2225 41157 2237 41191
rect 2271 41188 2283 41191
rect 7944 41188 7972 41228
rect 15102 41216 15108 41228
rect 15160 41216 15166 41268
rect 19521 41259 19579 41265
rect 19521 41225 19533 41259
rect 19567 41225 19579 41259
rect 19521 41219 19579 41225
rect 20073 41259 20131 41265
rect 20073 41225 20085 41259
rect 20119 41256 20131 41259
rect 20254 41256 20260 41268
rect 20119 41228 20260 41256
rect 20119 41225 20131 41228
rect 20073 41219 20131 41225
rect 12526 41188 12532 41200
rect 2271 41160 7972 41188
rect 10244 41160 12532 41188
rect 2271 41157 2283 41160
rect 2225 41151 2283 41157
rect 8831 41153 8889 41159
rect 1394 41080 1400 41132
rect 1452 41080 1458 41132
rect 2685 41123 2743 41129
rect 2685 41089 2697 41123
rect 2731 41089 2743 41123
rect 2685 41083 2743 41089
rect 2961 41123 3019 41129
rect 2961 41089 2973 41123
rect 3007 41089 3019 41123
rect 2961 41083 3019 41089
rect 474 41012 480 41064
rect 532 41052 538 41064
rect 2700 41052 2728 41083
rect 532 41024 2728 41052
rect 532 41012 538 41024
rect 382 40944 388 40996
rect 440 40984 446 40996
rect 2976 40984 3004 41083
rect 3234 41080 3240 41132
rect 3292 41080 3298 41132
rect 3418 41080 3424 41132
rect 3476 41120 3482 41132
rect 3787 41123 3845 41129
rect 3787 41120 3799 41123
rect 3476 41092 3799 41120
rect 3476 41080 3482 41092
rect 3787 41089 3799 41092
rect 3833 41120 3845 41123
rect 5167 41123 5225 41129
rect 3833 41092 4844 41120
rect 3833 41089 3845 41092
rect 3787 41083 3845 41089
rect 3510 41012 3516 41064
rect 3568 41012 3574 41064
rect 440 40956 3004 40984
rect 440 40944 446 40956
rect 1026 40876 1032 40928
rect 1084 40916 1090 40928
rect 3326 40916 3332 40928
rect 1084 40888 3332 40916
rect 1084 40876 1090 40888
rect 3326 40876 3332 40888
rect 3384 40876 3390 40928
rect 4522 40876 4528 40928
rect 4580 40876 4586 40928
rect 4816 40916 4844 41092
rect 5167 41089 5179 41123
rect 5213 41120 5225 41123
rect 5258 41120 5264 41132
rect 5213 41092 5264 41120
rect 5213 41089 5225 41092
rect 5167 41083 5225 41089
rect 5258 41080 5264 41092
rect 5316 41080 5322 41132
rect 7926 41080 7932 41132
rect 7984 41080 7990 41132
rect 8831 41119 8843 41153
rect 8877 41150 8889 41153
rect 8877 41120 8892 41150
rect 10244 41120 10272 41160
rect 12526 41148 12532 41160
rect 12584 41148 12590 41200
rect 8877 41119 10272 41120
rect 8831 41113 10272 41119
rect 8864 41092 10272 41113
rect 10319 41123 10377 41129
rect 10319 41089 10331 41123
rect 10365 41120 10377 41123
rect 19245 41123 19303 41129
rect 10365 41092 10732 41120
rect 10365 41089 10377 41092
rect 10319 41083 10377 41089
rect 4890 41012 4896 41064
rect 4948 41012 4954 41064
rect 8570 41012 8576 41064
rect 8628 41012 8634 41064
rect 10042 41052 10048 41064
rect 9232 41024 10048 41052
rect 5810 40916 5816 40928
rect 4816 40888 5816 40916
rect 5810 40876 5816 40888
rect 5868 40876 5874 40928
rect 5905 40919 5963 40925
rect 5905 40885 5917 40919
rect 5951 40916 5963 40919
rect 5994 40916 6000 40928
rect 5951 40888 6000 40916
rect 5951 40885 5963 40888
rect 5905 40879 5963 40885
rect 5994 40876 6000 40888
rect 6052 40876 6058 40928
rect 8588 40916 8616 41012
rect 9232 40916 9260 41024
rect 10042 41012 10048 41024
rect 10100 41012 10106 41064
rect 10704 40984 10732 41092
rect 19245 41089 19257 41123
rect 19291 41120 19303 41123
rect 19536 41120 19564 41219
rect 20254 41216 20260 41228
rect 20312 41216 20318 41268
rect 20625 41259 20683 41265
rect 20625 41225 20637 41259
rect 20671 41225 20683 41259
rect 20625 41219 20683 41225
rect 20901 41259 20959 41265
rect 20901 41225 20913 41259
rect 20947 41256 20959 41259
rect 21082 41256 21088 41268
rect 20947 41228 21088 41256
rect 20947 41225 20959 41228
rect 20901 41219 20959 41225
rect 20640 41188 20668 41219
rect 21082 41216 21088 41228
rect 21140 41216 21146 41268
rect 21174 41216 21180 41268
rect 21232 41216 21238 41268
rect 21266 41216 21272 41268
rect 21324 41256 21330 41268
rect 21453 41259 21511 41265
rect 21453 41256 21465 41259
rect 21324 41228 21465 41256
rect 21324 41216 21330 41228
rect 21453 41225 21465 41228
rect 21499 41225 21511 41259
rect 21453 41219 21511 41225
rect 21726 41216 21732 41268
rect 21784 41256 21790 41268
rect 21784 41228 22048 41256
rect 21784 41216 21790 41228
rect 21192 41188 21220 41216
rect 20640 41160 21220 41188
rect 21284 41160 21956 41188
rect 19291 41092 19564 41120
rect 19291 41089 19303 41092
rect 19245 41083 19303 41089
rect 19702 41080 19708 41132
rect 19760 41080 19766 41132
rect 19886 41080 19892 41132
rect 19944 41120 19950 41132
rect 19981 41123 20039 41129
rect 19981 41120 19993 41123
rect 19944 41092 19993 41120
rect 19944 41080 19950 41092
rect 19981 41089 19993 41092
rect 20027 41089 20039 41123
rect 19981 41083 20039 41089
rect 20257 41123 20315 41129
rect 20257 41089 20269 41123
rect 20303 41089 20315 41123
rect 20257 41083 20315 41089
rect 16298 41012 16304 41064
rect 16356 41052 16362 41064
rect 20272 41052 20300 41083
rect 20530 41080 20536 41132
rect 20588 41080 20594 41132
rect 20809 41123 20867 41129
rect 20809 41089 20821 41123
rect 20855 41089 20867 41123
rect 20809 41083 20867 41089
rect 16356 41024 20300 41052
rect 16356 41012 16362 41024
rect 20438 41012 20444 41064
rect 20496 41052 20502 41064
rect 20824 41052 20852 41083
rect 21082 41080 21088 41132
rect 21140 41080 21146 41132
rect 21174 41080 21180 41132
rect 21232 41120 21238 41132
rect 21284 41120 21312 41160
rect 21928 41132 21956 41160
rect 21232 41092 21312 41120
rect 21232 41080 21238 41092
rect 21358 41080 21364 41132
rect 21416 41080 21422 41132
rect 21542 41080 21548 41132
rect 21600 41080 21606 41132
rect 21637 41123 21695 41129
rect 21637 41089 21649 41123
rect 21683 41089 21695 41123
rect 21637 41083 21695 41089
rect 21560 41052 21588 41080
rect 20496 41024 20852 41052
rect 20916 41024 21588 41052
rect 21652 41052 21680 41083
rect 21910 41080 21916 41132
rect 21968 41080 21974 41132
rect 22020 41129 22048 41228
rect 22278 41216 22284 41268
rect 22336 41256 22342 41268
rect 22373 41259 22431 41265
rect 22373 41256 22385 41259
rect 22336 41228 22385 41256
rect 22336 41216 22342 41228
rect 22373 41225 22385 41228
rect 22419 41225 22431 41259
rect 22373 41219 22431 41225
rect 23109 41259 23167 41265
rect 23109 41225 23121 41259
rect 23155 41256 23167 41259
rect 23382 41256 23388 41268
rect 23155 41228 23388 41256
rect 23155 41225 23167 41228
rect 23109 41219 23167 41225
rect 23382 41216 23388 41228
rect 23440 41216 23446 41268
rect 24213 41259 24271 41265
rect 24213 41225 24225 41259
rect 24259 41256 24271 41259
rect 25038 41256 25044 41268
rect 24259 41228 25044 41256
rect 24259 41225 24271 41228
rect 24213 41219 24271 41225
rect 25038 41216 25044 41228
rect 25096 41216 25102 41268
rect 22094 41148 22100 41200
rect 22152 41188 22158 41200
rect 22152 41160 22876 41188
rect 22152 41148 22158 41160
rect 22005 41123 22063 41129
rect 22005 41089 22017 41123
rect 22051 41089 22063 41123
rect 22005 41083 22063 41089
rect 22186 41080 22192 41132
rect 22244 41120 22250 41132
rect 22281 41123 22339 41129
rect 22281 41120 22293 41123
rect 22244 41092 22293 41120
rect 22244 41080 22250 41092
rect 22281 41089 22293 41092
rect 22327 41089 22339 41123
rect 22281 41083 22339 41089
rect 22554 41080 22560 41132
rect 22612 41080 22618 41132
rect 22848 41129 22876 41160
rect 22833 41123 22891 41129
rect 22833 41089 22845 41123
rect 22879 41089 22891 41123
rect 22833 41083 22891 41089
rect 23106 41080 23112 41132
rect 23164 41120 23170 41132
rect 23385 41123 23443 41129
rect 23385 41120 23397 41123
rect 23164 41092 23397 41120
rect 23164 41080 23170 41092
rect 23385 41089 23397 41092
rect 23431 41089 23443 41123
rect 23385 41083 23443 41089
rect 23937 41123 23995 41129
rect 23937 41089 23949 41123
rect 23983 41089 23995 41123
rect 23937 41083 23995 41089
rect 22738 41052 22744 41064
rect 21652 41024 22744 41052
rect 20496 41012 20502 41024
rect 19702 40984 19708 40996
rect 10704 40956 19708 40984
rect 8588 40888 9260 40916
rect 9582 40876 9588 40928
rect 9640 40876 9646 40928
rect 9674 40876 9680 40928
rect 9732 40916 9738 40928
rect 10704 40916 10732 40956
rect 19702 40944 19708 40956
rect 19760 40944 19766 40996
rect 19978 40944 19984 40996
rect 20036 40984 20042 40996
rect 20349 40987 20407 40993
rect 20349 40984 20361 40987
rect 20036 40956 20361 40984
rect 20036 40944 20042 40956
rect 20349 40953 20361 40956
rect 20395 40953 20407 40987
rect 20349 40947 20407 40953
rect 20806 40944 20812 40996
rect 20864 40984 20870 40996
rect 20916 40984 20944 41024
rect 22738 41012 22744 41024
rect 22796 41012 22802 41064
rect 23198 41012 23204 41064
rect 23256 41052 23262 41064
rect 23952 41052 23980 41083
rect 23256 41024 23980 41052
rect 23256 41012 23262 41024
rect 20864 40956 20944 40984
rect 21177 40987 21235 40993
rect 20864 40944 20870 40956
rect 21177 40953 21189 40987
rect 21223 40984 21235 40987
rect 22002 40984 22008 40996
rect 21223 40956 22008 40984
rect 21223 40953 21235 40956
rect 21177 40947 21235 40953
rect 22002 40944 22008 40956
rect 22060 40944 22066 40996
rect 22097 40987 22155 40993
rect 22097 40953 22109 40987
rect 22143 40984 22155 40987
rect 22646 40984 22652 40996
rect 22143 40956 22652 40984
rect 22143 40953 22155 40956
rect 22097 40947 22155 40953
rect 22646 40944 22652 40956
rect 22704 40944 22710 40996
rect 9732 40888 10732 40916
rect 9732 40876 9738 40888
rect 11054 40876 11060 40928
rect 11112 40876 11118 40928
rect 19058 40876 19064 40928
rect 19116 40876 19122 40928
rect 19797 40919 19855 40925
rect 19797 40885 19809 40919
rect 19843 40916 19855 40919
rect 20622 40916 20628 40928
rect 19843 40888 20628 40916
rect 19843 40885 19855 40888
rect 19797 40879 19855 40885
rect 20622 40876 20628 40888
rect 20680 40876 20686 40928
rect 20714 40876 20720 40928
rect 20772 40916 20778 40928
rect 21821 40919 21879 40925
rect 21821 40916 21833 40919
rect 20772 40888 21833 40916
rect 20772 40876 20778 40888
rect 21821 40885 21833 40888
rect 21867 40885 21879 40919
rect 21821 40879 21879 40885
rect 21910 40876 21916 40928
rect 21968 40916 21974 40928
rect 22278 40916 22284 40928
rect 21968 40888 22284 40916
rect 21968 40876 21974 40888
rect 22278 40876 22284 40888
rect 22336 40876 22342 40928
rect 23658 40876 23664 40928
rect 23716 40876 23722 40928
rect 1104 40826 24840 40848
rect 1104 40774 3917 40826
rect 3969 40774 3981 40826
rect 4033 40774 4045 40826
rect 4097 40774 4109 40826
rect 4161 40774 4173 40826
rect 4225 40774 9851 40826
rect 9903 40774 9915 40826
rect 9967 40774 9979 40826
rect 10031 40774 10043 40826
rect 10095 40774 10107 40826
rect 10159 40774 15785 40826
rect 15837 40774 15849 40826
rect 15901 40774 15913 40826
rect 15965 40774 15977 40826
rect 16029 40774 16041 40826
rect 16093 40774 21719 40826
rect 21771 40774 21783 40826
rect 21835 40774 21847 40826
rect 21899 40774 21911 40826
rect 21963 40774 21975 40826
rect 22027 40774 24840 40826
rect 1104 40752 24840 40774
rect 3050 40672 3056 40724
rect 3108 40712 3114 40724
rect 3421 40715 3479 40721
rect 3421 40712 3433 40715
rect 3108 40684 3433 40712
rect 3108 40672 3114 40684
rect 3421 40681 3433 40684
rect 3467 40681 3479 40715
rect 3421 40675 3479 40681
rect 3896 40684 4844 40712
rect 3142 40604 3148 40656
rect 3200 40644 3206 40656
rect 3896 40644 3924 40684
rect 3200 40616 3924 40644
rect 3200 40604 3206 40616
rect 3510 40536 3516 40588
rect 3568 40576 3574 40588
rect 3786 40576 3792 40588
rect 3568 40548 3792 40576
rect 3568 40536 3574 40548
rect 3786 40536 3792 40548
rect 3844 40536 3850 40588
rect 3326 40468 3332 40520
rect 3384 40508 3390 40520
rect 3605 40511 3663 40517
rect 3605 40508 3617 40511
rect 3384 40480 3617 40508
rect 3384 40468 3390 40480
rect 3605 40477 3617 40480
rect 3651 40477 3663 40511
rect 3605 40471 3663 40477
rect 3970 40468 3976 40520
rect 4028 40508 4034 40520
rect 4063 40511 4121 40517
rect 4063 40508 4075 40511
rect 4028 40480 4075 40508
rect 4028 40468 4034 40480
rect 4063 40477 4075 40480
rect 4109 40477 4121 40511
rect 4816 40508 4844 40684
rect 5258 40672 5264 40724
rect 5316 40712 5322 40724
rect 5316 40684 7604 40712
rect 5316 40672 5322 40684
rect 7576 40644 7604 40684
rect 7650 40672 7656 40724
rect 7708 40712 7714 40724
rect 9674 40712 9680 40724
rect 7708 40684 9680 40712
rect 7708 40672 7714 40684
rect 9674 40672 9680 40684
rect 9732 40672 9738 40724
rect 9766 40672 9772 40724
rect 9824 40712 9830 40724
rect 11790 40712 11796 40724
rect 9824 40684 11796 40712
rect 9824 40672 9830 40684
rect 11790 40672 11796 40684
rect 11848 40672 11854 40724
rect 16298 40712 16304 40724
rect 11900 40684 16304 40712
rect 10318 40644 10324 40656
rect 7576 40616 9674 40644
rect 4890 40536 4896 40588
rect 4948 40576 4954 40588
rect 4948 40548 5580 40576
rect 4948 40536 4954 40548
rect 5552 40517 5580 40548
rect 5537 40511 5595 40517
rect 4816 40480 5488 40508
rect 4063 40471 4121 40477
rect 1394 40400 1400 40452
rect 1452 40400 1458 40452
rect 2222 40400 2228 40452
rect 2280 40400 2286 40452
rect 2409 40443 2467 40449
rect 2409 40409 2421 40443
rect 2455 40440 2467 40443
rect 2774 40440 2780 40452
rect 2455 40412 2780 40440
rect 2455 40409 2467 40412
rect 2409 40403 2467 40409
rect 2774 40400 2780 40412
rect 2832 40400 2838 40452
rect 3237 40443 3295 40449
rect 3237 40409 3249 40443
rect 3283 40440 3295 40443
rect 3510 40440 3516 40452
rect 3283 40412 3516 40440
rect 3283 40409 3295 40412
rect 3237 40403 3295 40409
rect 3510 40400 3516 40412
rect 3568 40400 3574 40452
rect 3786 40332 3792 40384
rect 3844 40372 3850 40384
rect 4801 40375 4859 40381
rect 4801 40372 4813 40375
rect 3844 40344 4813 40372
rect 3844 40332 3850 40344
rect 4801 40341 4813 40344
rect 4847 40341 4859 40375
rect 5460 40372 5488 40480
rect 5537 40477 5549 40511
rect 5583 40477 5595 40511
rect 5810 40508 5816 40520
rect 5771 40480 5816 40508
rect 5537 40471 5595 40477
rect 5552 40440 5580 40471
rect 5810 40468 5816 40480
rect 5868 40468 5874 40520
rect 6822 40468 6828 40520
rect 6880 40508 6886 40520
rect 6917 40511 6975 40517
rect 6917 40508 6929 40511
rect 6880 40480 6929 40508
rect 6880 40468 6886 40480
rect 6917 40477 6929 40480
rect 6963 40477 6975 40511
rect 6917 40471 6975 40477
rect 7191 40511 7249 40517
rect 7191 40477 7203 40511
rect 7237 40508 7249 40511
rect 7576 40508 7604 40616
rect 9306 40576 9312 40588
rect 7668 40548 9312 40576
rect 7668 40520 7696 40548
rect 9306 40536 9312 40548
rect 9364 40536 9370 40588
rect 9646 40576 9674 40616
rect 9876 40616 10324 40644
rect 9876 40576 9904 40616
rect 10318 40604 10324 40616
rect 10376 40604 10382 40656
rect 10502 40604 10508 40656
rect 10560 40604 10566 40656
rect 11900 40644 11928 40684
rect 16298 40672 16304 40684
rect 16356 40672 16362 40724
rect 16390 40672 16396 40724
rect 16448 40672 16454 40724
rect 19794 40672 19800 40724
rect 19852 40712 19858 40724
rect 20533 40715 20591 40721
rect 20533 40712 20545 40715
rect 19852 40684 20545 40712
rect 19852 40672 19858 40684
rect 20533 40681 20545 40684
rect 20579 40681 20591 40715
rect 20533 40675 20591 40681
rect 20806 40672 20812 40724
rect 20864 40672 20870 40724
rect 20990 40672 20996 40724
rect 21048 40712 21054 40724
rect 21361 40715 21419 40721
rect 21361 40712 21373 40715
rect 21048 40684 21373 40712
rect 21048 40672 21054 40684
rect 21361 40681 21373 40684
rect 21407 40681 21419 40715
rect 21361 40675 21419 40681
rect 21637 40715 21695 40721
rect 21637 40681 21649 40715
rect 21683 40712 21695 40715
rect 22094 40712 22100 40724
rect 21683 40684 22100 40712
rect 21683 40681 21695 40684
rect 21637 40675 21695 40681
rect 22094 40672 22100 40684
rect 22152 40672 22158 40724
rect 22189 40715 22247 40721
rect 22189 40681 22201 40715
rect 22235 40712 22247 40715
rect 22554 40712 22560 40724
rect 22235 40684 22560 40712
rect 22235 40681 22247 40684
rect 22189 40675 22247 40681
rect 22554 40672 22560 40684
rect 22612 40672 22618 40724
rect 22738 40672 22744 40724
rect 22796 40672 22802 40724
rect 23014 40672 23020 40724
rect 23072 40672 23078 40724
rect 23477 40715 23535 40721
rect 23477 40681 23489 40715
rect 23523 40712 23535 40715
rect 24026 40712 24032 40724
rect 23523 40684 24032 40712
rect 23523 40681 23535 40684
rect 23477 40675 23535 40681
rect 24026 40672 24032 40684
rect 24084 40672 24090 40724
rect 11808 40616 11928 40644
rect 16408 40644 16436 40672
rect 19981 40647 20039 40653
rect 19981 40644 19993 40647
rect 16408 40616 19993 40644
rect 9646 40548 9904 40576
rect 10042 40536 10048 40588
rect 10100 40536 10106 40588
rect 10870 40576 10876 40588
rect 10928 40585 10934 40588
rect 10928 40579 10956 40585
rect 10152 40548 10876 40576
rect 7237 40480 7604 40508
rect 7237 40477 7249 40480
rect 7191 40471 7249 40477
rect 7650 40468 7656 40520
rect 7708 40468 7714 40520
rect 9766 40508 9772 40520
rect 9646 40480 9772 40508
rect 6086 40440 6092 40452
rect 5552 40412 6092 40440
rect 6086 40400 6092 40412
rect 6144 40440 6150 40452
rect 6362 40440 6368 40452
rect 6144 40412 6368 40440
rect 6144 40400 6150 40412
rect 6362 40400 6368 40412
rect 6420 40400 6426 40452
rect 9646 40440 9674 40480
rect 9766 40468 9772 40480
rect 9824 40468 9830 40520
rect 9861 40511 9919 40517
rect 9861 40477 9873 40511
rect 9907 40477 9919 40511
rect 9861 40471 9919 40477
rect 6472 40412 9674 40440
rect 6472 40372 6500 40412
rect 5460 40344 6500 40372
rect 6549 40375 6607 40381
rect 4801 40335 4859 40341
rect 6549 40341 6561 40375
rect 6595 40372 6607 40375
rect 6638 40372 6644 40384
rect 6595 40344 6644 40372
rect 6595 40341 6607 40344
rect 6549 40335 6607 40341
rect 6638 40332 6644 40344
rect 6696 40332 6702 40384
rect 7926 40332 7932 40384
rect 7984 40332 7990 40384
rect 9122 40332 9128 40384
rect 9180 40372 9186 40384
rect 9766 40372 9772 40384
rect 9180 40344 9772 40372
rect 9180 40332 9186 40344
rect 9766 40332 9772 40344
rect 9824 40332 9830 40384
rect 9876 40372 9904 40471
rect 9950 40468 9956 40520
rect 10008 40508 10014 40520
rect 10152 40508 10180 40548
rect 10870 40536 10876 40548
rect 10944 40545 10956 40579
rect 10928 40539 10956 40545
rect 10928 40536 10934 40539
rect 11054 40536 11060 40588
rect 11112 40536 11118 40588
rect 10008 40480 10180 40508
rect 10008 40468 10014 40480
rect 10778 40468 10784 40520
rect 10836 40468 10842 40520
rect 11698 40468 11704 40520
rect 11756 40508 11762 40520
rect 11808 40517 11836 40616
rect 19981 40613 19993 40616
rect 20027 40613 20039 40647
rect 19981 40607 20039 40613
rect 20254 40604 20260 40656
rect 20312 40604 20318 40656
rect 22465 40647 22523 40653
rect 22465 40644 22477 40647
rect 20548 40616 22477 40644
rect 19058 40536 19064 40588
rect 19116 40576 19122 40588
rect 19116 40548 19380 40576
rect 19116 40536 19122 40548
rect 11793 40511 11851 40517
rect 11793 40508 11805 40511
rect 11756 40480 11805 40508
rect 11756 40468 11762 40480
rect 11793 40477 11805 40480
rect 11839 40477 11851 40511
rect 11793 40471 11851 40477
rect 12051 40481 12109 40487
rect 12051 40447 12063 40481
rect 12097 40478 12109 40481
rect 12097 40447 12112 40478
rect 12526 40468 12532 40520
rect 12584 40468 12590 40520
rect 12710 40468 12716 40520
rect 12768 40508 12774 40520
rect 19352 40517 19380 40548
rect 13357 40511 13415 40517
rect 13357 40508 13369 40511
rect 12768 40480 13369 40508
rect 12768 40468 12774 40480
rect 13357 40477 13369 40480
rect 13403 40477 13415 40511
rect 13357 40471 13415 40477
rect 19337 40511 19395 40517
rect 19337 40477 19349 40511
rect 19383 40477 19395 40511
rect 19337 40471 19395 40477
rect 19518 40468 19524 40520
rect 19576 40508 19582 40520
rect 19797 40511 19855 40517
rect 19797 40508 19809 40511
rect 19576 40480 19809 40508
rect 19576 40468 19582 40480
rect 19797 40477 19809 40480
rect 19843 40477 19855 40511
rect 19797 40471 19855 40477
rect 20162 40468 20168 40520
rect 20220 40468 20226 40520
rect 20441 40511 20499 40517
rect 20441 40477 20453 40511
rect 20487 40508 20499 40511
rect 20548 40508 20576 40616
rect 22465 40613 22477 40616
rect 22511 40613 22523 40647
rect 25314 40644 25320 40656
rect 22465 40607 22523 40613
rect 22664 40616 25320 40644
rect 21174 40536 21180 40588
rect 21232 40536 21238 40588
rect 21358 40536 21364 40588
rect 21416 40536 21422 40588
rect 22664 40576 22692 40616
rect 25314 40604 25320 40616
rect 25372 40604 25378 40656
rect 21560 40548 22048 40576
rect 20487 40480 20576 40508
rect 20717 40511 20775 40517
rect 20487 40477 20499 40480
rect 20441 40471 20499 40477
rect 20717 40477 20729 40511
rect 20763 40477 20775 40511
rect 20717 40471 20775 40477
rect 12051 40441 12112 40447
rect 12084 40440 12112 40441
rect 12544 40440 12572 40468
rect 13538 40440 13544 40452
rect 12084 40412 13544 40440
rect 13538 40400 13544 40412
rect 13596 40400 13602 40452
rect 19150 40400 19156 40452
rect 19208 40440 19214 40452
rect 20732 40440 20760 40471
rect 20990 40468 20996 40520
rect 21048 40468 21054 40520
rect 21192 40440 21220 40536
rect 21266 40468 21272 40520
rect 21324 40468 21330 40520
rect 19208 40412 20760 40440
rect 20824 40412 21220 40440
rect 21376 40440 21404 40536
rect 21560 40517 21588 40548
rect 21545 40511 21603 40517
rect 21545 40477 21557 40511
rect 21591 40477 21603 40511
rect 21545 40471 21603 40477
rect 21821 40511 21879 40517
rect 21821 40477 21833 40511
rect 21867 40508 21879 40511
rect 21867 40480 21956 40508
rect 21867 40477 21879 40480
rect 21821 40471 21879 40477
rect 21726 40440 21732 40452
rect 21376 40412 21732 40440
rect 19208 40400 19214 40412
rect 11514 40372 11520 40384
rect 9876 40344 11520 40372
rect 11514 40332 11520 40344
rect 11572 40332 11578 40384
rect 11701 40375 11759 40381
rect 11701 40341 11713 40375
rect 11747 40372 11759 40375
rect 12342 40372 12348 40384
rect 11747 40344 12348 40372
rect 11747 40341 11759 40344
rect 11701 40335 11759 40341
rect 12342 40332 12348 40344
rect 12400 40332 12406 40384
rect 12526 40332 12532 40384
rect 12584 40372 12590 40384
rect 12805 40375 12863 40381
rect 12805 40372 12817 40375
rect 12584 40344 12817 40372
rect 12584 40332 12590 40344
rect 12805 40341 12817 40344
rect 12851 40341 12863 40375
rect 12805 40335 12863 40341
rect 19426 40332 19432 40384
rect 19484 40332 19490 40384
rect 19610 40332 19616 40384
rect 19668 40332 19674 40384
rect 19794 40332 19800 40384
rect 19852 40372 19858 40384
rect 20824 40372 20852 40412
rect 21726 40400 21732 40412
rect 21784 40400 21790 40452
rect 19852 40344 20852 40372
rect 21085 40375 21143 40381
rect 19852 40332 19858 40344
rect 21085 40341 21097 40375
rect 21131 40372 21143 40375
rect 21634 40372 21640 40384
rect 21131 40344 21640 40372
rect 21131 40341 21143 40344
rect 21085 40335 21143 40341
rect 21634 40332 21640 40344
rect 21692 40332 21698 40384
rect 21928 40381 21956 40480
rect 21913 40375 21971 40381
rect 21913 40341 21925 40375
rect 21959 40341 21971 40375
rect 22020 40372 22048 40548
rect 22112 40548 22692 40576
rect 22112 40517 22140 40548
rect 22738 40536 22744 40588
rect 22796 40576 22802 40588
rect 22796 40548 23244 40576
rect 22796 40536 22802 40548
rect 22097 40511 22155 40517
rect 22097 40477 22109 40511
rect 22143 40477 22155 40511
rect 22097 40471 22155 40477
rect 22370 40468 22376 40520
rect 22428 40468 22434 40520
rect 22646 40468 22652 40520
rect 22704 40468 22710 40520
rect 22922 40468 22928 40520
rect 22980 40468 22986 40520
rect 23216 40517 23244 40548
rect 23201 40511 23259 40517
rect 23201 40477 23213 40511
rect 23247 40477 23259 40511
rect 23201 40471 23259 40477
rect 23658 40468 23664 40520
rect 23716 40468 23722 40520
rect 22278 40400 22284 40452
rect 22336 40440 22342 40452
rect 23845 40443 23903 40449
rect 23845 40440 23857 40443
rect 22336 40412 23857 40440
rect 22336 40400 22342 40412
rect 23845 40409 23857 40412
rect 23891 40409 23903 40443
rect 23845 40403 23903 40409
rect 24213 40443 24271 40449
rect 24213 40409 24225 40443
rect 24259 40440 24271 40443
rect 25130 40440 25136 40452
rect 24259 40412 25136 40440
rect 24259 40409 24271 40412
rect 24213 40403 24271 40409
rect 25130 40400 25136 40412
rect 25188 40400 25194 40452
rect 22922 40372 22928 40384
rect 22020 40344 22928 40372
rect 21913 40335 21971 40341
rect 22922 40332 22928 40344
rect 22980 40332 22986 40384
rect 1104 40282 25000 40304
rect 1104 40230 6884 40282
rect 6936 40230 6948 40282
rect 7000 40230 7012 40282
rect 7064 40230 7076 40282
rect 7128 40230 7140 40282
rect 7192 40230 12818 40282
rect 12870 40230 12882 40282
rect 12934 40230 12946 40282
rect 12998 40230 13010 40282
rect 13062 40230 13074 40282
rect 13126 40230 18752 40282
rect 18804 40230 18816 40282
rect 18868 40230 18880 40282
rect 18932 40230 18944 40282
rect 18996 40230 19008 40282
rect 19060 40230 24686 40282
rect 24738 40230 24750 40282
rect 24802 40230 24814 40282
rect 24866 40230 24878 40282
rect 24930 40230 24942 40282
rect 24994 40230 25000 40282
rect 1104 40208 25000 40230
rect 3142 40168 3148 40180
rect 1688 40140 3148 40168
rect 1688 40109 1716 40140
rect 3142 40128 3148 40140
rect 3200 40128 3206 40180
rect 3510 40128 3516 40180
rect 3568 40168 3574 40180
rect 3568 40140 7420 40168
rect 3568 40128 3574 40140
rect 1673 40103 1731 40109
rect 1673 40069 1685 40103
rect 1719 40069 1731 40103
rect 7392 40100 7420 40140
rect 7466 40128 7472 40180
rect 7524 40128 7530 40180
rect 8018 40128 8024 40180
rect 8076 40168 8082 40180
rect 8076 40140 9260 40168
rect 8076 40128 8082 40140
rect 9232 40112 9260 40140
rect 9306 40128 9312 40180
rect 9364 40168 9370 40180
rect 9364 40140 19196 40168
rect 9364 40128 9370 40140
rect 7558 40100 7564 40112
rect 1673 40063 1731 40069
rect 2746 40072 3464 40100
rect 2223 40045 2281 40051
rect 1397 40035 1455 40041
rect 1397 40001 1409 40035
rect 1443 40032 1455 40035
rect 1578 40032 1584 40044
rect 1443 40004 1584 40032
rect 1443 40001 1455 40004
rect 1397 39995 1455 40001
rect 1578 39992 1584 40004
rect 1636 39992 1642 40044
rect 2223 40011 2235 40045
rect 2269 40032 2281 40045
rect 2746 40032 2774 40072
rect 3436 40044 3464 40072
rect 3988 40072 4844 40100
rect 2269 40011 2774 40032
rect 2223 40005 2774 40011
rect 2240 40004 2774 40005
rect 3142 39992 3148 40044
rect 3200 40032 3206 40044
rect 3329 40035 3387 40041
rect 3329 40032 3341 40035
rect 3200 40004 3341 40032
rect 3200 39992 3206 40004
rect 3329 40001 3341 40004
rect 3375 40001 3387 40035
rect 3329 39995 3387 40001
rect 3418 39992 3424 40044
rect 3476 39992 3482 40044
rect 1854 39924 1860 39976
rect 1912 39964 1918 39976
rect 1949 39967 2007 39973
rect 1949 39964 1961 39967
rect 1912 39936 1961 39964
rect 1912 39924 1918 39936
rect 1949 39933 1961 39936
rect 1995 39933 2007 39967
rect 1949 39927 2007 39933
rect 3050 39924 3056 39976
rect 3108 39964 3114 39976
rect 3513 39967 3571 39973
rect 3513 39964 3525 39967
rect 3108 39936 3525 39964
rect 3108 39924 3114 39936
rect 3513 39933 3525 39936
rect 3559 39933 3571 39967
rect 3513 39927 3571 39933
rect 3988 39908 4016 40072
rect 4816 40042 4844 40072
rect 5644 40072 7328 40100
rect 7392 40072 7564 40100
rect 4816 40032 5028 40042
rect 5135 40035 5193 40041
rect 5135 40032 5147 40035
rect 4816 40014 5147 40032
rect 5000 40004 5147 40014
rect 5135 40001 5147 40004
rect 5181 40032 5193 40035
rect 5644 40032 5672 40072
rect 5181 40004 5672 40032
rect 7300 40032 7328 40072
rect 7558 40060 7564 40072
rect 7616 40060 7622 40112
rect 7837 40103 7895 40109
rect 7837 40069 7849 40103
rect 7883 40100 7895 40103
rect 8386 40100 8392 40112
rect 7883 40072 8392 40100
rect 7883 40069 7895 40072
rect 7837 40063 7895 40069
rect 8386 40060 8392 40072
rect 8444 40060 8450 40112
rect 8573 40103 8631 40109
rect 8573 40069 8585 40103
rect 8619 40100 8631 40103
rect 8619 40072 9076 40100
rect 8619 40069 8631 40072
rect 8573 40063 8631 40069
rect 7650 40032 7656 40044
rect 7300 40004 7656 40032
rect 5181 40001 5193 40004
rect 5135 39995 5193 40001
rect 7650 39992 7656 40004
rect 7708 39992 7714 40044
rect 7745 40035 7803 40041
rect 7745 40001 7757 40035
rect 7791 40032 7803 40035
rect 8018 40032 8024 40044
rect 7791 40004 8024 40032
rect 7791 40001 7803 40004
rect 7745 39995 7803 40001
rect 8018 39992 8024 40004
rect 8076 39992 8082 40044
rect 8110 39992 8116 40044
rect 8168 40032 8174 40044
rect 8205 40035 8263 40041
rect 8205 40032 8217 40035
rect 8168 40004 8217 40032
rect 8168 39992 8174 40004
rect 8205 40001 8217 40004
rect 8251 40001 8263 40035
rect 9048 40032 9076 40072
rect 9122 40060 9128 40112
rect 9180 40060 9186 40112
rect 9214 40060 9220 40112
rect 9272 40100 9278 40112
rect 9401 40103 9459 40109
rect 9401 40100 9413 40103
rect 9272 40072 9413 40100
rect 9272 40060 9278 40072
rect 9401 40069 9413 40072
rect 9447 40069 9459 40103
rect 9401 40063 9459 40069
rect 9490 40060 9496 40112
rect 9548 40060 9554 40112
rect 9766 40100 9772 40112
rect 9600 40072 9772 40100
rect 9600 40032 9628 40072
rect 9766 40060 9772 40072
rect 9824 40100 9830 40112
rect 10042 40100 10048 40112
rect 9824 40072 10048 40100
rect 9824 40060 9830 40072
rect 10042 40060 10048 40072
rect 10100 40100 10106 40112
rect 10229 40103 10287 40109
rect 10229 40100 10241 40103
rect 10100 40072 10241 40100
rect 10100 40060 10106 40072
rect 10229 40069 10241 40072
rect 10275 40069 10287 40103
rect 10229 40063 10287 40069
rect 10318 40060 10324 40112
rect 10376 40100 10382 40112
rect 10686 40100 10692 40112
rect 10376 40072 10692 40100
rect 10376 40060 10382 40072
rect 10686 40060 10692 40072
rect 10744 40060 10750 40112
rect 10778 40060 10784 40112
rect 10836 40100 10842 40112
rect 10836 40072 11100 40100
rect 10836 40060 10842 40072
rect 9048 40004 9628 40032
rect 8205 39995 8263 40001
rect 9674 39992 9680 40044
rect 9732 40032 9738 40044
rect 11072 40041 11100 40072
rect 9861 40035 9919 40041
rect 9861 40032 9873 40035
rect 9732 40004 9873 40032
rect 9732 39992 9738 40004
rect 9861 40001 9873 40004
rect 9907 40001 9919 40035
rect 9861 39995 9919 40001
rect 11057 40035 11115 40041
rect 11057 40001 11069 40035
rect 11103 40001 11115 40035
rect 11057 39995 11115 40001
rect 12710 39992 12716 40044
rect 12768 39992 12774 40044
rect 19168 40032 19196 40140
rect 19610 40128 19616 40180
rect 19668 40128 19674 40180
rect 19794 40128 19800 40180
rect 19852 40128 19858 40180
rect 20070 40128 20076 40180
rect 20128 40128 20134 40180
rect 20901 40171 20959 40177
rect 20901 40168 20913 40171
rect 20272 40140 20913 40168
rect 19245 40103 19303 40109
rect 19245 40069 19257 40103
rect 19291 40100 19303 40103
rect 19628 40100 19656 40128
rect 19291 40072 19656 40100
rect 19291 40069 19303 40072
rect 19245 40063 19303 40069
rect 19168 40004 19334 40032
rect 4338 39924 4344 39976
rect 4396 39964 4402 39976
rect 4433 39967 4491 39973
rect 4433 39964 4445 39967
rect 4396 39936 4445 39964
rect 4396 39924 4402 39936
rect 4433 39933 4445 39936
rect 4479 39964 4491 39967
rect 4798 39964 4804 39976
rect 4479 39936 4804 39964
rect 4479 39933 4491 39936
rect 4433 39927 4491 39933
rect 4798 39924 4804 39936
rect 4856 39924 4862 39976
rect 4890 39924 4896 39976
rect 4948 39924 4954 39976
rect 7926 39924 7932 39976
rect 7984 39924 7990 39976
rect 9582 39924 9588 39976
rect 9640 39924 9646 39976
rect 11422 39924 11428 39976
rect 11480 39964 11486 39976
rect 11793 39967 11851 39973
rect 11793 39964 11805 39967
rect 11480 39936 11805 39964
rect 11480 39924 11486 39936
rect 11793 39933 11805 39936
rect 11839 39933 11851 39967
rect 11793 39927 11851 39933
rect 11882 39924 11888 39976
rect 11940 39964 11946 39976
rect 11977 39967 12035 39973
rect 11977 39964 11989 39967
rect 11940 39936 11989 39964
rect 11940 39924 11946 39936
rect 11977 39933 11989 39936
rect 12023 39933 12035 39967
rect 11977 39927 12035 39933
rect 12342 39924 12348 39976
rect 12400 39964 12406 39976
rect 12830 39967 12888 39973
rect 12830 39964 12842 39967
rect 12400 39936 12842 39964
rect 12400 39924 12406 39936
rect 12830 39933 12842 39936
rect 12876 39933 12888 39967
rect 12830 39927 12888 39933
rect 12989 39967 13047 39973
rect 12989 39933 13001 39967
rect 13035 39964 13047 39967
rect 13354 39964 13360 39976
rect 13035 39936 13360 39964
rect 13035 39933 13047 39936
rect 12989 39927 13047 39933
rect 13354 39924 13360 39936
rect 13412 39924 13418 39976
rect 19306 39964 19334 40004
rect 19978 39992 19984 40044
rect 20036 39992 20042 40044
rect 20272 40041 20300 40140
rect 20901 40137 20913 40140
rect 20947 40137 20959 40171
rect 20901 40131 20959 40137
rect 21177 40171 21235 40177
rect 21177 40137 21189 40171
rect 21223 40168 21235 40171
rect 21223 40140 23428 40168
rect 21223 40137 21235 40140
rect 21177 40131 21235 40137
rect 20714 40100 20720 40112
rect 20456 40072 20720 40100
rect 20257 40035 20315 40041
rect 20257 40001 20269 40035
rect 20303 40001 20315 40035
rect 20456 40032 20484 40072
rect 20714 40060 20720 40072
rect 20772 40060 20778 40112
rect 21542 40060 21548 40112
rect 21600 40100 21606 40112
rect 21600 40072 22048 40100
rect 21600 40060 21606 40072
rect 20525 40035 20583 40041
rect 20525 40032 20537 40035
rect 20456 40004 20537 40032
rect 20257 39995 20315 40001
rect 20525 40001 20537 40004
rect 20571 40001 20583 40035
rect 20525 39995 20583 40001
rect 20806 39992 20812 40044
rect 20864 39992 20870 40044
rect 21082 39992 21088 40044
rect 21140 39992 21146 40044
rect 21358 39992 21364 40044
rect 21416 39992 21422 40044
rect 21637 40035 21695 40041
rect 21637 40001 21649 40035
rect 21683 40001 21695 40035
rect 21637 39995 21695 40001
rect 21652 39964 21680 39995
rect 21726 39992 21732 40044
rect 21784 39992 21790 40044
rect 22020 40041 22048 40072
rect 22112 40072 22692 40100
rect 22005 40035 22063 40041
rect 22005 40001 22017 40035
rect 22051 40001 22063 40035
rect 22005 39995 22063 40001
rect 19306 39936 21680 39964
rect 21744 39964 21772 39992
rect 22112 39964 22140 40072
rect 22281 40035 22339 40041
rect 22281 40001 22293 40035
rect 22327 40032 22339 40035
rect 22462 40032 22468 40044
rect 22327 40004 22468 40032
rect 22327 40001 22339 40004
rect 22281 39995 22339 40001
rect 22462 39992 22468 40004
rect 22520 39992 22526 40044
rect 22557 40035 22615 40041
rect 22557 40001 22569 40035
rect 22603 40001 22615 40035
rect 22557 39995 22615 40001
rect 21744 39936 22140 39964
rect 2866 39856 2872 39908
rect 2924 39896 2930 39908
rect 3970 39896 3976 39908
rect 2924 39868 3976 39896
rect 2924 39856 2930 39868
rect 3970 39856 3976 39868
rect 4028 39856 4034 39908
rect 12437 39899 12495 39905
rect 12437 39865 12449 39899
rect 12483 39896 12495 39899
rect 12526 39896 12532 39908
rect 12483 39868 12532 39896
rect 12483 39865 12495 39868
rect 12437 39859 12495 39865
rect 12526 39856 12532 39868
rect 12584 39856 12590 39908
rect 19426 39856 19432 39908
rect 19484 39856 19490 39908
rect 20625 39899 20683 39905
rect 20625 39865 20637 39899
rect 20671 39896 20683 39899
rect 20806 39896 20812 39908
rect 20671 39868 20812 39896
rect 20671 39865 20683 39868
rect 20625 39859 20683 39865
rect 20806 39856 20812 39868
rect 20864 39856 20870 39908
rect 22572 39896 22600 39995
rect 22664 39905 22692 40072
rect 22833 40035 22891 40041
rect 22833 40001 22845 40035
rect 22879 40032 22891 40035
rect 23014 40032 23020 40044
rect 22879 40004 23020 40032
rect 22879 40001 22891 40004
rect 22833 39995 22891 40001
rect 23014 39992 23020 40004
rect 23072 39992 23078 40044
rect 23400 40041 23428 40140
rect 23842 40128 23848 40180
rect 23900 40128 23906 40180
rect 23860 40100 23888 40128
rect 23492 40072 23888 40100
rect 23109 40035 23167 40041
rect 23109 40001 23121 40035
rect 23155 40001 23167 40035
rect 23109 39995 23167 40001
rect 23385 40035 23443 40041
rect 23385 40001 23397 40035
rect 23431 40001 23443 40035
rect 23385 39995 23443 40001
rect 23124 39964 23152 39995
rect 23032 39936 23152 39964
rect 23032 39908 23060 39936
rect 21008 39868 22600 39896
rect 22649 39899 22707 39905
rect 2314 39788 2320 39840
rect 2372 39828 2378 39840
rect 2961 39831 3019 39837
rect 2961 39828 2973 39831
rect 2372 39800 2973 39828
rect 2372 39788 2378 39800
rect 2961 39797 2973 39800
rect 3007 39797 3019 39831
rect 2961 39791 3019 39797
rect 3418 39788 3424 39840
rect 3476 39828 3482 39840
rect 4065 39831 4123 39837
rect 4065 39828 4077 39831
rect 3476 39800 4077 39828
rect 3476 39788 3482 39800
rect 4065 39797 4077 39800
rect 4111 39797 4123 39831
rect 4065 39791 4123 39797
rect 4246 39788 4252 39840
rect 4304 39828 4310 39840
rect 5350 39828 5356 39840
rect 4304 39800 5356 39828
rect 4304 39788 4310 39800
rect 5350 39788 5356 39800
rect 5408 39788 5414 39840
rect 5902 39788 5908 39840
rect 5960 39788 5966 39840
rect 8662 39788 8668 39840
rect 8720 39828 8726 39840
rect 8757 39831 8815 39837
rect 8757 39828 8769 39831
rect 8720 39800 8769 39828
rect 8720 39788 8726 39800
rect 8757 39797 8769 39800
rect 8803 39797 8815 39831
rect 8757 39791 8815 39797
rect 10318 39788 10324 39840
rect 10376 39828 10382 39840
rect 10413 39831 10471 39837
rect 10413 39828 10425 39831
rect 10376 39800 10425 39828
rect 10376 39788 10382 39800
rect 10413 39797 10425 39800
rect 10459 39797 10471 39831
rect 10413 39791 10471 39797
rect 13630 39788 13636 39840
rect 13688 39788 13694 39840
rect 20349 39831 20407 39837
rect 20349 39797 20361 39831
rect 20395 39828 20407 39831
rect 21008 39828 21036 39868
rect 22649 39865 22661 39899
rect 22695 39865 22707 39899
rect 22649 39859 22707 39865
rect 22830 39856 22836 39908
rect 22888 39856 22894 39908
rect 23014 39856 23020 39908
rect 23072 39856 23078 39908
rect 23201 39899 23259 39905
rect 23201 39865 23213 39899
rect 23247 39896 23259 39899
rect 23492 39896 23520 40072
rect 23750 39992 23756 40044
rect 23808 40032 23814 40044
rect 23845 40035 23903 40041
rect 23845 40032 23857 40035
rect 23808 40004 23857 40032
rect 23808 39992 23814 40004
rect 23845 40001 23857 40004
rect 23891 40001 23903 40035
rect 23845 39995 23903 40001
rect 24026 39992 24032 40044
rect 24084 40032 24090 40044
rect 24121 40035 24179 40041
rect 24121 40032 24133 40035
rect 24084 40004 24133 40032
rect 24084 39992 24090 40004
rect 24121 40001 24133 40004
rect 24167 40001 24179 40035
rect 24121 39995 24179 40001
rect 23247 39868 23520 39896
rect 23247 39865 23259 39868
rect 23201 39859 23259 39865
rect 20395 39800 21036 39828
rect 20395 39797 20407 39800
rect 20349 39791 20407 39797
rect 21082 39788 21088 39840
rect 21140 39828 21146 39840
rect 21453 39831 21511 39837
rect 21453 39828 21465 39831
rect 21140 39800 21465 39828
rect 21140 39788 21146 39800
rect 21453 39797 21465 39800
rect 21499 39797 21511 39831
rect 21453 39791 21511 39797
rect 21634 39788 21640 39840
rect 21692 39828 21698 39840
rect 21821 39831 21879 39837
rect 21821 39828 21833 39831
rect 21692 39800 21833 39828
rect 21692 39788 21698 39800
rect 21821 39797 21833 39800
rect 21867 39797 21879 39831
rect 21821 39791 21879 39797
rect 22097 39831 22155 39837
rect 22097 39797 22109 39831
rect 22143 39828 22155 39831
rect 22278 39828 22284 39840
rect 22143 39800 22284 39828
rect 22143 39797 22155 39800
rect 22097 39791 22155 39797
rect 22278 39788 22284 39800
rect 22336 39788 22342 39840
rect 22373 39831 22431 39837
rect 22373 39797 22385 39831
rect 22419 39828 22431 39831
rect 22848 39828 22876 39856
rect 22419 39800 22876 39828
rect 22419 39797 22431 39800
rect 22373 39791 22431 39797
rect 22922 39788 22928 39840
rect 22980 39788 22986 39840
rect 23661 39831 23719 39837
rect 23661 39797 23673 39831
rect 23707 39828 23719 39831
rect 23934 39828 23940 39840
rect 23707 39800 23940 39828
rect 23707 39797 23719 39800
rect 23661 39791 23719 39797
rect 23934 39788 23940 39800
rect 23992 39788 23998 39840
rect 24394 39788 24400 39840
rect 24452 39788 24458 39840
rect 1104 39738 24840 39760
rect 1104 39686 3917 39738
rect 3969 39686 3981 39738
rect 4033 39686 4045 39738
rect 4097 39686 4109 39738
rect 4161 39686 4173 39738
rect 4225 39686 9851 39738
rect 9903 39686 9915 39738
rect 9967 39686 9979 39738
rect 10031 39686 10043 39738
rect 10095 39686 10107 39738
rect 10159 39686 15785 39738
rect 15837 39686 15849 39738
rect 15901 39686 15913 39738
rect 15965 39686 15977 39738
rect 16029 39686 16041 39738
rect 16093 39686 21719 39738
rect 21771 39686 21783 39738
rect 21835 39686 21847 39738
rect 21899 39686 21911 39738
rect 21963 39686 21975 39738
rect 22027 39686 24840 39738
rect 1104 39664 24840 39686
rect 3418 39584 3424 39636
rect 3476 39584 3482 39636
rect 5902 39584 5908 39636
rect 5960 39624 5966 39636
rect 6730 39624 6736 39636
rect 5960 39596 6132 39624
rect 5960 39584 5966 39596
rect 3234 39516 3240 39568
rect 3292 39516 3298 39568
rect 2682 39448 2688 39500
rect 2740 39448 2746 39500
rect 2225 39423 2283 39429
rect 2225 39389 2237 39423
rect 2271 39420 2283 39423
rect 3436 39420 3464 39584
rect 6104 39565 6132 39596
rect 6196 39596 6736 39624
rect 5261 39559 5319 39565
rect 5261 39556 5273 39559
rect 5092 39528 5273 39556
rect 3792 39500 3844 39506
rect 5092 39500 5120 39528
rect 5261 39525 5273 39528
rect 5307 39525 5319 39559
rect 5261 39519 5319 39525
rect 6089 39559 6147 39565
rect 6089 39525 6101 39559
rect 6135 39525 6147 39559
rect 6089 39519 6147 39525
rect 5074 39448 5080 39500
rect 5132 39448 5138 39500
rect 5442 39448 5448 39500
rect 5500 39448 5506 39500
rect 6196 39488 6224 39596
rect 6730 39584 6736 39596
rect 6788 39624 6794 39636
rect 6788 39596 8340 39624
rect 6788 39584 6794 39596
rect 8312 39556 8340 39596
rect 8386 39584 8392 39636
rect 8444 39584 8450 39636
rect 9490 39584 9496 39636
rect 9548 39624 9554 39636
rect 10505 39627 10563 39633
rect 10505 39624 10517 39627
rect 9548 39596 10517 39624
rect 9548 39584 9554 39596
rect 10505 39593 10517 39596
rect 10551 39593 10563 39627
rect 10505 39587 10563 39593
rect 13354 39584 13360 39636
rect 13412 39584 13418 39636
rect 13630 39584 13636 39636
rect 13688 39584 13694 39636
rect 20717 39627 20775 39633
rect 20717 39593 20729 39627
rect 20763 39624 20775 39627
rect 20898 39624 20904 39636
rect 20763 39596 20904 39624
rect 20763 39593 20775 39596
rect 20717 39587 20775 39593
rect 20898 39584 20904 39596
rect 20956 39584 20962 39636
rect 20990 39584 20996 39636
rect 21048 39624 21054 39636
rect 21545 39627 21603 39633
rect 21545 39624 21557 39627
rect 21048 39596 21557 39624
rect 21048 39584 21054 39596
rect 21545 39593 21557 39596
rect 21591 39593 21603 39627
rect 21545 39587 21603 39593
rect 21821 39627 21879 39633
rect 21821 39593 21833 39627
rect 21867 39624 21879 39627
rect 22186 39624 22192 39636
rect 21867 39596 22192 39624
rect 21867 39593 21879 39596
rect 21821 39587 21879 39593
rect 22186 39584 22192 39596
rect 22244 39584 22250 39636
rect 22370 39584 22376 39636
rect 22428 39584 22434 39636
rect 22830 39584 22836 39636
rect 22888 39584 22894 39636
rect 8662 39556 8668 39568
rect 8312 39528 8668 39556
rect 8662 39516 8668 39528
rect 8720 39516 8726 39568
rect 13648 39556 13676 39584
rect 21174 39556 21180 39568
rect 13648 39528 21180 39556
rect 21174 39516 21180 39528
rect 21232 39516 21238 39568
rect 21358 39516 21364 39568
rect 21416 39556 21422 39568
rect 23201 39559 23259 39565
rect 23201 39556 23213 39559
rect 21416 39528 23213 39556
rect 21416 39516 21422 39528
rect 23201 39525 23213 39528
rect 23247 39525 23259 39559
rect 23201 39519 23259 39525
rect 6482 39491 6540 39497
rect 6482 39488 6494 39491
rect 6196 39460 6494 39488
rect 6482 39457 6494 39460
rect 6528 39457 6540 39491
rect 6482 39451 6540 39457
rect 6638 39448 6644 39500
rect 6696 39448 6702 39500
rect 6822 39448 6828 39500
rect 6880 39488 6886 39500
rect 7374 39488 7380 39500
rect 6880 39460 7380 39488
rect 6880 39448 6886 39460
rect 7374 39448 7380 39460
rect 7432 39448 7438 39500
rect 11698 39448 11704 39500
rect 11756 39488 11762 39500
rect 12345 39491 12403 39497
rect 12345 39488 12357 39491
rect 11756 39460 12357 39488
rect 11756 39448 11762 39460
rect 12345 39457 12357 39460
rect 12391 39457 12403 39491
rect 12345 39451 12403 39457
rect 20438 39448 20444 39500
rect 20496 39488 20502 39500
rect 20714 39488 20720 39500
rect 20496 39460 20720 39488
rect 20496 39448 20502 39460
rect 20714 39448 20720 39460
rect 20772 39448 20778 39500
rect 20824 39460 23428 39488
rect 3792 39442 3844 39448
rect 2271 39392 3464 39420
rect 4341 39423 4399 39429
rect 2271 39389 2283 39392
rect 2225 39383 2283 39389
rect 4341 39389 4353 39423
rect 4387 39420 4399 39423
rect 4522 39420 4528 39432
rect 4387 39392 4528 39420
rect 4387 39389 4399 39392
rect 4341 39383 4399 39389
rect 4522 39380 4528 39392
rect 4580 39380 4586 39432
rect 5460 39420 5488 39448
rect 4632 39392 5488 39420
rect 5629 39423 5687 39429
rect 1486 39312 1492 39364
rect 1544 39312 1550 39364
rect 1670 39312 1676 39364
rect 1728 39312 1734 39364
rect 2314 39312 2320 39364
rect 2372 39312 2378 39364
rect 2590 39312 2596 39364
rect 2648 39352 2654 39364
rect 2685 39355 2743 39361
rect 2685 39352 2697 39355
rect 2648 39324 2697 39352
rect 2648 39312 2654 39324
rect 2685 39321 2697 39324
rect 2731 39321 2743 39355
rect 2685 39315 2743 39321
rect 3053 39355 3111 39361
rect 3053 39321 3065 39355
rect 3099 39352 3111 39355
rect 3099 39324 4200 39352
rect 3099 39321 3111 39324
rect 3053 39315 3111 39321
rect 4172 39296 4200 39324
rect 4246 39312 4252 39364
rect 4304 39352 4310 39364
rect 4632 39352 4660 39392
rect 5629 39389 5641 39423
rect 5675 39389 5687 39423
rect 5629 39383 5687 39389
rect 4304 39324 4660 39352
rect 4709 39355 4767 39361
rect 4304 39312 4310 39324
rect 4709 39321 4721 39355
rect 4755 39352 4767 39355
rect 5644 39352 5672 39383
rect 6362 39380 6368 39432
rect 6420 39380 6426 39432
rect 7558 39380 7564 39432
rect 7616 39420 7622 39432
rect 7651 39423 7709 39429
rect 7651 39420 7663 39423
rect 7616 39392 7663 39420
rect 7616 39380 7622 39392
rect 7651 39389 7663 39392
rect 7697 39389 7709 39423
rect 7651 39383 7709 39389
rect 8570 39380 8576 39432
rect 8628 39420 8634 39432
rect 9493 39423 9551 39429
rect 9493 39420 9505 39423
rect 8628 39392 9505 39420
rect 8628 39380 8634 39392
rect 9493 39389 9505 39392
rect 9539 39389 9551 39423
rect 9493 39383 9551 39389
rect 9767 39423 9825 39429
rect 9767 39389 9779 39423
rect 9813 39420 9825 39423
rect 10226 39420 10232 39432
rect 9813 39392 10232 39420
rect 9813 39389 9825 39392
rect 9767 39383 9825 39389
rect 10226 39380 10232 39392
rect 10284 39420 10290 39432
rect 12587 39423 12645 39429
rect 12587 39420 12599 39423
rect 10284 39392 12599 39420
rect 10284 39380 10290 39392
rect 12587 39389 12599 39392
rect 12633 39389 12645 39423
rect 12587 39383 12645 39389
rect 16482 39380 16488 39432
rect 16540 39420 16546 39432
rect 20824 39420 20852 39460
rect 16540 39392 20852 39420
rect 16540 39380 16546 39392
rect 20898 39380 20904 39432
rect 20956 39380 20962 39432
rect 21269 39423 21327 39429
rect 21269 39420 21281 39423
rect 21008 39392 21281 39420
rect 4755 39324 5672 39352
rect 4755 39321 4767 39324
rect 4709 39315 4767 39321
rect 1949 39287 2007 39293
rect 1949 39253 1961 39287
rect 1995 39284 2007 39287
rect 3602 39284 3608 39296
rect 1995 39256 3608 39284
rect 1995 39253 2007 39256
rect 1949 39247 2007 39253
rect 3602 39244 3608 39256
rect 3660 39284 3666 39296
rect 3973 39287 4031 39293
rect 3973 39284 3985 39287
rect 3660 39256 3985 39284
rect 3660 39244 3666 39256
rect 3973 39253 3985 39256
rect 4019 39284 4031 39287
rect 4062 39284 4068 39296
rect 4019 39256 4068 39284
rect 4019 39253 4031 39256
rect 3973 39247 4031 39253
rect 4062 39244 4068 39256
rect 4120 39244 4126 39296
rect 4154 39244 4160 39296
rect 4212 39244 4218 39296
rect 4522 39244 4528 39296
rect 4580 39284 4586 39296
rect 4724 39284 4752 39315
rect 8018 39312 8024 39364
rect 8076 39352 8082 39364
rect 10318 39352 10324 39364
rect 8076 39324 10324 39352
rect 8076 39312 8082 39324
rect 10318 39312 10324 39324
rect 10376 39352 10382 39364
rect 11974 39352 11980 39364
rect 10376 39324 11980 39352
rect 10376 39312 10382 39324
rect 11974 39312 11980 39324
rect 12032 39312 12038 39364
rect 20070 39312 20076 39364
rect 20128 39352 20134 39364
rect 20806 39352 20812 39364
rect 20128 39324 20812 39352
rect 20128 39312 20134 39324
rect 20806 39312 20812 39324
rect 20864 39312 20870 39364
rect 4580 39256 4752 39284
rect 4580 39244 4586 39256
rect 4890 39244 4896 39296
rect 4948 39284 4954 39296
rect 5077 39287 5135 39293
rect 5077 39284 5089 39287
rect 4948 39256 5089 39284
rect 4948 39244 4954 39256
rect 5077 39253 5089 39256
rect 5123 39253 5135 39287
rect 5077 39247 5135 39253
rect 5350 39244 5356 39296
rect 5408 39284 5414 39296
rect 7285 39287 7343 39293
rect 7285 39284 7297 39287
rect 5408 39256 7297 39284
rect 5408 39244 5414 39256
rect 7285 39253 7297 39256
rect 7331 39253 7343 39287
rect 7285 39247 7343 39253
rect 20438 39244 20444 39296
rect 20496 39284 20502 39296
rect 21008 39284 21036 39392
rect 21269 39389 21281 39392
rect 21315 39389 21327 39423
rect 21269 39383 21327 39389
rect 21450 39380 21456 39432
rect 21508 39420 21514 39432
rect 21729 39423 21787 39429
rect 21729 39420 21741 39423
rect 21508 39392 21741 39420
rect 21508 39380 21514 39392
rect 21729 39389 21741 39392
rect 21775 39389 21787 39423
rect 21729 39383 21787 39389
rect 22002 39380 22008 39432
rect 22060 39380 22066 39432
rect 22278 39380 22284 39432
rect 22336 39380 22342 39432
rect 22554 39380 22560 39432
rect 22612 39380 22618 39432
rect 23400 39429 23428 39460
rect 23017 39423 23075 39429
rect 23017 39389 23029 39423
rect 23063 39389 23075 39423
rect 23017 39383 23075 39389
rect 23385 39423 23443 39429
rect 23385 39389 23397 39423
rect 23431 39389 23443 39423
rect 23385 39383 23443 39389
rect 20496 39256 21036 39284
rect 21085 39287 21143 39293
rect 20496 39244 20502 39256
rect 21085 39253 21097 39287
rect 21131 39284 21143 39287
rect 21450 39284 21456 39296
rect 21131 39256 21456 39284
rect 21131 39253 21143 39256
rect 21085 39247 21143 39253
rect 21450 39244 21456 39256
rect 21508 39244 21514 39296
rect 22097 39287 22155 39293
rect 22097 39253 22109 39287
rect 22143 39284 22155 39287
rect 23032 39284 23060 39383
rect 23842 39380 23848 39432
rect 23900 39380 23906 39432
rect 23934 39380 23940 39432
rect 23992 39380 23998 39432
rect 22143 39256 23060 39284
rect 23661 39287 23719 39293
rect 22143 39253 22155 39256
rect 22097 39247 22155 39253
rect 23661 39253 23673 39287
rect 23707 39284 23719 39287
rect 23934 39284 23940 39296
rect 23707 39256 23940 39284
rect 23707 39253 23719 39256
rect 23661 39247 23719 39253
rect 23934 39244 23940 39256
rect 23992 39244 23998 39296
rect 24121 39287 24179 39293
rect 24121 39253 24133 39287
rect 24167 39284 24179 39287
rect 25222 39284 25228 39296
rect 24167 39256 25228 39284
rect 24167 39253 24179 39256
rect 24121 39247 24179 39253
rect 25222 39244 25228 39256
rect 25280 39244 25286 39296
rect 1104 39194 25000 39216
rect 1104 39142 6884 39194
rect 6936 39142 6948 39194
rect 7000 39142 7012 39194
rect 7064 39142 7076 39194
rect 7128 39142 7140 39194
rect 7192 39142 12818 39194
rect 12870 39142 12882 39194
rect 12934 39142 12946 39194
rect 12998 39142 13010 39194
rect 13062 39142 13074 39194
rect 13126 39142 18752 39194
rect 18804 39142 18816 39194
rect 18868 39142 18880 39194
rect 18932 39142 18944 39194
rect 18996 39142 19008 39194
rect 19060 39142 24686 39194
rect 24738 39142 24750 39194
rect 24802 39142 24814 39194
rect 24866 39142 24878 39194
rect 24930 39142 24942 39194
rect 24994 39142 25000 39194
rect 1104 39120 25000 39142
rect 1486 39040 1492 39092
rect 1544 39040 1550 39092
rect 4154 39040 4160 39092
rect 4212 39080 4218 39092
rect 4890 39080 4896 39092
rect 4212 39052 4896 39080
rect 4212 39040 4218 39052
rect 4890 39040 4896 39052
rect 4948 39040 4954 39092
rect 5350 39040 5356 39092
rect 5408 39040 5414 39092
rect 6362 39040 6368 39092
rect 6420 39080 6426 39092
rect 8018 39080 8024 39092
rect 6420 39052 8024 39080
rect 6420 39040 6426 39052
rect 8018 39040 8024 39052
rect 8076 39040 8082 39092
rect 11698 39080 11704 39092
rect 8312 39052 11704 39080
rect 1504 39012 1532 39040
rect 5368 39012 5396 39040
rect 8312 39024 8340 39052
rect 11698 39040 11704 39052
rect 11756 39040 11762 39092
rect 20438 39040 20444 39092
rect 20496 39040 20502 39092
rect 20717 39083 20775 39089
rect 20717 39049 20729 39083
rect 20763 39080 20775 39083
rect 20898 39080 20904 39092
rect 20763 39052 20904 39080
rect 20763 39049 20775 39052
rect 20717 39043 20775 39049
rect 20898 39040 20904 39052
rect 20956 39040 20962 39092
rect 21450 39040 21456 39092
rect 21508 39080 21514 39092
rect 23385 39083 23443 39089
rect 21508 39052 23152 39080
rect 21508 39040 21514 39052
rect 8294 39012 8300 39024
rect 1504 38984 5396 39012
rect 8036 38984 8300 39012
rect 1854 38944 1860 38956
rect 1688 38916 1860 38944
rect 1688 38885 1716 38916
rect 1854 38904 1860 38916
rect 1912 38904 1918 38956
rect 1947 38947 2005 38953
rect 1947 38913 1959 38947
rect 1993 38944 2005 38947
rect 2866 38944 2872 38956
rect 1993 38916 2872 38944
rect 1993 38913 2005 38916
rect 1947 38907 2005 38913
rect 2866 38904 2872 38916
rect 2924 38904 2930 38956
rect 3050 38904 3056 38956
rect 3108 38904 3114 38956
rect 3418 38904 3424 38956
rect 3476 38944 3482 38956
rect 4065 38947 4123 38953
rect 4065 38944 4077 38947
rect 3476 38916 4077 38944
rect 3476 38904 3482 38916
rect 4065 38913 4077 38916
rect 4111 38913 4123 38947
rect 4617 38947 4675 38953
rect 4617 38944 4629 38947
rect 4065 38907 4123 38913
rect 4172 38916 4629 38944
rect 1673 38879 1731 38885
rect 1673 38845 1685 38879
rect 1719 38845 1731 38879
rect 1673 38839 1731 38845
rect 2682 38836 2688 38888
rect 2740 38836 2746 38888
rect 3510 38836 3516 38888
rect 3568 38876 3574 38888
rect 3789 38879 3847 38885
rect 3789 38876 3801 38879
rect 3568 38848 3801 38876
rect 3568 38836 3574 38848
rect 3789 38845 3801 38848
rect 3835 38845 3847 38879
rect 3789 38839 3847 38845
rect 3878 38836 3884 38888
rect 3936 38876 3942 38888
rect 4172 38876 4200 38916
rect 4617 38913 4629 38916
rect 4663 38913 4675 38947
rect 4617 38907 4675 38913
rect 4893 38947 4951 38953
rect 4893 38913 4905 38947
rect 4939 38944 4951 38947
rect 5258 38944 5264 38956
rect 4939 38916 5264 38944
rect 4939 38913 4951 38916
rect 4893 38907 4951 38913
rect 5258 38904 5264 38916
rect 5316 38904 5322 38956
rect 7374 38904 7380 38956
rect 7432 38904 7438 38956
rect 3936 38848 4200 38876
rect 4341 38879 4399 38885
rect 3936 38836 3942 38848
rect 4341 38845 4353 38879
rect 4387 38876 4399 38879
rect 5902 38876 5908 38888
rect 4387 38848 5908 38876
rect 4387 38845 4399 38848
rect 4341 38839 4399 38845
rect 5902 38836 5908 38848
rect 5960 38876 5966 38888
rect 6822 38876 6828 38888
rect 5960 38848 6828 38876
rect 5960 38836 5966 38848
rect 6822 38836 6828 38848
rect 6880 38836 6886 38888
rect 7392 38876 7420 38904
rect 8036 38876 8064 38984
rect 8294 38972 8300 38984
rect 8352 38972 8358 39024
rect 8662 38972 8668 39024
rect 8720 39012 8726 39024
rect 16482 39012 16488 39024
rect 8720 38984 16488 39012
rect 8720 38972 8726 38984
rect 16482 38972 16488 38984
rect 16540 38972 16546 39024
rect 21174 38972 21180 39024
rect 21232 38972 21238 39024
rect 8386 38944 8392 38956
rect 8347 38916 8392 38944
rect 8386 38904 8392 38916
rect 8444 38944 8450 38956
rect 11759 38947 11817 38953
rect 11759 38944 11771 38947
rect 8444 38916 11771 38944
rect 8444 38904 8450 38916
rect 11759 38913 11771 38916
rect 11805 38913 11817 38947
rect 11759 38907 11817 38913
rect 19242 38904 19248 38956
rect 19300 38904 19306 38956
rect 8113 38879 8171 38885
rect 8113 38876 8125 38879
rect 7392 38848 8125 38876
rect 8113 38845 8125 38848
rect 8159 38845 8171 38879
rect 8113 38839 8171 38845
rect 11514 38836 11520 38888
rect 11572 38836 11578 38888
rect 19260 38876 19288 38904
rect 20622 38888 20628 38940
rect 20680 38888 20686 38940
rect 20898 38904 20904 38956
rect 20956 38904 20962 38956
rect 21192 38944 21220 38972
rect 21637 38947 21695 38953
rect 21637 38944 21649 38947
rect 21192 38916 21649 38944
rect 21637 38913 21649 38916
rect 21683 38944 21695 38947
rect 22077 38947 22135 38953
rect 22077 38944 22089 38947
rect 21683 38916 22089 38944
rect 21683 38913 21695 38916
rect 21637 38907 21695 38913
rect 22077 38913 22089 38916
rect 22123 38913 22135 38947
rect 22077 38907 22135 38913
rect 20438 38876 20444 38888
rect 19260 38848 20444 38876
rect 20438 38836 20444 38848
rect 20496 38836 20502 38888
rect 21818 38836 21824 38888
rect 21876 38836 21882 38888
rect 23124 38876 23152 39052
rect 23385 39049 23397 39083
rect 23431 39049 23443 39083
rect 23385 39043 23443 39049
rect 23661 39083 23719 39089
rect 23661 39049 23673 39083
rect 23707 39080 23719 39083
rect 23842 39080 23848 39092
rect 23707 39052 23848 39080
rect 23707 39049 23719 39052
rect 23661 39043 23719 39049
rect 23400 39012 23428 39043
rect 23842 39040 23848 39052
rect 23900 39040 23906 39092
rect 24121 39015 24179 39021
rect 24121 39012 24133 39015
rect 23400 38984 24133 39012
rect 24121 38981 24133 38984
rect 24167 38981 24179 39015
rect 24121 38975 24179 38981
rect 23566 38904 23572 38956
rect 23624 38904 23630 38956
rect 23658 38904 23664 38956
rect 23716 38944 23722 38956
rect 23845 38947 23903 38953
rect 23845 38944 23857 38947
rect 23716 38916 23857 38944
rect 23716 38904 23722 38916
rect 23845 38913 23857 38916
rect 23891 38913 23903 38947
rect 23845 38907 23903 38913
rect 24026 38904 24032 38956
rect 24084 38904 24090 38956
rect 24044 38876 24072 38904
rect 23124 38848 24072 38876
rect 2700 38749 2728 38836
rect 16666 38768 16672 38820
rect 16724 38808 16730 38820
rect 20070 38808 20076 38820
rect 16724 38780 20076 38808
rect 16724 38768 16730 38780
rect 20070 38768 20076 38780
rect 20128 38768 20134 38820
rect 23201 38811 23259 38817
rect 23201 38777 23213 38811
rect 23247 38808 23259 38811
rect 23474 38808 23480 38820
rect 23247 38780 23480 38808
rect 23247 38777 23259 38780
rect 23201 38771 23259 38777
rect 23474 38768 23480 38780
rect 23532 38768 23538 38820
rect 2685 38743 2743 38749
rect 2685 38709 2697 38743
rect 2731 38709 2743 38743
rect 2685 38703 2743 38709
rect 5258 38700 5264 38752
rect 5316 38740 5322 38752
rect 8570 38740 8576 38752
rect 5316 38712 8576 38740
rect 5316 38700 5322 38712
rect 8570 38700 8576 38712
rect 8628 38700 8634 38752
rect 9122 38700 9128 38752
rect 9180 38700 9186 38752
rect 12526 38700 12532 38752
rect 12584 38700 12590 38752
rect 17126 38700 17132 38752
rect 17184 38740 17190 38752
rect 20898 38740 20904 38752
rect 17184 38712 20904 38740
rect 17184 38700 17190 38712
rect 20898 38700 20904 38712
rect 20956 38700 20962 38752
rect 21453 38743 21511 38749
rect 21453 38709 21465 38743
rect 21499 38740 21511 38743
rect 22094 38740 22100 38752
rect 21499 38712 22100 38740
rect 21499 38709 21511 38712
rect 21453 38703 21511 38709
rect 22094 38700 22100 38712
rect 22152 38700 22158 38752
rect 24394 38700 24400 38752
rect 24452 38700 24458 38752
rect 1104 38650 24840 38672
rect 1104 38598 3917 38650
rect 3969 38598 3981 38650
rect 4033 38598 4045 38650
rect 4097 38598 4109 38650
rect 4161 38598 4173 38650
rect 4225 38598 9851 38650
rect 9903 38598 9915 38650
rect 9967 38598 9979 38650
rect 10031 38598 10043 38650
rect 10095 38598 10107 38650
rect 10159 38598 15785 38650
rect 15837 38598 15849 38650
rect 15901 38598 15913 38650
rect 15965 38598 15977 38650
rect 16029 38598 16041 38650
rect 16093 38598 21719 38650
rect 21771 38598 21783 38650
rect 21835 38598 21847 38650
rect 21899 38598 21911 38650
rect 21963 38598 21975 38650
rect 22027 38598 24840 38650
rect 1104 38576 24840 38598
rect 5258 38536 5264 38548
rect 3804 38508 5264 38536
rect 1854 38292 1860 38344
rect 1912 38332 1918 38344
rect 3804 38341 3832 38508
rect 5258 38496 5264 38508
rect 5316 38496 5322 38548
rect 9214 38536 9220 38548
rect 5368 38508 9220 38536
rect 3789 38335 3847 38341
rect 3789 38332 3801 38335
rect 1912 38304 3801 38332
rect 1912 38292 1918 38304
rect 3789 38301 3801 38304
rect 3835 38301 3847 38335
rect 3789 38295 3847 38301
rect 4047 38305 4105 38311
rect 750 38224 756 38276
rect 808 38264 814 38276
rect 1397 38267 1455 38273
rect 1397 38264 1409 38267
rect 808 38236 1409 38264
rect 808 38224 814 38236
rect 1397 38233 1409 38236
rect 1443 38233 1455 38267
rect 1397 38227 1455 38233
rect 2222 38224 2228 38276
rect 2280 38224 2286 38276
rect 2409 38267 2467 38273
rect 2409 38233 2421 38267
rect 2455 38233 2467 38267
rect 2409 38227 2467 38233
rect 1210 38156 1216 38208
rect 1268 38196 1274 38208
rect 2424 38196 2452 38227
rect 2866 38224 2872 38276
rect 2924 38264 2930 38276
rect 3050 38264 3056 38276
rect 2924 38236 3056 38264
rect 2924 38224 2930 38236
rect 3050 38224 3056 38236
rect 3108 38264 3114 38276
rect 3145 38267 3203 38273
rect 3145 38264 3157 38267
rect 3108 38236 3157 38264
rect 3108 38224 3114 38236
rect 3145 38233 3157 38236
rect 3191 38233 3203 38267
rect 4047 38271 4059 38305
rect 4093 38302 4105 38305
rect 4093 38271 4106 38302
rect 5074 38292 5080 38344
rect 5132 38292 5138 38344
rect 5368 38341 5396 38508
rect 9214 38496 9220 38508
rect 9272 38496 9278 38548
rect 11698 38496 11704 38548
rect 11756 38536 11762 38548
rect 12526 38536 12532 38548
rect 11756 38508 12020 38536
rect 11756 38496 11762 38508
rect 5994 38428 6000 38480
rect 6052 38428 6058 38480
rect 11330 38428 11336 38480
rect 11388 38428 11394 38480
rect 11882 38428 11888 38480
rect 11940 38428 11946 38480
rect 6390 38403 6448 38409
rect 6390 38400 6402 38403
rect 5460 38372 6402 38400
rect 5353 38335 5411 38341
rect 5353 38301 5365 38335
rect 5399 38301 5411 38335
rect 5353 38295 5411 38301
rect 4047 38265 4106 38271
rect 4078 38264 4106 38265
rect 5092 38264 5120 38292
rect 5460 38264 5488 38372
rect 6390 38369 6402 38372
rect 6436 38369 6448 38403
rect 6390 38363 6448 38369
rect 8294 38360 8300 38412
rect 8352 38400 8358 38412
rect 8662 38400 8668 38412
rect 8352 38372 8668 38400
rect 8352 38360 8358 38372
rect 8662 38360 8668 38372
rect 8720 38400 8726 38412
rect 9125 38403 9183 38409
rect 9125 38400 9137 38403
rect 8720 38372 9137 38400
rect 8720 38360 8726 38372
rect 9125 38369 9137 38372
rect 9171 38369 9183 38403
rect 11348 38400 11376 38428
rect 9125 38363 9183 38369
rect 9784 38372 11376 38400
rect 11609 38403 11667 38409
rect 5534 38292 5540 38344
rect 5592 38292 5598 38344
rect 6270 38292 6276 38344
rect 6328 38292 6334 38344
rect 6546 38292 6552 38344
rect 6604 38292 6610 38344
rect 7650 38292 7656 38344
rect 7708 38332 7714 38344
rect 9399 38335 9457 38341
rect 9399 38332 9411 38335
rect 7708 38304 9411 38332
rect 7708 38292 7714 38304
rect 9399 38301 9411 38304
rect 9445 38332 9457 38335
rect 9490 38332 9496 38344
rect 9445 38304 9496 38332
rect 9445 38301 9457 38304
rect 9399 38295 9457 38301
rect 9490 38292 9496 38304
rect 9548 38292 9554 38344
rect 4078 38236 4936 38264
rect 5092 38236 5488 38264
rect 7024 38236 7604 38264
rect 3145 38227 3203 38233
rect 1268 38168 2452 38196
rect 1268 38156 1274 38168
rect 4798 38156 4804 38208
rect 4856 38156 4862 38208
rect 4908 38196 4936 38236
rect 5350 38196 5356 38208
rect 4908 38168 5356 38196
rect 5350 38156 5356 38168
rect 5408 38156 5414 38208
rect 6822 38156 6828 38208
rect 6880 38196 6886 38208
rect 7024 38196 7052 38236
rect 6880 38168 7052 38196
rect 7193 38199 7251 38205
rect 6880 38156 6886 38168
rect 7193 38165 7205 38199
rect 7239 38196 7251 38199
rect 7466 38196 7472 38208
rect 7239 38168 7472 38196
rect 7239 38165 7251 38168
rect 7193 38159 7251 38165
rect 7466 38156 7472 38168
rect 7524 38156 7530 38208
rect 7576 38196 7604 38236
rect 7926 38224 7932 38276
rect 7984 38264 7990 38276
rect 9784 38264 9812 38372
rect 11609 38369 11621 38403
rect 11655 38400 11667 38403
rect 11900 38400 11928 38428
rect 11992 38412 12020 38508
rect 12084 38508 12532 38536
rect 12084 38477 12112 38508
rect 12526 38496 12532 38508
rect 12584 38496 12590 38548
rect 13262 38496 13268 38548
rect 13320 38496 13326 38548
rect 19889 38539 19947 38545
rect 19889 38505 19901 38539
rect 19935 38536 19947 38539
rect 20622 38536 20628 38548
rect 19935 38508 20628 38536
rect 19935 38505 19947 38508
rect 19889 38499 19947 38505
rect 20622 38496 20628 38508
rect 20680 38496 20686 38548
rect 21082 38496 21088 38548
rect 21140 38536 21146 38548
rect 22465 38539 22523 38545
rect 22465 38536 22477 38539
rect 21140 38508 22477 38536
rect 21140 38496 21146 38508
rect 22465 38505 22477 38508
rect 22511 38505 22523 38539
rect 22465 38499 22523 38505
rect 22922 38496 22928 38548
rect 22980 38536 22986 38548
rect 23293 38539 23351 38545
rect 23293 38536 23305 38539
rect 22980 38508 23305 38536
rect 22980 38496 22986 38508
rect 23293 38505 23305 38508
rect 23339 38505 23351 38539
rect 23293 38499 23351 38505
rect 23566 38496 23572 38548
rect 23624 38536 23630 38548
rect 23661 38539 23719 38545
rect 23661 38536 23673 38539
rect 23624 38508 23673 38536
rect 23624 38496 23630 38508
rect 23661 38505 23673 38508
rect 23707 38505 23719 38539
rect 23661 38499 23719 38505
rect 23750 38496 23756 38548
rect 23808 38496 23814 38548
rect 12069 38471 12127 38477
rect 12069 38437 12081 38471
rect 12115 38437 12127 38471
rect 12069 38431 12127 38437
rect 20714 38428 20720 38480
rect 20772 38468 20778 38480
rect 22738 38468 22744 38480
rect 20772 38440 22744 38468
rect 20772 38428 20778 38440
rect 22738 38428 22744 38440
rect 22796 38428 22802 38480
rect 23017 38471 23075 38477
rect 23017 38437 23029 38471
rect 23063 38468 23075 38471
rect 23768 38468 23796 38496
rect 23063 38440 23796 38468
rect 23063 38437 23075 38440
rect 23017 38431 23075 38437
rect 11655 38372 11928 38400
rect 11655 38369 11667 38372
rect 11609 38363 11667 38369
rect 11974 38360 11980 38412
rect 12032 38400 12038 38412
rect 12462 38403 12520 38409
rect 12462 38400 12474 38403
rect 12032 38372 12474 38400
rect 12032 38360 12038 38372
rect 12462 38369 12474 38372
rect 12508 38369 12520 38403
rect 12462 38363 12520 38369
rect 23106 38360 23112 38412
rect 23164 38400 23170 38412
rect 23164 38372 23888 38400
rect 23164 38360 23170 38372
rect 11330 38292 11336 38344
rect 11388 38332 11394 38344
rect 11425 38335 11483 38341
rect 11425 38332 11437 38335
rect 11388 38304 11437 38332
rect 11388 38292 11394 38304
rect 11425 38301 11437 38304
rect 11471 38301 11483 38335
rect 11425 38295 11483 38301
rect 12342 38292 12348 38344
rect 12400 38292 12406 38344
rect 12618 38292 12624 38344
rect 12676 38292 12682 38344
rect 20073 38335 20131 38341
rect 20073 38301 20085 38335
rect 20119 38301 20131 38335
rect 20073 38295 20131 38301
rect 7984 38236 9812 38264
rect 9876 38236 10272 38264
rect 7984 38224 7990 38236
rect 9876 38196 9904 38236
rect 7576 38168 9904 38196
rect 10134 38156 10140 38208
rect 10192 38156 10198 38208
rect 10244 38196 10272 38236
rect 20088 38196 20116 38295
rect 22094 38292 22100 38344
rect 22152 38292 22158 38344
rect 22646 38292 22652 38344
rect 22704 38292 22710 38344
rect 22741 38335 22799 38341
rect 22741 38301 22753 38335
rect 22787 38332 22799 38335
rect 22787 38304 22876 38332
rect 22787 38301 22799 38304
rect 22741 38295 22799 38301
rect 22848 38208 22876 38304
rect 22922 38292 22928 38344
rect 22980 38292 22986 38344
rect 23201 38335 23259 38341
rect 23201 38322 23213 38335
rect 23124 38301 23213 38322
rect 23247 38301 23259 38335
rect 23124 38295 23259 38301
rect 23124 38294 23244 38295
rect 23014 38224 23020 38276
rect 23072 38264 23078 38276
rect 23124 38264 23152 38294
rect 23474 38292 23480 38344
rect 23532 38292 23538 38344
rect 23860 38341 23888 38372
rect 23845 38335 23903 38341
rect 23845 38301 23857 38335
rect 23891 38301 23903 38335
rect 23845 38295 23903 38301
rect 23934 38292 23940 38344
rect 23992 38292 23998 38344
rect 23072 38236 23152 38264
rect 23072 38224 23078 38236
rect 10244 38168 20116 38196
rect 22186 38156 22192 38208
rect 22244 38156 22250 38208
rect 22830 38156 22836 38208
rect 22888 38156 22894 38208
rect 22922 38156 22928 38208
rect 22980 38156 22986 38208
rect 24121 38199 24179 38205
rect 24121 38165 24133 38199
rect 24167 38196 24179 38199
rect 25222 38196 25228 38208
rect 24167 38168 25228 38196
rect 24167 38165 24179 38168
rect 24121 38159 24179 38165
rect 25222 38156 25228 38168
rect 25280 38156 25286 38208
rect 1104 38106 25000 38128
rect 1104 38054 6884 38106
rect 6936 38054 6948 38106
rect 7000 38054 7012 38106
rect 7064 38054 7076 38106
rect 7128 38054 7140 38106
rect 7192 38054 12818 38106
rect 12870 38054 12882 38106
rect 12934 38054 12946 38106
rect 12998 38054 13010 38106
rect 13062 38054 13074 38106
rect 13126 38054 18752 38106
rect 18804 38054 18816 38106
rect 18868 38054 18880 38106
rect 18932 38054 18944 38106
rect 18996 38054 19008 38106
rect 19060 38054 24686 38106
rect 24738 38054 24750 38106
rect 24802 38054 24814 38106
rect 24866 38054 24878 38106
rect 24930 38054 24942 38106
rect 24994 38054 25000 38106
rect 1104 38032 25000 38054
rect 4798 37992 4804 38004
rect 3896 37964 4804 37992
rect 1673 37927 1731 37933
rect 1673 37893 1685 37927
rect 1719 37924 1731 37927
rect 2038 37924 2044 37936
rect 1719 37896 2044 37924
rect 1719 37893 1731 37896
rect 1673 37887 1731 37893
rect 2038 37884 2044 37896
rect 2096 37884 2102 37936
rect 3510 37884 3516 37936
rect 3568 37884 3574 37936
rect 3896 37933 3924 37964
rect 4798 37952 4804 37964
rect 4856 37952 4862 38004
rect 6546 37952 6552 38004
rect 6604 37992 6610 38004
rect 7377 37995 7435 38001
rect 7377 37992 7389 37995
rect 6604 37964 7389 37992
rect 6604 37952 6610 37964
rect 7377 37961 7389 37964
rect 7423 37961 7435 37995
rect 7377 37955 7435 37961
rect 8294 37952 8300 38004
rect 8352 37992 8358 38004
rect 8938 37992 8944 38004
rect 8352 37964 8944 37992
rect 8352 37952 8358 37964
rect 8938 37952 8944 37964
rect 8996 37952 9002 38004
rect 10134 37992 10140 38004
rect 9324 37964 10140 37992
rect 3881 37927 3939 37933
rect 3881 37893 3893 37927
rect 3927 37893 3939 37927
rect 4522 37924 4528 37936
rect 3881 37887 3939 37893
rect 4264 37896 4528 37924
rect 1394 37816 1400 37868
rect 1452 37816 1458 37868
rect 2191 37859 2249 37865
rect 2191 37856 2203 37859
rect 1504 37828 2203 37856
rect 1118 37748 1124 37800
rect 1176 37788 1182 37800
rect 1504 37788 1532 37828
rect 2191 37825 2203 37828
rect 2237 37825 2249 37859
rect 2191 37819 2249 37825
rect 3602 37816 3608 37868
rect 3660 37856 3666 37868
rect 3789 37859 3847 37865
rect 3789 37856 3801 37859
rect 3660 37828 3801 37856
rect 3660 37816 3666 37828
rect 3789 37825 3801 37828
rect 3835 37856 3847 37859
rect 4154 37856 4160 37868
rect 3835 37828 4160 37856
rect 3835 37825 3847 37828
rect 3789 37819 3847 37825
rect 4154 37816 4160 37828
rect 4212 37816 4218 37868
rect 4264 37865 4292 37896
rect 4522 37884 4528 37896
rect 4580 37884 4586 37936
rect 4617 37927 4675 37933
rect 4617 37893 4629 37927
rect 4663 37893 4675 37927
rect 4617 37887 4675 37893
rect 5813 37927 5871 37933
rect 5813 37893 5825 37927
rect 5859 37924 5871 37927
rect 7834 37924 7840 37936
rect 5859 37896 7840 37924
rect 5859 37893 5871 37896
rect 5813 37887 5871 37893
rect 4249 37859 4307 37865
rect 4249 37825 4261 37859
rect 4295 37825 4307 37859
rect 4632 37856 4660 37887
rect 7834 37884 7840 37896
rect 7892 37884 7898 37936
rect 8110 37884 8116 37936
rect 8168 37924 8174 37936
rect 8754 37924 8760 37936
rect 8168 37896 8760 37924
rect 8168 37884 8174 37896
rect 8754 37884 8760 37896
rect 8812 37884 8818 37936
rect 9214 37884 9220 37936
rect 9272 37884 9278 37936
rect 9324 37933 9352 37964
rect 10134 37952 10140 37964
rect 10192 37952 10198 38004
rect 11974 37952 11980 38004
rect 12032 37992 12038 38004
rect 12342 37992 12348 38004
rect 12032 37964 12348 37992
rect 12032 37952 12038 37964
rect 12342 37952 12348 37964
rect 12400 37952 12406 38004
rect 12618 37952 12624 38004
rect 12676 37992 12682 38004
rect 13081 37995 13139 38001
rect 13081 37992 13093 37995
rect 12676 37964 13093 37992
rect 12676 37952 12682 37964
rect 13081 37961 13093 37964
rect 13127 37961 13139 37995
rect 13081 37955 13139 37961
rect 20162 37952 20168 38004
rect 20220 37992 20226 38004
rect 21453 37995 21511 38001
rect 21453 37992 21465 37995
rect 20220 37964 21465 37992
rect 20220 37952 20226 37964
rect 21453 37961 21465 37964
rect 21499 37961 21511 37995
rect 21453 37955 21511 37961
rect 22186 37952 22192 38004
rect 22244 37992 22250 38004
rect 22244 37964 22692 37992
rect 22244 37952 22250 37964
rect 9309 37927 9367 37933
rect 9309 37893 9321 37927
rect 9355 37893 9367 37927
rect 9309 37887 9367 37893
rect 9490 37884 9496 37936
rect 9548 37924 9554 37936
rect 22554 37924 22560 37936
rect 9548 37896 12296 37924
rect 9548 37884 9554 37896
rect 4798 37856 4804 37868
rect 4632 37828 4804 37856
rect 4249 37819 4307 37825
rect 4798 37816 4804 37828
rect 4856 37816 4862 37868
rect 4982 37816 4988 37868
rect 5040 37816 5046 37868
rect 5537 37859 5595 37865
rect 5537 37856 5549 37859
rect 5092 37828 5549 37856
rect 1176 37760 1532 37788
rect 1176 37748 1182 37760
rect 1854 37748 1860 37800
rect 1912 37788 1918 37800
rect 1949 37791 2007 37797
rect 1949 37788 1961 37791
rect 1912 37760 1961 37788
rect 1912 37748 1918 37760
rect 1949 37757 1961 37760
rect 1995 37757 2007 37791
rect 1949 37751 2007 37757
rect 2976 37760 3358 37788
rect 2976 37729 3004 37760
rect 4890 37748 4896 37800
rect 4948 37788 4954 37800
rect 5092 37788 5120 37828
rect 5537 37825 5549 37828
rect 5583 37825 5595 37859
rect 5537 37819 5595 37825
rect 6639 37859 6697 37865
rect 6639 37825 6651 37859
rect 6685 37856 6697 37859
rect 7558 37856 7564 37868
rect 6685 37828 7564 37856
rect 6685 37825 6697 37828
rect 6639 37819 6697 37825
rect 7558 37816 7564 37828
rect 7616 37816 7622 37868
rect 8772 37856 8800 37884
rect 9674 37856 9680 37868
rect 8772 37828 9680 37856
rect 9674 37816 9680 37828
rect 9732 37816 9738 37868
rect 9766 37816 9772 37868
rect 9824 37856 9830 37868
rect 10059 37859 10117 37865
rect 10059 37856 10071 37859
rect 9824 37828 10071 37856
rect 9824 37816 9830 37828
rect 10059 37825 10071 37828
rect 10105 37825 10117 37859
rect 10059 37819 10117 37825
rect 11514 37816 11520 37868
rect 11572 37856 11578 37868
rect 12069 37859 12127 37865
rect 12069 37856 12081 37859
rect 11572 37828 12081 37856
rect 11572 37816 11578 37828
rect 12069 37825 12081 37828
rect 12115 37825 12127 37859
rect 12268 37856 12296 37896
rect 21836 37896 22560 37924
rect 12343 37859 12401 37865
rect 12343 37856 12355 37859
rect 12268 37828 12355 37856
rect 12069 37819 12127 37825
rect 12343 37825 12355 37828
rect 12389 37856 12401 37859
rect 13630 37856 13636 37868
rect 12389 37828 13636 37856
rect 12389 37825 12401 37828
rect 12343 37819 12401 37825
rect 4948 37760 5120 37788
rect 5261 37791 5319 37797
rect 4948 37748 4954 37760
rect 5261 37757 5273 37791
rect 5307 37757 5319 37791
rect 5261 37751 5319 37757
rect 2961 37723 3019 37729
rect 2961 37689 2973 37723
rect 3007 37689 3019 37723
rect 5276 37720 5304 37751
rect 6086 37748 6092 37800
rect 6144 37788 6150 37800
rect 6365 37791 6423 37797
rect 6365 37788 6377 37791
rect 6144 37760 6377 37788
rect 6144 37748 6150 37760
rect 6365 37757 6377 37760
rect 6411 37757 6423 37791
rect 6365 37751 6423 37757
rect 9122 37748 9128 37800
rect 9180 37748 9186 37800
rect 5276 37692 6500 37720
rect 2961 37683 3019 37689
rect 4801 37655 4859 37661
rect 4801 37621 4813 37655
rect 4847 37652 4859 37655
rect 5258 37652 5264 37664
rect 4847 37624 5264 37652
rect 4847 37621 4859 37624
rect 4801 37615 4859 37621
rect 5258 37612 5264 37624
rect 5316 37652 5322 37664
rect 6270 37652 6276 37664
rect 5316 37624 6276 37652
rect 5316 37612 5322 37624
rect 6270 37612 6276 37624
rect 6328 37612 6334 37664
rect 6472 37652 6500 37692
rect 7374 37652 7380 37664
rect 6472 37624 7380 37652
rect 7374 37612 7380 37624
rect 7432 37612 7438 37664
rect 8662 37612 8668 37664
rect 8720 37652 8726 37664
rect 8938 37652 8944 37664
rect 8720 37624 8944 37652
rect 8720 37612 8726 37624
rect 8938 37612 8944 37624
rect 8996 37612 9002 37664
rect 10229 37655 10287 37661
rect 10229 37621 10241 37655
rect 10275 37652 10287 37655
rect 10594 37652 10600 37664
rect 10275 37624 10600 37652
rect 10275 37621 10287 37624
rect 10229 37615 10287 37621
rect 10594 37612 10600 37624
rect 10652 37612 10658 37664
rect 12084 37652 12112 37819
rect 13630 37816 13636 37828
rect 13688 37816 13694 37868
rect 15286 37816 15292 37868
rect 15344 37856 15350 37868
rect 21637 37859 21695 37865
rect 21637 37856 21649 37859
rect 15344 37828 21649 37856
rect 15344 37816 15350 37828
rect 21637 37825 21649 37828
rect 21683 37825 21695 37859
rect 21637 37819 21695 37825
rect 20254 37788 20260 37800
rect 14108 37760 20260 37788
rect 14108 37664 14136 37760
rect 20254 37748 20260 37760
rect 20312 37788 20318 37800
rect 21836 37797 21864 37896
rect 22554 37884 22560 37896
rect 22612 37884 22618 37936
rect 22095 37859 22153 37865
rect 22095 37825 22107 37859
rect 22141 37856 22153 37859
rect 22664 37856 22692 37964
rect 22738 37952 22744 38004
rect 22796 37952 22802 38004
rect 22922 37952 22928 38004
rect 22980 37992 22986 38004
rect 23845 37995 23903 38001
rect 22980 37964 23796 37992
rect 22980 37952 22986 37964
rect 22756 37924 22784 37952
rect 23768 37933 23796 37964
rect 23845 37961 23857 37995
rect 23891 37961 23903 37995
rect 23845 37955 23903 37961
rect 23753 37927 23811 37933
rect 22756 37896 23520 37924
rect 23385 37859 23443 37865
rect 23385 37856 23397 37859
rect 22141 37828 22600 37856
rect 22664 37828 23397 37856
rect 22141 37825 22153 37828
rect 22095 37819 22153 37825
rect 21821 37791 21879 37797
rect 21821 37788 21833 37791
rect 20312 37760 21833 37788
rect 20312 37748 20318 37760
rect 21821 37757 21833 37760
rect 21867 37757 21879 37791
rect 22572 37788 22600 37828
rect 23385 37825 23397 37828
rect 23431 37825 23443 37859
rect 23492 37856 23520 37896
rect 23753 37893 23765 37927
rect 23799 37893 23811 37927
rect 23753 37887 23811 37893
rect 23860 37856 23888 37955
rect 23492 37828 23888 37856
rect 23385 37819 23443 37825
rect 24026 37816 24032 37868
rect 24084 37816 24090 37868
rect 24213 37859 24271 37865
rect 24213 37825 24225 37859
rect 24259 37825 24271 37859
rect 24213 37819 24271 37825
rect 22922 37788 22928 37800
rect 22572 37760 22928 37788
rect 21821 37751 21879 37757
rect 22922 37748 22928 37760
rect 22980 37748 22986 37800
rect 23201 37791 23259 37797
rect 23201 37757 23213 37791
rect 23247 37757 23259 37791
rect 24228 37788 24256 37819
rect 23201 37751 23259 37757
rect 23308 37760 24256 37788
rect 22830 37680 22836 37732
rect 22888 37720 22894 37732
rect 23216 37720 23244 37751
rect 22888 37692 23244 37720
rect 22888 37680 22894 37692
rect 14090 37652 14096 37664
rect 12084 37624 14096 37652
rect 14090 37612 14096 37624
rect 14148 37612 14154 37664
rect 21634 37612 21640 37664
rect 21692 37652 21698 37664
rect 23308 37652 23336 37760
rect 23661 37723 23719 37729
rect 23661 37689 23673 37723
rect 23707 37720 23719 37723
rect 23707 37692 25452 37720
rect 23707 37689 23719 37692
rect 23661 37683 23719 37689
rect 25424 37664 25452 37692
rect 21692 37624 23336 37652
rect 21692 37612 21698 37624
rect 24394 37612 24400 37664
rect 24452 37612 24458 37664
rect 25406 37612 25412 37664
rect 25464 37612 25470 37664
rect 1104 37562 24840 37584
rect 1104 37510 3917 37562
rect 3969 37510 3981 37562
rect 4033 37510 4045 37562
rect 4097 37510 4109 37562
rect 4161 37510 4173 37562
rect 4225 37510 9851 37562
rect 9903 37510 9915 37562
rect 9967 37510 9979 37562
rect 10031 37510 10043 37562
rect 10095 37510 10107 37562
rect 10159 37510 15785 37562
rect 15837 37510 15849 37562
rect 15901 37510 15913 37562
rect 15965 37510 15977 37562
rect 16029 37510 16041 37562
rect 16093 37510 21719 37562
rect 21771 37510 21783 37562
rect 21835 37510 21847 37562
rect 21899 37510 21911 37562
rect 21963 37510 21975 37562
rect 22027 37510 24840 37562
rect 1104 37488 24840 37510
rect 3878 37408 3884 37460
rect 3936 37448 3942 37460
rect 4982 37448 4988 37460
rect 3936 37420 4988 37448
rect 3936 37408 3942 37420
rect 4982 37408 4988 37420
rect 5040 37408 5046 37460
rect 5626 37408 5632 37460
rect 5684 37448 5690 37460
rect 6546 37448 6552 37460
rect 5684 37420 6552 37448
rect 5684 37408 5690 37420
rect 6546 37408 6552 37420
rect 6604 37448 6610 37460
rect 6604 37420 16252 37448
rect 6604 37408 6610 37420
rect 7374 37340 7380 37392
rect 7432 37380 7438 37392
rect 8110 37380 8116 37392
rect 7432 37352 8116 37380
rect 7432 37340 7438 37352
rect 8110 37340 8116 37352
rect 8168 37380 8174 37392
rect 16224 37380 16252 37420
rect 21634 37408 21640 37460
rect 21692 37408 21698 37460
rect 21913 37451 21971 37457
rect 21913 37417 21925 37451
rect 21959 37448 21971 37451
rect 22557 37451 22615 37457
rect 21959 37420 22232 37448
rect 21959 37417 21971 37420
rect 21913 37411 21971 37417
rect 22204 37380 22232 37420
rect 22557 37417 22569 37451
rect 22603 37448 22615 37451
rect 22646 37448 22652 37460
rect 22603 37420 22652 37448
rect 22603 37417 22615 37420
rect 22557 37411 22615 37417
rect 22646 37408 22652 37420
rect 22704 37408 22710 37460
rect 22833 37451 22891 37457
rect 22833 37417 22845 37451
rect 22879 37448 22891 37451
rect 23106 37448 23112 37460
rect 22879 37420 23112 37448
rect 22879 37417 22891 37420
rect 22833 37411 22891 37417
rect 23106 37408 23112 37420
rect 23164 37408 23170 37460
rect 23014 37380 23020 37392
rect 8168 37352 9674 37380
rect 16224 37352 22048 37380
rect 22204 37352 23020 37380
rect 8168 37340 8174 37352
rect 1946 37272 1952 37324
rect 2004 37312 2010 37324
rect 8205 37315 8263 37321
rect 2004 37284 3832 37312
rect 2004 37272 2010 37284
rect 2501 37247 2559 37253
rect 2501 37213 2513 37247
rect 2547 37244 2559 37247
rect 2866 37244 2872 37256
rect 2547 37216 2872 37244
rect 2547 37213 2559 37216
rect 2501 37207 2559 37213
rect 2866 37204 2872 37216
rect 2924 37204 2930 37256
rect 3804 37253 3832 37284
rect 8205 37281 8217 37315
rect 8251 37312 8263 37315
rect 8389 37315 8447 37321
rect 8389 37312 8401 37315
rect 8251 37284 8401 37312
rect 8251 37281 8263 37284
rect 8205 37275 8263 37281
rect 8389 37281 8401 37284
rect 8435 37281 8447 37315
rect 8389 37275 8447 37281
rect 3789 37247 3847 37253
rect 3789 37213 3801 37247
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 4709 37247 4767 37253
rect 4709 37213 4721 37247
rect 4755 37213 4767 37247
rect 4982 37244 4988 37256
rect 4943 37216 4988 37244
rect 4709 37207 4767 37213
rect 1397 37179 1455 37185
rect 1397 37145 1409 37179
rect 1443 37176 1455 37179
rect 1486 37176 1492 37188
rect 1443 37148 1492 37176
rect 1443 37145 1455 37148
rect 1397 37139 1455 37145
rect 1486 37136 1492 37148
rect 1544 37136 1550 37188
rect 2222 37136 2228 37188
rect 2280 37136 2286 37188
rect 2774 37136 2780 37188
rect 2832 37136 2838 37188
rect 3145 37179 3203 37185
rect 3145 37176 3157 37179
rect 2884 37148 3157 37176
rect 1670 37068 1676 37120
rect 1728 37108 1734 37120
rect 2884 37108 2912 37148
rect 3145 37145 3157 37148
rect 3191 37145 3203 37179
rect 4062 37176 4068 37188
rect 3145 37139 3203 37145
rect 3344 37148 4068 37176
rect 1728 37080 2912 37108
rect 1728 37068 1734 37080
rect 2958 37068 2964 37120
rect 3016 37108 3022 37120
rect 3344 37108 3372 37148
rect 4062 37136 4068 37148
rect 4120 37136 4126 37188
rect 4724 37176 4752 37207
rect 4982 37204 4988 37216
rect 5040 37244 5046 37256
rect 5350 37244 5356 37256
rect 5040 37216 5356 37244
rect 5040 37204 5046 37216
rect 5350 37204 5356 37216
rect 5408 37204 5414 37256
rect 5718 37204 5724 37256
rect 5776 37204 5782 37256
rect 6549 37247 6607 37253
rect 6549 37213 6561 37247
rect 6595 37213 6607 37247
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 6549 37207 6607 37213
rect 6807 37217 6865 37223
rect 5736 37176 5764 37204
rect 6564 37176 6592 37207
rect 6807 37183 6819 37217
rect 6853 37214 6865 37217
rect 7576 37216 7941 37244
rect 6853 37183 6868 37214
rect 6807 37177 6868 37183
rect 4724 37148 6592 37176
rect 3016 37080 3372 37108
rect 3016 37068 3022 37080
rect 3418 37068 3424 37120
rect 3476 37108 3482 37120
rect 4614 37108 4620 37120
rect 3476 37080 4620 37108
rect 3476 37068 3482 37080
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 5442 37068 5448 37120
rect 5500 37108 5506 37120
rect 5721 37111 5779 37117
rect 5721 37108 5733 37111
rect 5500 37080 5733 37108
rect 5500 37068 5506 37080
rect 5721 37077 5733 37080
rect 5767 37077 5779 37111
rect 5721 37071 5779 37077
rect 5902 37068 5908 37120
rect 5960 37108 5966 37120
rect 6840 37108 6868 37177
rect 7576 37117 7604 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 7929 37207 7987 37213
rect 7944 37176 7972 37207
rect 8018 37204 8024 37256
rect 8076 37204 8082 37256
rect 8297 37247 8355 37253
rect 8297 37213 8309 37247
rect 8343 37213 8355 37247
rect 8297 37207 8355 37213
rect 8312 37176 8340 37207
rect 8478 37204 8484 37256
rect 8536 37204 8542 37256
rect 9030 37204 9036 37256
rect 9088 37204 9094 37256
rect 7944 37148 8340 37176
rect 5960 37080 6868 37108
rect 7561 37111 7619 37117
rect 5960 37068 5966 37080
rect 7561 37077 7573 37111
rect 7607 37077 7619 37111
rect 7561 37071 7619 37077
rect 8205 37111 8263 37117
rect 8205 37077 8217 37111
rect 8251 37108 8263 37111
rect 9048 37108 9076 37204
rect 8251 37080 9076 37108
rect 9646 37108 9674 37352
rect 10704 37284 10916 37312
rect 10042 37204 10048 37256
rect 10100 37204 10106 37256
rect 10704 37244 10732 37284
rect 10318 37223 10732 37244
rect 10303 37217 10732 37223
rect 10303 37214 10315 37217
rect 9766 37136 9772 37188
rect 9824 37176 9830 37188
rect 10302 37183 10315 37214
rect 10349 37216 10732 37217
rect 10888 37244 10916 37284
rect 16390 37272 16396 37324
rect 16448 37312 16454 37324
rect 16758 37312 16764 37324
rect 16448 37284 16764 37312
rect 16448 37272 16454 37284
rect 16758 37272 16764 37284
rect 16816 37272 16822 37324
rect 18506 37272 18512 37324
rect 18564 37312 18570 37324
rect 19334 37312 19340 37324
rect 18564 37284 19340 37312
rect 18564 37272 18570 37284
rect 19334 37272 19340 37284
rect 19392 37272 19398 37324
rect 22020 37312 22048 37352
rect 23014 37340 23020 37352
rect 23072 37340 23078 37392
rect 22278 37312 22284 37324
rect 20456 37284 20852 37312
rect 14366 37244 14372 37256
rect 10888 37216 14372 37244
rect 10349 37183 10361 37216
rect 14366 37204 14372 37216
rect 14424 37204 14430 37256
rect 17218 37204 17224 37256
rect 17276 37244 17282 37256
rect 20456 37244 20484 37284
rect 17276 37216 20484 37244
rect 17276 37204 17282 37216
rect 20714 37204 20720 37256
rect 20772 37204 20778 37256
rect 20824 37244 20852 37284
rect 21744 37284 21956 37312
rect 22020 37284 22284 37312
rect 21744 37244 21772 37284
rect 20824 37216 21772 37244
rect 21818 37204 21824 37256
rect 21876 37204 21882 37256
rect 10302 37177 10361 37183
rect 10302 37176 10330 37177
rect 21928 37176 21956 37284
rect 22278 37272 22284 37284
rect 22336 37272 22342 37324
rect 22664 37284 22876 37312
rect 22094 37204 22100 37256
rect 22152 37204 22158 37256
rect 22186 37204 22192 37256
rect 22244 37244 22250 37256
rect 22664 37244 22692 37284
rect 22244 37216 22692 37244
rect 22244 37204 22250 37216
rect 22738 37204 22744 37256
rect 22796 37204 22802 37256
rect 22848 37244 22876 37284
rect 24118 37272 24124 37324
rect 24176 37272 24182 37324
rect 23017 37247 23075 37253
rect 23017 37244 23029 37247
rect 22848 37216 23029 37244
rect 23017 37213 23029 37216
rect 23063 37213 23075 37247
rect 23293 37247 23351 37253
rect 23293 37244 23305 37247
rect 23017 37207 23075 37213
rect 23124 37216 23305 37244
rect 23124 37176 23152 37216
rect 23293 37213 23305 37216
rect 23339 37213 23351 37247
rect 23293 37207 23351 37213
rect 23566 37204 23572 37256
rect 23624 37204 23630 37256
rect 23658 37204 23664 37256
rect 23716 37204 23722 37256
rect 23934 37204 23940 37256
rect 23992 37204 23998 37256
rect 23676 37176 23704 37204
rect 9824 37148 10330 37176
rect 10888 37148 21772 37176
rect 21928 37148 23152 37176
rect 23308 37148 23704 37176
rect 9824 37136 9830 37148
rect 10888 37108 10916 37148
rect 9646 37080 10916 37108
rect 8251 37077 8263 37080
rect 8205 37071 8263 37077
rect 11054 37068 11060 37120
rect 11112 37068 11118 37120
rect 11238 37068 11244 37120
rect 11296 37108 11302 37120
rect 18138 37108 18144 37120
rect 11296 37080 18144 37108
rect 11296 37068 11302 37080
rect 18138 37068 18144 37080
rect 18196 37068 18202 37120
rect 20530 37068 20536 37120
rect 20588 37068 20594 37120
rect 21744 37108 21772 37148
rect 22186 37108 22192 37120
rect 21744 37080 22192 37108
rect 22186 37068 22192 37080
rect 22244 37068 22250 37120
rect 23109 37111 23167 37117
rect 23109 37077 23121 37111
rect 23155 37108 23167 37111
rect 23308 37108 23336 37148
rect 23842 37136 23848 37188
rect 23900 37136 23906 37188
rect 23155 37080 23336 37108
rect 23385 37111 23443 37117
rect 23155 37077 23167 37080
rect 23109 37071 23167 37077
rect 23385 37077 23397 37111
rect 23431 37108 23443 37111
rect 23952 37108 23980 37204
rect 23431 37080 23980 37108
rect 23431 37077 23443 37080
rect 23385 37071 23443 37077
rect 1104 37018 25000 37040
rect 1104 36966 6884 37018
rect 6936 36966 6948 37018
rect 7000 36966 7012 37018
rect 7064 36966 7076 37018
rect 7128 36966 7140 37018
rect 7192 36966 12818 37018
rect 12870 36966 12882 37018
rect 12934 36966 12946 37018
rect 12998 36966 13010 37018
rect 13062 36966 13074 37018
rect 13126 36966 18752 37018
rect 18804 36966 18816 37018
rect 18868 36966 18880 37018
rect 18932 36966 18944 37018
rect 18996 36966 19008 37018
rect 19060 36966 24686 37018
rect 24738 36966 24750 37018
rect 24802 36966 24814 37018
rect 24866 36966 24878 37018
rect 24930 36966 24942 37018
rect 24994 36966 25000 37018
rect 1104 36944 25000 36966
rect 5905 36907 5963 36913
rect 5905 36904 5917 36907
rect 3804 36876 5917 36904
rect 1581 36839 1639 36845
rect 1581 36805 1593 36839
rect 1627 36836 1639 36839
rect 3421 36839 3479 36845
rect 1627 36808 2774 36836
rect 1627 36805 1639 36808
rect 1581 36799 1639 36805
rect 2131 36771 2189 36777
rect 2131 36737 2143 36771
rect 2177 36768 2189 36771
rect 2498 36768 2504 36780
rect 2177 36740 2504 36768
rect 2177 36737 2189 36740
rect 2131 36731 2189 36737
rect 2498 36728 2504 36740
rect 2556 36728 2562 36780
rect 2746 36768 2774 36808
rect 3421 36805 3433 36839
rect 3467 36836 3479 36839
rect 3510 36836 3516 36848
rect 3467 36808 3516 36836
rect 3467 36805 3479 36808
rect 3421 36799 3479 36805
rect 3510 36796 3516 36808
rect 3568 36796 3574 36848
rect 3602 36796 3608 36848
rect 3660 36836 3666 36848
rect 3804 36845 3832 36876
rect 5905 36873 5917 36876
rect 5951 36873 5963 36907
rect 5905 36867 5963 36873
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 8018 36904 8024 36916
rect 7055 36876 8024 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 8018 36864 8024 36876
rect 8076 36864 8082 36916
rect 8202 36864 8208 36916
rect 8260 36904 8266 36916
rect 8478 36904 8484 36916
rect 8260 36876 8484 36904
rect 8260 36864 8266 36876
rect 8478 36864 8484 36876
rect 8536 36864 8542 36916
rect 17218 36904 17224 36916
rect 12406 36876 17224 36904
rect 3697 36839 3755 36845
rect 3697 36836 3709 36839
rect 3660 36808 3709 36836
rect 3660 36796 3666 36808
rect 3697 36805 3709 36808
rect 3743 36805 3755 36839
rect 3697 36799 3755 36805
rect 3789 36839 3847 36845
rect 3789 36805 3801 36839
rect 3835 36805 3847 36839
rect 7466 36836 7472 36848
rect 3789 36799 3847 36805
rect 3896 36808 7472 36836
rect 3896 36768 3924 36808
rect 7466 36796 7472 36808
rect 7524 36796 7530 36848
rect 9766 36836 9772 36848
rect 9140 36808 9772 36836
rect 9140 36780 9168 36808
rect 9766 36796 9772 36808
rect 9824 36796 9830 36848
rect 2746 36740 3924 36768
rect 4157 36771 4215 36777
rect 4157 36737 4169 36771
rect 4203 36768 4215 36771
rect 4338 36768 4344 36780
rect 4203 36740 4344 36768
rect 4203 36737 4215 36740
rect 4157 36731 4215 36737
rect 4338 36728 4344 36740
rect 4396 36728 4402 36780
rect 4539 36771 4597 36777
rect 4539 36737 4551 36771
rect 4585 36737 4597 36771
rect 4539 36731 4597 36737
rect 1857 36703 1915 36709
rect 1857 36669 1869 36703
rect 1903 36669 1915 36703
rect 4554 36700 4582 36731
rect 4706 36728 4712 36780
rect 4764 36768 4770 36780
rect 5167 36771 5225 36777
rect 5167 36768 5179 36771
rect 4764 36740 5179 36768
rect 4764 36728 4770 36740
rect 5167 36737 5179 36740
rect 5213 36768 5225 36771
rect 5213 36740 5948 36768
rect 5213 36737 5225 36740
rect 5167 36731 5225 36737
rect 4798 36700 4804 36712
rect 1857 36663 1915 36669
rect 1762 36592 1768 36644
rect 1820 36592 1826 36644
rect 1872 36564 1900 36663
rect 2869 36635 2927 36641
rect 2869 36601 2881 36635
rect 2915 36632 2927 36635
rect 3252 36632 3280 36686
rect 4554 36672 4804 36700
rect 4798 36660 4804 36672
rect 4856 36660 4862 36712
rect 4893 36703 4951 36709
rect 4893 36669 4905 36703
rect 4939 36669 4951 36703
rect 5920 36700 5948 36740
rect 6914 36728 6920 36780
rect 6972 36728 6978 36780
rect 7006 36728 7012 36780
rect 7064 36728 7070 36780
rect 7098 36728 7104 36780
rect 7156 36768 7162 36780
rect 7377 36771 7435 36777
rect 7377 36768 7389 36771
rect 7156 36740 7389 36768
rect 7156 36728 7162 36740
rect 7377 36737 7389 36740
rect 7423 36737 7435 36771
rect 7742 36768 7748 36780
rect 7703 36740 7748 36768
rect 7377 36731 7435 36737
rect 7742 36728 7748 36740
rect 7800 36768 7806 36780
rect 9122 36768 9128 36780
rect 7800 36740 9128 36768
rect 7800 36728 7806 36740
rect 9122 36728 9128 36740
rect 9180 36728 9186 36780
rect 9306 36728 9312 36780
rect 9364 36768 9370 36780
rect 11759 36771 11817 36777
rect 11759 36768 11771 36771
rect 9364 36740 11771 36768
rect 9364 36728 9370 36740
rect 11759 36737 11771 36740
rect 11805 36768 11817 36771
rect 12406 36768 12434 36876
rect 17218 36864 17224 36876
rect 17276 36864 17282 36916
rect 19613 36907 19671 36913
rect 19613 36873 19625 36907
rect 19659 36904 19671 36907
rect 20349 36907 20407 36913
rect 19659 36876 20300 36904
rect 19659 36873 19671 36876
rect 19613 36867 19671 36873
rect 14366 36796 14372 36848
rect 14424 36836 14430 36848
rect 19334 36836 19340 36848
rect 14424 36808 19340 36836
rect 14424 36796 14430 36808
rect 19334 36796 19340 36808
rect 19392 36796 19398 36848
rect 20272 36836 20300 36876
rect 20349 36873 20361 36907
rect 20395 36904 20407 36907
rect 20714 36904 20720 36916
rect 20395 36876 20720 36904
rect 20395 36873 20407 36876
rect 20349 36867 20407 36873
rect 20714 36864 20720 36876
rect 20772 36864 20778 36916
rect 20901 36907 20959 36913
rect 20901 36873 20913 36907
rect 20947 36904 20959 36907
rect 21818 36904 21824 36916
rect 20947 36876 21824 36904
rect 20947 36873 20959 36876
rect 20901 36867 20959 36873
rect 21818 36864 21824 36876
rect 21876 36864 21882 36916
rect 23842 36904 23848 36916
rect 22066 36876 23848 36904
rect 20272 36808 20852 36836
rect 11805 36740 12434 36768
rect 11805 36737 11817 36740
rect 11759 36731 11817 36737
rect 16666 36728 16672 36780
rect 16724 36728 16730 36780
rect 17773 36771 17831 36777
rect 17773 36737 17785 36771
rect 17819 36737 17831 36771
rect 19153 36771 19211 36777
rect 19153 36768 19165 36771
rect 17773 36731 17831 36737
rect 18248 36740 19165 36768
rect 7024 36700 7052 36728
rect 7466 36700 7472 36712
rect 5920 36672 7052 36700
rect 7114 36672 7472 36700
rect 4893 36663 4951 36669
rect 4908 36632 4936 36663
rect 2915 36604 3280 36632
rect 4632 36604 4936 36632
rect 2915 36601 2927 36604
rect 2869 36595 2927 36601
rect 4632 36576 4660 36604
rect 2314 36564 2320 36576
rect 1872 36536 2320 36564
rect 2314 36524 2320 36536
rect 2372 36524 2378 36576
rect 4614 36524 4620 36576
rect 4672 36524 4678 36576
rect 4709 36567 4767 36573
rect 4709 36533 4721 36567
rect 4755 36564 4767 36567
rect 4798 36564 4804 36576
rect 4755 36536 4804 36564
rect 4755 36533 4767 36536
rect 4709 36527 4767 36533
rect 4798 36524 4804 36536
rect 4856 36524 4862 36576
rect 4908 36564 4936 36604
rect 7114 36564 7142 36672
rect 7466 36660 7472 36672
rect 7524 36660 7530 36712
rect 8202 36660 8208 36712
rect 8260 36660 8266 36712
rect 10042 36660 10048 36712
rect 10100 36700 10106 36712
rect 10778 36700 10784 36712
rect 10100 36672 10784 36700
rect 10100 36660 10106 36672
rect 10778 36660 10784 36672
rect 10836 36700 10842 36712
rect 11517 36703 11575 36709
rect 11517 36700 11529 36703
rect 10836 36672 11529 36700
rect 10836 36660 10842 36672
rect 11517 36669 11529 36672
rect 11563 36669 11575 36703
rect 11517 36663 11575 36669
rect 4908 36536 7142 36564
rect 7193 36567 7251 36573
rect 7193 36533 7205 36567
rect 7239 36564 7251 36567
rect 8220 36564 8248 36660
rect 7239 36536 8248 36564
rect 7239 36533 7251 36536
rect 7193 36527 7251 36533
rect 8386 36524 8392 36576
rect 8444 36564 8450 36576
rect 8481 36567 8539 36573
rect 8481 36564 8493 36567
rect 8444 36536 8493 36564
rect 8444 36524 8450 36536
rect 8481 36533 8493 36536
rect 8527 36533 8539 36567
rect 8481 36527 8539 36533
rect 8938 36524 8944 36576
rect 8996 36564 9002 36576
rect 10502 36564 10508 36576
rect 8996 36536 10508 36564
rect 8996 36524 9002 36536
rect 10502 36524 10508 36536
rect 10560 36524 10566 36576
rect 11532 36564 11560 36663
rect 16684 36632 16712 36728
rect 17402 36660 17408 36712
rect 17460 36700 17466 36712
rect 17788 36700 17816 36731
rect 17460 36672 17816 36700
rect 17460 36660 17466 36672
rect 18248 36644 18276 36740
rect 19153 36737 19165 36740
rect 19199 36737 19211 36771
rect 19153 36731 19211 36737
rect 19797 36775 19855 36781
rect 19797 36741 19809 36775
rect 19843 36741 19855 36775
rect 20257 36771 20315 36777
rect 20257 36768 20269 36771
rect 19797 36735 19855 36741
rect 19904 36740 20269 36768
rect 19812 36700 19840 36735
rect 18984 36672 19840 36700
rect 12174 36604 16712 36632
rect 12174 36564 12202 36604
rect 17310 36592 17316 36644
rect 17368 36592 17374 36644
rect 17492 36604 18092 36632
rect 11532 36536 12202 36564
rect 12526 36524 12532 36576
rect 12584 36524 12590 36576
rect 17328 36564 17356 36592
rect 17492 36564 17520 36604
rect 17328 36536 17520 36564
rect 17589 36567 17647 36573
rect 17589 36533 17601 36567
rect 17635 36564 17647 36567
rect 17954 36564 17960 36576
rect 17635 36536 17960 36564
rect 17635 36533 17647 36536
rect 17589 36527 17647 36533
rect 17954 36524 17960 36536
rect 18012 36524 18018 36576
rect 18064 36564 18092 36604
rect 18230 36592 18236 36644
rect 18288 36592 18294 36644
rect 18984 36641 19012 36672
rect 18969 36635 19027 36641
rect 18969 36601 18981 36635
rect 19015 36601 19027 36635
rect 18969 36595 19027 36601
rect 19334 36592 19340 36644
rect 19392 36632 19398 36644
rect 19702 36632 19708 36644
rect 19392 36604 19708 36632
rect 19392 36592 19398 36604
rect 19702 36592 19708 36604
rect 19760 36632 19766 36644
rect 19904 36632 19932 36740
rect 20257 36737 20269 36740
rect 20303 36737 20315 36771
rect 20257 36731 20315 36737
rect 20530 36728 20536 36780
rect 20588 36728 20594 36780
rect 20824 36777 20852 36808
rect 20809 36771 20867 36777
rect 20809 36737 20821 36771
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36737 21143 36771
rect 21085 36731 21143 36737
rect 21100 36700 21128 36731
rect 20364 36672 21128 36700
rect 19760 36604 19932 36632
rect 20073 36635 20131 36641
rect 19760 36592 19766 36604
rect 20073 36601 20085 36635
rect 20119 36632 20131 36635
rect 20364 36632 20392 36672
rect 22066 36632 22094 36876
rect 23842 36864 23848 36876
rect 23900 36864 23906 36916
rect 23937 36907 23995 36913
rect 23937 36873 23949 36907
rect 23983 36904 23995 36907
rect 24026 36904 24032 36916
rect 23983 36876 24032 36904
rect 23983 36873 23995 36876
rect 23937 36867 23995 36873
rect 24026 36864 24032 36876
rect 24084 36864 24090 36916
rect 23661 36839 23719 36845
rect 23661 36805 23673 36839
rect 23707 36836 23719 36839
rect 23707 36808 25636 36836
rect 23707 36805 23719 36808
rect 23661 36799 23719 36805
rect 23014 36728 23020 36780
rect 23072 36728 23078 36780
rect 23293 36771 23351 36777
rect 23293 36737 23305 36771
rect 23339 36768 23351 36771
rect 24026 36768 24032 36780
rect 23339 36740 24032 36768
rect 23339 36737 23351 36740
rect 23293 36731 23351 36737
rect 24026 36728 24032 36740
rect 24084 36728 24090 36780
rect 24136 36777 24164 36808
rect 25608 36780 25636 36808
rect 24121 36771 24179 36777
rect 24121 36737 24133 36771
rect 24167 36737 24179 36771
rect 24121 36731 24179 36737
rect 24213 36771 24271 36777
rect 24213 36737 24225 36771
rect 24259 36737 24271 36771
rect 24213 36731 24271 36737
rect 22370 36660 22376 36712
rect 22428 36700 22434 36712
rect 24228 36700 24256 36731
rect 25590 36728 25596 36780
rect 25648 36728 25654 36780
rect 22428 36672 24256 36700
rect 22428 36660 22434 36672
rect 20119 36604 20392 36632
rect 20640 36604 22094 36632
rect 23109 36635 23167 36641
rect 20119 36601 20131 36604
rect 20073 36595 20131 36601
rect 20530 36564 20536 36576
rect 18064 36536 20536 36564
rect 20530 36524 20536 36536
rect 20588 36524 20594 36576
rect 20640 36573 20668 36604
rect 23109 36601 23121 36635
rect 23155 36632 23167 36635
rect 24210 36632 24216 36644
rect 23155 36604 24216 36632
rect 23155 36601 23167 36604
rect 23109 36595 23167 36601
rect 24210 36592 24216 36604
rect 24268 36592 24274 36644
rect 20625 36567 20683 36573
rect 20625 36533 20637 36567
rect 20671 36533 20683 36567
rect 20625 36527 20683 36533
rect 22830 36524 22836 36576
rect 22888 36524 22894 36576
rect 24394 36524 24400 36576
rect 24452 36524 24458 36576
rect 1104 36474 24840 36496
rect 1104 36422 3917 36474
rect 3969 36422 3981 36474
rect 4033 36422 4045 36474
rect 4097 36422 4109 36474
rect 4161 36422 4173 36474
rect 4225 36422 9851 36474
rect 9903 36422 9915 36474
rect 9967 36422 9979 36474
rect 10031 36422 10043 36474
rect 10095 36422 10107 36474
rect 10159 36422 15785 36474
rect 15837 36422 15849 36474
rect 15901 36422 15913 36474
rect 15965 36422 15977 36474
rect 16029 36422 16041 36474
rect 16093 36422 21719 36474
rect 21771 36422 21783 36474
rect 21835 36422 21847 36474
rect 21899 36422 21911 36474
rect 21963 36422 21975 36474
rect 22027 36422 24840 36474
rect 1104 36400 24840 36422
rect 1762 36320 1768 36372
rect 1820 36360 1826 36372
rect 2498 36360 2504 36372
rect 1820 36332 2504 36360
rect 1820 36320 1826 36332
rect 2498 36320 2504 36332
rect 2556 36360 2562 36372
rect 4709 36363 4767 36369
rect 4709 36360 4721 36363
rect 2556 36332 4721 36360
rect 2556 36320 2562 36332
rect 4709 36329 4721 36332
rect 4755 36360 4767 36363
rect 4755 36332 6682 36360
rect 4755 36329 4767 36332
rect 4709 36323 4767 36329
rect 3142 36252 3148 36304
rect 3200 36292 3206 36304
rect 3418 36292 3424 36304
rect 3200 36264 3424 36292
rect 3200 36252 3206 36264
rect 3418 36252 3424 36264
rect 3476 36252 3482 36304
rect 3786 36252 3792 36304
rect 3844 36292 3850 36304
rect 4614 36292 4620 36304
rect 3844 36264 4620 36292
rect 3844 36252 3850 36264
rect 4614 36252 4620 36264
rect 4672 36252 4678 36304
rect 4798 36252 4804 36304
rect 4856 36292 4862 36304
rect 4856 36264 5304 36292
rect 4856 36252 4862 36264
rect 2792 36196 3280 36224
rect 1489 36159 1547 36165
rect 1489 36125 1501 36159
rect 1535 36156 1547 36159
rect 1670 36156 1676 36168
rect 1535 36128 1676 36156
rect 1535 36125 1547 36128
rect 1489 36119 1547 36125
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 1763 36159 1821 36165
rect 1763 36125 1775 36159
rect 1809 36156 1821 36159
rect 2792 36156 2820 36196
rect 1809 36128 2820 36156
rect 1809 36125 1821 36128
rect 1763 36119 1821 36125
rect 2866 36116 2872 36168
rect 2924 36116 2930 36168
rect 3145 36091 3203 36097
rect 3145 36088 3157 36091
rect 2056 36060 3157 36088
rect 2056 36032 2084 36060
rect 3145 36057 3157 36060
rect 3191 36057 3203 36091
rect 3145 36051 3203 36057
rect 2038 35980 2044 36032
rect 2096 35980 2102 36032
rect 2501 36023 2559 36029
rect 2501 35989 2513 36023
rect 2547 36020 2559 36023
rect 2682 36020 2688 36032
rect 2547 35992 2688 36020
rect 2547 35989 2559 35992
rect 2501 35983 2559 35989
rect 2682 35980 2688 35992
rect 2740 35980 2746 36032
rect 3050 35980 3056 36032
rect 3108 36020 3114 36032
rect 3252 36020 3280 36196
rect 4338 36184 4344 36236
rect 4396 36224 4402 36236
rect 4522 36224 4528 36236
rect 4396 36196 4528 36224
rect 4396 36184 4402 36196
rect 4522 36184 4528 36196
rect 4580 36224 4586 36236
rect 4706 36224 4712 36236
rect 4580 36196 4712 36224
rect 4580 36184 4586 36196
rect 4706 36184 4712 36196
rect 4764 36184 4770 36236
rect 3786 36116 3792 36168
rect 3844 36116 3850 36168
rect 4798 36116 4804 36168
rect 4856 36156 4862 36168
rect 5074 36156 5080 36168
rect 4856 36128 5080 36156
rect 4856 36116 4862 36128
rect 5074 36116 5080 36128
rect 5132 36116 5138 36168
rect 5276 36165 5304 36264
rect 5442 36252 5448 36304
rect 5500 36292 5506 36304
rect 5721 36295 5779 36301
rect 5721 36292 5733 36295
rect 5500 36264 5733 36292
rect 5500 36252 5506 36264
rect 5721 36261 5733 36264
rect 5767 36261 5779 36295
rect 6654 36292 6682 36332
rect 6914 36320 6920 36372
rect 6972 36360 6978 36372
rect 7009 36363 7067 36369
rect 7009 36360 7021 36363
rect 6972 36332 7021 36360
rect 6972 36320 6978 36332
rect 7009 36329 7021 36332
rect 7055 36329 7067 36363
rect 7009 36323 7067 36329
rect 7834 36320 7840 36372
rect 7892 36360 7898 36372
rect 8018 36360 8024 36372
rect 7892 36332 8024 36360
rect 7892 36320 7898 36332
rect 8018 36320 8024 36332
rect 8076 36360 8082 36372
rect 22094 36360 22100 36372
rect 8076 36332 22100 36360
rect 8076 36320 8082 36332
rect 22094 36320 22100 36332
rect 22152 36320 22158 36372
rect 22370 36320 22376 36372
rect 22428 36320 22434 36372
rect 22830 36320 22836 36372
rect 22888 36320 22894 36372
rect 23385 36363 23443 36369
rect 23385 36329 23397 36363
rect 23431 36360 23443 36363
rect 23566 36360 23572 36372
rect 23431 36332 23572 36360
rect 23431 36329 23443 36332
rect 23385 36323 23443 36329
rect 23566 36320 23572 36332
rect 23624 36320 23630 36372
rect 10965 36295 11023 36301
rect 6654 36264 7328 36292
rect 5721 36255 5779 36261
rect 5350 36184 5356 36236
rect 5408 36224 5414 36236
rect 6135 36227 6193 36233
rect 6135 36224 6147 36227
rect 5408 36196 6147 36224
rect 5408 36184 5414 36196
rect 6135 36193 6147 36196
rect 6181 36193 6193 36227
rect 6135 36187 6193 36193
rect 6273 36227 6331 36233
rect 6273 36193 6285 36227
rect 6319 36224 6331 36227
rect 6454 36224 6460 36236
rect 6319 36196 6460 36224
rect 6319 36193 6331 36196
rect 6273 36187 6331 36193
rect 6454 36184 6460 36196
rect 6512 36184 6518 36236
rect 6638 36184 6644 36236
rect 6696 36224 6702 36236
rect 6696 36196 7236 36224
rect 6696 36184 6702 36196
rect 5261 36159 5319 36165
rect 5261 36125 5273 36159
rect 5307 36125 5319 36159
rect 5261 36119 5319 36125
rect 4062 36048 4068 36100
rect 4120 36048 4126 36100
rect 4433 36091 4491 36097
rect 4433 36057 4445 36091
rect 4479 36057 4491 36091
rect 4433 36051 4491 36057
rect 3108 35992 3280 36020
rect 3108 35980 3114 35992
rect 3602 35980 3608 36032
rect 3660 36020 3666 36032
rect 4448 36020 4476 36051
rect 3660 35992 4476 36020
rect 3660 35980 3666 35992
rect 4890 35980 4896 36032
rect 4948 36020 4954 36032
rect 5074 36020 5080 36032
rect 4948 35992 5080 36020
rect 4948 35980 4954 35992
rect 5074 35980 5080 35992
rect 5132 35980 5138 36032
rect 5276 36020 5304 36119
rect 5994 36116 6000 36168
rect 6052 36116 6058 36168
rect 6917 36159 6975 36165
rect 6917 36125 6929 36159
rect 6963 36156 6975 36159
rect 7098 36156 7104 36168
rect 6963 36128 7104 36156
rect 6963 36125 6975 36128
rect 6917 36119 6975 36125
rect 7098 36116 7104 36128
rect 7156 36116 7162 36168
rect 7208 36165 7236 36196
rect 7193 36159 7251 36165
rect 7193 36125 7205 36159
rect 7239 36125 7251 36159
rect 7193 36119 7251 36125
rect 7300 36088 7328 36264
rect 10965 36261 10977 36295
rect 11011 36292 11023 36295
rect 11054 36292 11060 36304
rect 11011 36264 11060 36292
rect 11011 36261 11023 36264
rect 10965 36255 11023 36261
rect 11054 36252 11060 36264
rect 11112 36252 11118 36304
rect 12526 36292 12532 36304
rect 12406 36264 12532 36292
rect 7466 36184 7472 36236
rect 7524 36224 7530 36236
rect 8938 36224 8944 36236
rect 7524 36196 8944 36224
rect 7524 36184 7530 36196
rect 8938 36184 8944 36196
rect 8996 36184 9002 36236
rect 9858 36184 9864 36236
rect 9916 36224 9922 36236
rect 10594 36224 10600 36236
rect 9916 36196 10600 36224
rect 9916 36184 9922 36196
rect 10594 36184 10600 36196
rect 10652 36224 10658 36236
rect 11517 36227 11575 36233
rect 10652 36196 11284 36224
rect 10652 36184 10658 36196
rect 11256 36168 11284 36196
rect 11517 36193 11529 36227
rect 11563 36224 11575 36227
rect 12406 36224 12434 36264
rect 12526 36252 12532 36264
rect 12584 36252 12590 36304
rect 22848 36224 22876 36320
rect 11563 36196 12434 36224
rect 18708 36196 19288 36224
rect 22848 36196 23888 36224
rect 11563 36193 11575 36196
rect 11517 36187 11575 36193
rect 7374 36116 7380 36168
rect 7432 36156 7438 36168
rect 8662 36156 8668 36168
rect 7432 36128 8668 36156
rect 7432 36116 7438 36128
rect 8662 36116 8668 36128
rect 8720 36156 8726 36168
rect 9183 36159 9241 36165
rect 9183 36156 9195 36159
rect 8720 36128 9195 36156
rect 8720 36116 8726 36128
rect 9183 36125 9195 36128
rect 9229 36156 9241 36159
rect 9306 36156 9312 36168
rect 9229 36128 9312 36156
rect 9229 36125 9241 36128
rect 9183 36119 9241 36125
rect 9306 36116 9312 36128
rect 9364 36116 9370 36168
rect 9674 36116 9680 36168
rect 9732 36156 9738 36168
rect 10321 36159 10379 36165
rect 10321 36156 10333 36159
rect 9732 36128 10333 36156
rect 9732 36116 9738 36128
rect 10321 36125 10333 36128
rect 10367 36125 10379 36159
rect 10321 36119 10379 36125
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36125 10563 36159
rect 10505 36119 10563 36125
rect 7300 36060 10102 36088
rect 5534 36020 5540 36032
rect 5276 35992 5540 36020
rect 5534 35980 5540 35992
rect 5592 35980 5598 36032
rect 7006 35980 7012 36032
rect 7064 36020 7070 36032
rect 7374 36020 7380 36032
rect 7064 35992 7380 36020
rect 7064 35980 7070 35992
rect 7374 35980 7380 35992
rect 7432 35980 7438 36032
rect 7742 35980 7748 36032
rect 7800 36020 7806 36032
rect 9858 36020 9864 36032
rect 7800 35992 9864 36020
rect 7800 35980 7806 35992
rect 9858 35980 9864 35992
rect 9916 35980 9922 36032
rect 9950 35980 9956 36032
rect 10008 35980 10014 36032
rect 10074 36020 10102 36060
rect 10134 36048 10140 36100
rect 10192 36088 10198 36100
rect 10520 36088 10548 36119
rect 11238 36116 11244 36168
rect 11296 36116 11302 36168
rect 11422 36165 11428 36168
rect 11379 36159 11428 36165
rect 11379 36125 11391 36159
rect 11425 36125 11428 36159
rect 11379 36119 11428 36125
rect 11422 36116 11428 36119
rect 11480 36116 11486 36168
rect 17129 36159 17187 36165
rect 17129 36125 17141 36159
rect 17175 36156 17187 36159
rect 18708 36156 18736 36196
rect 19260 36168 19288 36196
rect 17175 36128 18736 36156
rect 18785 36159 18843 36165
rect 17175 36125 17187 36128
rect 17129 36119 17187 36125
rect 18785 36125 18797 36159
rect 18831 36125 18843 36159
rect 18785 36119 18843 36125
rect 17402 36097 17408 36100
rect 10192 36060 10548 36088
rect 12161 36091 12219 36097
rect 10192 36048 10198 36060
rect 12161 36057 12173 36091
rect 12207 36088 12219 36091
rect 17374 36091 17408 36097
rect 17374 36088 17386 36091
rect 12207 36060 17386 36088
rect 12207 36057 12219 36060
rect 12161 36051 12219 36057
rect 17374 36057 17386 36060
rect 17374 36051 17408 36057
rect 17402 36048 17408 36051
rect 17460 36048 17466 36100
rect 18800 36088 18828 36119
rect 19242 36116 19248 36168
rect 19300 36116 19306 36168
rect 20254 36116 20260 36168
rect 20312 36156 20318 36168
rect 21177 36159 21235 36165
rect 21177 36156 21189 36159
rect 20312 36128 21189 36156
rect 20312 36116 20318 36128
rect 21177 36125 21189 36128
rect 21223 36125 21235 36159
rect 21177 36119 21235 36125
rect 21821 36159 21879 36165
rect 21821 36125 21833 36159
rect 21867 36125 21879 36159
rect 22557 36159 22615 36165
rect 22557 36156 22569 36159
rect 21821 36119 21879 36125
rect 22066 36128 22569 36156
rect 21836 36088 21864 36119
rect 18524 36060 18828 36088
rect 21008 36060 21864 36088
rect 14274 36020 14280 36032
rect 10074 35992 14280 36020
rect 14274 35980 14280 35992
rect 14332 35980 14338 36032
rect 18524 36029 18552 36060
rect 18509 36023 18567 36029
rect 18509 35989 18521 36023
rect 18555 35989 18567 36023
rect 18509 35983 18567 35989
rect 18601 36023 18659 36029
rect 18601 35989 18613 36023
rect 18647 36020 18659 36023
rect 19334 36020 19340 36032
rect 18647 35992 19340 36020
rect 18647 35989 18659 35992
rect 18601 35983 18659 35989
rect 19334 35980 19340 35992
rect 19392 35980 19398 36032
rect 21008 36029 21036 36060
rect 20993 36023 21051 36029
rect 20993 35989 21005 36023
rect 21039 35989 21051 36023
rect 20993 35983 21051 35989
rect 21637 36023 21695 36029
rect 21637 35989 21649 36023
rect 21683 36020 21695 36023
rect 22066 36020 22094 36128
rect 22557 36125 22569 36128
rect 22603 36125 22615 36159
rect 22557 36119 22615 36125
rect 23566 36116 23572 36168
rect 23624 36116 23630 36168
rect 23860 36165 23888 36196
rect 23845 36159 23903 36165
rect 23845 36125 23857 36159
rect 23891 36125 23903 36159
rect 23845 36119 23903 36125
rect 24213 36091 24271 36097
rect 24213 36057 24225 36091
rect 24259 36088 24271 36091
rect 25130 36088 25136 36100
rect 24259 36060 25136 36088
rect 24259 36057 24271 36060
rect 24213 36051 24271 36057
rect 25130 36048 25136 36060
rect 25188 36048 25194 36100
rect 21683 35992 22094 36020
rect 21683 35989 21695 35992
rect 21637 35983 21695 35989
rect 1104 35930 25000 35952
rect 1104 35878 6884 35930
rect 6936 35878 6948 35930
rect 7000 35878 7012 35930
rect 7064 35878 7076 35930
rect 7128 35878 7140 35930
rect 7192 35878 12818 35930
rect 12870 35878 12882 35930
rect 12934 35878 12946 35930
rect 12998 35878 13010 35930
rect 13062 35878 13074 35930
rect 13126 35878 18752 35930
rect 18804 35878 18816 35930
rect 18868 35878 18880 35930
rect 18932 35878 18944 35930
rect 18996 35878 19008 35930
rect 19060 35878 24686 35930
rect 24738 35878 24750 35930
rect 24802 35878 24814 35930
rect 24866 35878 24878 35930
rect 24930 35878 24942 35930
rect 24994 35878 25000 35930
rect 1104 35856 25000 35878
rect 1688 35788 3280 35816
rect 1688 35689 1716 35788
rect 3252 35748 3280 35788
rect 3326 35776 3332 35828
rect 3384 35776 3390 35828
rect 4522 35776 4528 35828
rect 4580 35816 4586 35828
rect 5258 35816 5264 35828
rect 4580 35788 5264 35816
rect 4580 35776 4586 35788
rect 5258 35776 5264 35788
rect 5316 35776 5322 35828
rect 6181 35819 6239 35825
rect 6181 35785 6193 35819
rect 6227 35816 6239 35819
rect 6638 35816 6644 35828
rect 6227 35788 6644 35816
rect 6227 35785 6239 35788
rect 6181 35779 6239 35785
rect 6638 35776 6644 35788
rect 6696 35776 6702 35828
rect 9950 35816 9956 35828
rect 8588 35788 9956 35816
rect 3252 35720 4568 35748
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35649 1731 35683
rect 1673 35643 1731 35649
rect 2682 35640 2688 35692
rect 2740 35640 2746 35692
rect 3418 35640 3424 35692
rect 3476 35640 3482 35692
rect 4540 35689 4568 35720
rect 8202 35708 8208 35760
rect 8260 35708 8266 35760
rect 8588 35757 8616 35788
rect 9950 35776 9956 35788
rect 10008 35776 10014 35828
rect 11698 35776 11704 35828
rect 11756 35776 11762 35828
rect 14185 35819 14243 35825
rect 14185 35816 14197 35819
rect 12084 35788 14197 35816
rect 8573 35751 8631 35757
rect 8573 35717 8585 35751
rect 8619 35717 8631 35751
rect 9214 35748 9220 35760
rect 8573 35711 8631 35717
rect 8680 35720 9220 35748
rect 4525 35683 4583 35689
rect 4525 35649 4537 35683
rect 4571 35649 4583 35683
rect 4525 35643 4583 35649
rect 8481 35683 8539 35689
rect 8481 35649 8493 35683
rect 8527 35680 8539 35683
rect 8680 35680 8708 35720
rect 9214 35708 9220 35720
rect 9272 35708 9278 35760
rect 9309 35751 9367 35757
rect 9309 35717 9321 35751
rect 9355 35748 9367 35751
rect 9355 35720 9628 35748
rect 9355 35717 9367 35720
rect 9309 35711 9367 35717
rect 9600 35692 9628 35720
rect 11238 35708 11244 35760
rect 11296 35748 11302 35760
rect 11422 35748 11428 35760
rect 11296 35720 11428 35748
rect 11296 35708 11302 35720
rect 11422 35708 11428 35720
rect 11480 35708 11486 35760
rect 11974 35708 11980 35760
rect 12032 35708 12038 35760
rect 12084 35757 12112 35788
rect 14185 35785 14197 35788
rect 14231 35785 14243 35819
rect 14185 35779 14243 35785
rect 15194 35776 15200 35828
rect 15252 35816 15258 35828
rect 18230 35816 18236 35828
rect 15252 35788 18236 35816
rect 15252 35776 15258 35788
rect 18230 35776 18236 35788
rect 18288 35776 18294 35828
rect 19334 35776 19340 35828
rect 19392 35776 19398 35828
rect 21821 35819 21879 35825
rect 21821 35785 21833 35819
rect 21867 35816 21879 35819
rect 21867 35788 22600 35816
rect 21867 35785 21879 35788
rect 21821 35779 21879 35785
rect 12069 35751 12127 35757
rect 12069 35717 12081 35751
rect 12115 35717 12127 35751
rect 12069 35711 12127 35717
rect 12342 35708 12348 35760
rect 12400 35748 12406 35760
rect 12400 35720 12572 35748
rect 12400 35708 12406 35720
rect 8527 35652 8708 35680
rect 8527 35649 8539 35652
rect 8481 35643 8539 35649
rect 1210 35572 1216 35624
rect 1268 35612 1274 35624
rect 1489 35615 1547 35621
rect 1489 35612 1501 35615
rect 1268 35584 1501 35612
rect 1268 35572 1274 35584
rect 1489 35581 1501 35584
rect 1535 35581 1547 35615
rect 2409 35615 2467 35621
rect 2409 35612 2421 35615
rect 1489 35575 1547 35581
rect 2240 35584 2421 35612
rect 2130 35504 2136 35556
rect 2188 35504 2194 35556
rect 1946 35436 1952 35488
rect 2004 35476 2010 35488
rect 2240 35476 2268 35584
rect 2409 35581 2421 35584
rect 2455 35581 2467 35615
rect 2409 35575 2467 35581
rect 2498 35572 2504 35624
rect 2556 35621 2562 35624
rect 2556 35615 2584 35621
rect 2572 35581 2584 35615
rect 2556 35575 2584 35581
rect 2556 35572 2562 35575
rect 3050 35572 3056 35624
rect 3108 35612 3114 35624
rect 3602 35612 3608 35624
rect 3108 35584 3608 35612
rect 3108 35572 3114 35584
rect 3602 35572 3608 35584
rect 3660 35572 3666 35624
rect 4341 35615 4399 35621
rect 4341 35581 4353 35615
rect 4387 35581 4399 35615
rect 4540 35612 4568 35643
rect 8754 35640 8760 35692
rect 8812 35680 8818 35692
rect 8941 35683 8999 35689
rect 8941 35680 8953 35683
rect 8812 35652 8953 35680
rect 8812 35640 8818 35652
rect 8941 35649 8953 35652
rect 8987 35649 8999 35683
rect 8941 35643 8999 35649
rect 9582 35640 9588 35692
rect 9640 35640 9646 35692
rect 9951 35683 10009 35689
rect 9951 35649 9963 35683
rect 9997 35680 10009 35683
rect 10410 35680 10416 35692
rect 9997 35652 10416 35680
rect 9997 35649 10009 35652
rect 9951 35643 10009 35649
rect 10410 35640 10416 35652
rect 10468 35640 10474 35692
rect 10962 35640 10968 35692
rect 11020 35680 11026 35692
rect 12437 35683 12495 35689
rect 12437 35680 12449 35683
rect 11020 35652 12449 35680
rect 11020 35640 11026 35652
rect 12437 35649 12449 35652
rect 12483 35649 12495 35683
rect 12544 35680 12572 35720
rect 12618 35708 12624 35760
rect 12676 35748 12682 35760
rect 12805 35751 12863 35757
rect 12805 35748 12817 35751
rect 12676 35720 12817 35748
rect 12676 35708 12682 35720
rect 12805 35717 12817 35720
rect 12851 35717 12863 35751
rect 12805 35711 12863 35717
rect 18414 35708 18420 35760
rect 18472 35748 18478 35760
rect 19245 35751 19303 35757
rect 19245 35748 19257 35751
rect 18472 35720 19257 35748
rect 18472 35708 18478 35720
rect 19245 35717 19257 35720
rect 19291 35717 19303 35751
rect 19352 35748 19380 35776
rect 19352 35720 19564 35748
rect 19245 35711 19303 35717
rect 13447 35683 13505 35689
rect 13447 35680 13459 35683
rect 12544 35652 13459 35680
rect 12437 35643 12495 35649
rect 13447 35649 13459 35652
rect 13493 35680 13505 35683
rect 13493 35652 15976 35680
rect 13493 35649 13505 35652
rect 13447 35643 13505 35649
rect 4614 35612 4620 35624
rect 4540 35584 4620 35612
rect 4341 35575 4399 35581
rect 4356 35544 4384 35575
rect 4614 35572 4620 35584
rect 4672 35572 4678 35624
rect 5258 35572 5264 35624
rect 5316 35572 5322 35624
rect 5350 35572 5356 35624
rect 5408 35621 5414 35624
rect 5408 35615 5436 35621
rect 5424 35581 5436 35615
rect 5408 35575 5436 35581
rect 5537 35615 5595 35621
rect 5537 35581 5549 35615
rect 5583 35612 5595 35615
rect 5583 35584 6408 35612
rect 5583 35581 5595 35584
rect 5537 35575 5595 35581
rect 5408 35572 5414 35575
rect 6380 35556 6408 35584
rect 8386 35572 8392 35624
rect 8444 35572 8450 35624
rect 9306 35572 9312 35624
rect 9364 35572 9370 35624
rect 9677 35615 9735 35621
rect 9677 35581 9689 35615
rect 9723 35581 9735 35615
rect 12802 35612 12808 35624
rect 12742 35584 12808 35612
rect 9677 35575 9735 35581
rect 4890 35544 4896 35556
rect 4356 35516 4896 35544
rect 4890 35504 4896 35516
rect 4948 35504 4954 35556
rect 4985 35547 5043 35553
rect 4985 35513 4997 35547
rect 5031 35513 5043 35547
rect 4985 35507 5043 35513
rect 2004 35448 2268 35476
rect 2004 35436 2010 35448
rect 2498 35436 2504 35488
rect 2556 35476 2562 35488
rect 4522 35476 4528 35488
rect 2556 35448 4528 35476
rect 2556 35436 2562 35448
rect 4522 35436 4528 35448
rect 4580 35436 4586 35488
rect 5000 35476 5028 35507
rect 6362 35504 6368 35556
rect 6420 35504 6426 35556
rect 9324 35544 9352 35572
rect 9493 35547 9551 35553
rect 9493 35544 9505 35547
rect 9324 35516 9505 35544
rect 9493 35513 9505 35516
rect 9539 35513 9551 35547
rect 9692 35544 9720 35575
rect 12802 35572 12808 35584
rect 12860 35572 12866 35624
rect 12894 35572 12900 35624
rect 12952 35612 12958 35624
rect 13173 35615 13231 35621
rect 13173 35612 13185 35615
rect 12952 35584 13185 35612
rect 12952 35572 12958 35584
rect 13173 35581 13185 35584
rect 13219 35581 13231 35615
rect 13173 35575 13231 35581
rect 9692 35516 9812 35544
rect 9493 35507 9551 35513
rect 9784 35488 9812 35516
rect 5442 35476 5448 35488
rect 5000 35448 5448 35476
rect 5442 35436 5448 35448
rect 5500 35436 5506 35488
rect 5994 35436 6000 35488
rect 6052 35476 6058 35488
rect 6454 35476 6460 35488
rect 6052 35448 6460 35476
rect 6052 35436 6058 35448
rect 6454 35436 6460 35448
rect 6512 35436 6518 35488
rect 7745 35479 7803 35485
rect 7745 35445 7757 35479
rect 7791 35476 7803 35479
rect 7834 35476 7840 35488
rect 7791 35448 7840 35476
rect 7791 35445 7803 35448
rect 7745 35439 7803 35445
rect 7834 35436 7840 35448
rect 7892 35436 7898 35488
rect 9766 35436 9772 35488
rect 9824 35436 9830 35488
rect 10594 35436 10600 35488
rect 10652 35476 10658 35488
rect 10689 35479 10747 35485
rect 10689 35476 10701 35479
rect 10652 35448 10701 35476
rect 10652 35436 10658 35448
rect 10689 35445 10701 35448
rect 10735 35445 10747 35479
rect 10689 35439 10747 35445
rect 12986 35436 12992 35488
rect 13044 35436 13050 35488
rect 15948 35476 15976 35652
rect 16758 35640 16764 35692
rect 16816 35680 16822 35692
rect 19536 35689 19564 35720
rect 22572 35689 22600 35788
rect 23014 35776 23020 35828
rect 23072 35816 23078 35828
rect 23109 35819 23167 35825
rect 23109 35816 23121 35819
rect 23072 35788 23121 35816
rect 23072 35776 23078 35788
rect 23109 35785 23121 35788
rect 23155 35785 23167 35819
rect 23109 35779 23167 35785
rect 23477 35819 23535 35825
rect 23477 35785 23489 35819
rect 23523 35816 23535 35819
rect 23566 35816 23572 35828
rect 23523 35788 23572 35816
rect 23523 35785 23535 35788
rect 23477 35779 23535 35785
rect 23566 35776 23572 35788
rect 23624 35776 23630 35828
rect 25130 35748 25136 35760
rect 23676 35720 25136 35748
rect 17831 35683 17889 35689
rect 17831 35680 17843 35683
rect 16816 35652 17843 35680
rect 16816 35640 16822 35652
rect 17831 35649 17843 35652
rect 17877 35649 17889 35683
rect 18969 35683 19027 35689
rect 18969 35680 18981 35683
rect 17831 35643 17889 35649
rect 18616 35652 18981 35680
rect 17586 35572 17592 35624
rect 17644 35572 17650 35624
rect 18616 35553 18644 35652
rect 18969 35649 18981 35652
rect 19015 35680 19027 35683
rect 19337 35683 19395 35689
rect 19337 35680 19349 35683
rect 19015 35652 19349 35680
rect 19015 35649 19027 35652
rect 18969 35643 19027 35649
rect 19337 35649 19349 35652
rect 19383 35649 19395 35683
rect 19337 35643 19395 35649
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 21269 35683 21327 35689
rect 21269 35680 21281 35683
rect 19521 35643 19579 35649
rect 19628 35652 21281 35680
rect 19058 35572 19064 35624
rect 19116 35572 19122 35624
rect 19245 35615 19303 35621
rect 19245 35581 19257 35615
rect 19291 35612 19303 35615
rect 19429 35615 19487 35621
rect 19429 35612 19441 35615
rect 19291 35584 19441 35612
rect 19291 35581 19303 35584
rect 19245 35575 19303 35581
rect 19429 35581 19441 35584
rect 19475 35581 19487 35615
rect 19429 35575 19487 35581
rect 18601 35547 18659 35553
rect 18601 35513 18613 35547
rect 18647 35513 18659 35547
rect 18601 35507 18659 35513
rect 18874 35504 18880 35556
rect 18932 35544 18938 35556
rect 19628 35544 19656 35652
rect 21269 35649 21281 35652
rect 21315 35649 21327 35683
rect 21269 35643 21327 35649
rect 22005 35683 22063 35689
rect 22005 35649 22017 35683
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 22557 35683 22615 35689
rect 22557 35649 22569 35683
rect 22603 35649 22615 35683
rect 22833 35683 22891 35689
rect 22833 35680 22845 35683
rect 22557 35643 22615 35649
rect 22664 35652 22845 35680
rect 22020 35612 22048 35643
rect 22664 35612 22692 35652
rect 22833 35649 22845 35652
rect 22879 35680 22891 35683
rect 23198 35680 23204 35692
rect 22879 35652 23204 35680
rect 22879 35649 22891 35652
rect 22833 35643 22891 35649
rect 23198 35640 23204 35652
rect 23256 35640 23262 35692
rect 23676 35689 23704 35720
rect 25130 35708 25136 35720
rect 25188 35708 25194 35760
rect 23293 35683 23351 35689
rect 23293 35649 23305 35683
rect 23339 35649 23351 35683
rect 23293 35643 23351 35649
rect 23661 35683 23719 35689
rect 23661 35649 23673 35683
rect 23707 35649 23719 35683
rect 23661 35643 23719 35649
rect 21100 35584 22048 35612
rect 22296 35584 22692 35612
rect 21100 35553 21128 35584
rect 18932 35516 19656 35544
rect 21085 35547 21143 35553
rect 18932 35504 18938 35516
rect 21085 35513 21097 35547
rect 21131 35513 21143 35547
rect 21085 35507 21143 35513
rect 22296 35476 22324 35584
rect 22649 35547 22707 35553
rect 22649 35513 22661 35547
rect 22695 35544 22707 35547
rect 23308 35544 23336 35643
rect 23934 35640 23940 35692
rect 23992 35640 23998 35692
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 24121 35643 24179 35649
rect 24136 35612 24164 35643
rect 22695 35516 23336 35544
rect 23676 35584 24164 35612
rect 22695 35513 22707 35516
rect 22649 35507 22707 35513
rect 15948 35448 22324 35476
rect 22373 35479 22431 35485
rect 22373 35445 22385 35479
rect 22419 35476 22431 35479
rect 23676 35476 23704 35584
rect 22419 35448 23704 35476
rect 22419 35445 22431 35448
rect 22373 35439 22431 35445
rect 23750 35436 23756 35488
rect 23808 35436 23814 35488
rect 24394 35436 24400 35488
rect 24452 35436 24458 35488
rect 1104 35386 24840 35408
rect 1104 35334 3917 35386
rect 3969 35334 3981 35386
rect 4033 35334 4045 35386
rect 4097 35334 4109 35386
rect 4161 35334 4173 35386
rect 4225 35334 9851 35386
rect 9903 35334 9915 35386
rect 9967 35334 9979 35386
rect 10031 35334 10043 35386
rect 10095 35334 10107 35386
rect 10159 35334 15785 35386
rect 15837 35334 15849 35386
rect 15901 35334 15913 35386
rect 15965 35334 15977 35386
rect 16029 35334 16041 35386
rect 16093 35334 21719 35386
rect 21771 35334 21783 35386
rect 21835 35334 21847 35386
rect 21899 35334 21911 35386
rect 21963 35334 21975 35386
rect 22027 35334 24840 35386
rect 1104 35312 24840 35334
rect 1946 35232 1952 35284
rect 2004 35272 2010 35284
rect 2004 35244 3280 35272
rect 2004 35232 2010 35244
rect 3252 35148 3280 35244
rect 5460 35244 6130 35272
rect 5460 35216 5488 35244
rect 3329 35207 3387 35213
rect 3329 35173 3341 35207
rect 3375 35173 3387 35207
rect 3329 35167 3387 35173
rect 2314 35096 2320 35148
rect 2372 35096 2378 35148
rect 3234 35096 3240 35148
rect 3292 35096 3298 35148
rect 3344 35136 3372 35167
rect 5442 35164 5448 35216
rect 5500 35164 5506 35216
rect 6102 35204 6130 35244
rect 6362 35232 6368 35284
rect 6420 35272 6426 35284
rect 6457 35275 6515 35281
rect 6457 35272 6469 35275
rect 6420 35244 6469 35272
rect 6420 35232 6426 35244
rect 6457 35241 6469 35244
rect 6503 35241 6515 35275
rect 7650 35272 7656 35284
rect 6457 35235 6515 35241
rect 6564 35244 7656 35272
rect 6564 35204 6592 35244
rect 7650 35232 7656 35244
rect 7708 35232 7714 35284
rect 7834 35232 7840 35284
rect 7892 35272 7898 35284
rect 9582 35272 9588 35284
rect 7892 35244 9588 35272
rect 7892 35232 7898 35244
rect 9582 35232 9588 35244
rect 9640 35232 9646 35284
rect 11606 35272 11612 35284
rect 9784 35244 11612 35272
rect 6102 35176 6592 35204
rect 7374 35164 7380 35216
rect 7432 35204 7438 35216
rect 9784 35204 9812 35244
rect 11606 35232 11612 35244
rect 11664 35232 11670 35284
rect 11790 35232 11796 35284
rect 11848 35272 11854 35284
rect 12066 35272 12072 35284
rect 11848 35244 12072 35272
rect 11848 35232 11854 35244
rect 12066 35232 12072 35244
rect 12124 35232 12130 35284
rect 12802 35232 12808 35284
rect 12860 35232 12866 35284
rect 13630 35232 13636 35284
rect 13688 35272 13694 35284
rect 18233 35275 18291 35281
rect 13688 35244 16344 35272
rect 13688 35232 13694 35244
rect 7432 35176 9812 35204
rect 7432 35164 7438 35176
rect 10410 35164 10416 35216
rect 10468 35164 10474 35216
rect 10505 35207 10563 35213
rect 10505 35173 10517 35207
rect 10551 35204 10563 35207
rect 10594 35204 10600 35216
rect 10551 35176 10600 35204
rect 10551 35173 10563 35176
rect 10505 35167 10563 35173
rect 10594 35164 10600 35176
rect 10652 35164 10658 35216
rect 16316 35204 16344 35244
rect 18233 35241 18245 35275
rect 18279 35272 18291 35275
rect 19058 35272 19064 35284
rect 18279 35244 19064 35272
rect 18279 35241 18291 35244
rect 18233 35235 18291 35241
rect 19058 35232 19064 35244
rect 19116 35232 19122 35284
rect 19306 35244 21128 35272
rect 19306 35204 19334 35244
rect 16316 35176 19334 35204
rect 19889 35207 19947 35213
rect 19889 35173 19901 35207
rect 19935 35173 19947 35207
rect 19889 35167 19947 35173
rect 5460 35136 5488 35164
rect 3344 35108 3818 35136
rect 5368 35108 5488 35136
rect 750 35028 756 35080
rect 808 35068 814 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 808 35040 1409 35068
rect 808 35028 814 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 2038 35028 2044 35080
rect 2096 35068 2102 35080
rect 2559 35071 2617 35077
rect 2559 35068 2571 35071
rect 2096 35040 2571 35068
rect 2096 35028 2102 35040
rect 2559 35037 2571 35040
rect 2605 35037 2617 35071
rect 2559 35031 2617 35037
rect 4246 35028 4252 35080
rect 4304 35028 4310 35080
rect 5368 35068 5396 35108
rect 6638 35096 6644 35148
rect 6696 35136 6702 35148
rect 10045 35139 10103 35145
rect 10045 35136 10057 35139
rect 6696 35108 10057 35136
rect 6696 35096 6702 35108
rect 10045 35105 10057 35108
rect 10091 35136 10103 35139
rect 10134 35136 10140 35148
rect 10091 35108 10140 35136
rect 10091 35105 10103 35108
rect 10045 35099 10103 35105
rect 10134 35096 10140 35108
rect 10192 35096 10198 35148
rect 10428 35136 10456 35164
rect 10781 35139 10839 35145
rect 10781 35136 10793 35139
rect 10244 35108 10793 35136
rect 4632 35040 5396 35068
rect 1673 35003 1731 35009
rect 1673 34969 1685 35003
rect 1719 35000 1731 35003
rect 1719 34972 4292 35000
rect 1719 34969 1731 34972
rect 1673 34963 1731 34969
rect 3510 34892 3516 34944
rect 3568 34932 3574 34944
rect 3973 34935 4031 34941
rect 3973 34932 3985 34935
rect 3568 34904 3985 34932
rect 3568 34892 3574 34904
rect 3973 34901 3985 34904
rect 4019 34901 4031 34935
rect 4264 34932 4292 34972
rect 4338 34960 4344 35012
rect 4396 34960 4402 35012
rect 4632 34932 4660 35040
rect 5442 35028 5448 35080
rect 5500 35028 5506 35080
rect 5626 35028 5632 35080
rect 5684 35068 5690 35080
rect 5719 35071 5777 35077
rect 5719 35068 5731 35071
rect 5684 35040 5731 35068
rect 5684 35028 5690 35040
rect 5719 35037 5731 35040
rect 5765 35037 5777 35071
rect 5719 35031 5777 35037
rect 8570 35028 8576 35080
rect 8628 35068 8634 35080
rect 9674 35068 9680 35080
rect 8628 35040 9680 35068
rect 8628 35028 8634 35040
rect 9674 35028 9680 35040
rect 9732 35068 9738 35080
rect 9861 35071 9919 35077
rect 9861 35068 9873 35071
rect 9732 35040 9873 35068
rect 9732 35028 9738 35040
rect 9861 35037 9873 35040
rect 9907 35037 9919 35071
rect 10244 35068 10272 35108
rect 10781 35105 10793 35108
rect 10827 35105 10839 35139
rect 10781 35099 10839 35105
rect 11238 35096 11244 35148
rect 11296 35136 11302 35148
rect 11793 35139 11851 35145
rect 11793 35136 11805 35139
rect 11296 35108 11805 35136
rect 11296 35096 11302 35108
rect 10962 35077 10968 35080
rect 9861 35031 9919 35037
rect 10074 35040 10272 35068
rect 10919 35071 10968 35077
rect 4706 34960 4712 35012
rect 4764 35000 4770 35012
rect 9950 35000 9956 35012
rect 4764 34972 9956 35000
rect 4764 34960 4770 34972
rect 9950 34960 9956 34972
rect 10008 34960 10014 35012
rect 4264 34904 4660 34932
rect 3973 34895 4031 34901
rect 5074 34892 5080 34944
rect 5132 34892 5138 34944
rect 5258 34892 5264 34944
rect 5316 34892 5322 34944
rect 5442 34892 5448 34944
rect 5500 34932 5506 34944
rect 5718 34932 5724 34944
rect 5500 34904 5724 34932
rect 5500 34892 5506 34904
rect 5718 34892 5724 34904
rect 5776 34892 5782 34944
rect 6730 34892 6736 34944
rect 6788 34932 6794 34944
rect 10074 34932 10102 35040
rect 10919 35037 10931 35071
rect 10965 35037 10968 35071
rect 10919 35031 10968 35037
rect 10934 35030 10968 35031
rect 10962 35028 10968 35030
rect 11020 35028 11026 35080
rect 11054 35028 11060 35080
rect 11112 35028 11118 35080
rect 6788 34904 10102 34932
rect 11624 34932 11652 35108
rect 11793 35105 11805 35108
rect 11839 35105 11851 35139
rect 11793 35099 11851 35105
rect 15286 35096 15292 35148
rect 15344 35136 15350 35148
rect 15657 35139 15715 35145
rect 15657 35136 15669 35139
rect 15344 35108 15669 35136
rect 15344 35096 15350 35108
rect 15657 35105 15669 35108
rect 15703 35105 15715 35139
rect 15657 35099 15715 35105
rect 16482 35096 16488 35148
rect 16540 35136 16546 35148
rect 18046 35136 18052 35148
rect 16540 35108 18052 35136
rect 16540 35096 16546 35108
rect 18046 35096 18052 35108
rect 18104 35096 18110 35148
rect 19904 35136 19932 35167
rect 21100 35136 21128 35244
rect 22462 35232 22468 35284
rect 22520 35272 22526 35284
rect 23201 35275 23259 35281
rect 23201 35272 23213 35275
rect 22520 35244 23213 35272
rect 22520 35232 22526 35244
rect 23201 35241 23213 35244
rect 23247 35241 23259 35275
rect 23201 35235 23259 35241
rect 23658 35232 23664 35284
rect 23716 35272 23722 35284
rect 24578 35272 24584 35284
rect 23716 35244 24584 35272
rect 23716 35232 23722 35244
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 19904 35108 21036 35136
rect 21100 35108 23704 35136
rect 11974 35028 11980 35080
rect 12032 35070 12038 35080
rect 12067 35071 12125 35077
rect 12067 35070 12079 35071
rect 12032 35042 12079 35070
rect 12032 35028 12038 35042
rect 12067 35037 12079 35042
rect 12113 35037 12125 35071
rect 12067 35031 12125 35037
rect 12894 35028 12900 35080
rect 12952 35068 12958 35080
rect 14093 35071 14151 35077
rect 14093 35068 14105 35071
rect 12952 35040 14105 35068
rect 12952 35028 12958 35040
rect 14093 35037 14105 35040
rect 14139 35037 14151 35071
rect 14093 35031 14151 35037
rect 14366 35028 14372 35080
rect 14424 35068 14430 35080
rect 15194 35068 15200 35080
rect 14424 35040 15200 35068
rect 14424 35028 14430 35040
rect 15194 35028 15200 35040
rect 15252 35028 15258 35080
rect 15931 35071 15989 35077
rect 15931 35037 15943 35071
rect 15977 35068 15989 35071
rect 16298 35068 16304 35080
rect 15977 35040 16304 35068
rect 15977 35037 15989 35040
rect 15931 35031 15989 35037
rect 16298 35028 16304 35040
rect 16356 35028 16362 35080
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 18141 35071 18199 35077
rect 18141 35068 18153 35071
rect 18012 35040 18153 35068
rect 18012 35028 18018 35040
rect 18141 35037 18153 35040
rect 18187 35037 18199 35071
rect 19334 35068 19340 35080
rect 18141 35031 18199 35037
rect 18246 35040 19340 35068
rect 11701 35003 11759 35009
rect 11701 34969 11713 35003
rect 11747 35000 11759 35003
rect 18246 35000 18274 35040
rect 19334 35028 19340 35040
rect 19392 35068 19398 35080
rect 21008 35077 21036 35108
rect 19705 35071 19763 35077
rect 19705 35068 19717 35071
rect 19392 35040 19717 35068
rect 19392 35028 19398 35040
rect 19705 35037 19717 35040
rect 19751 35037 19763 35071
rect 20993 35071 21051 35077
rect 19705 35031 19763 35037
rect 19810 35044 20024 35068
rect 20073 35047 20131 35053
rect 20073 35044 20085 35047
rect 19810 35040 20085 35044
rect 11747 34972 14136 35000
rect 11747 34969 11759 34972
rect 11701 34963 11759 34969
rect 12894 34932 12900 34944
rect 11624 34904 12900 34932
rect 6788 34892 6794 34904
rect 12894 34892 12900 34904
rect 12952 34892 12958 34944
rect 14108 34932 14136 34972
rect 14384 34972 18274 35000
rect 14384 34932 14412 34972
rect 19150 34960 19156 35012
rect 19208 35000 19214 35012
rect 19810 35000 19838 35040
rect 19996 35016 20085 35040
rect 20073 35013 20085 35016
rect 20119 35013 20131 35047
rect 20993 35037 21005 35071
rect 21039 35037 21051 35071
rect 20993 35031 21051 35037
rect 23382 35028 23388 35080
rect 23440 35028 23446 35080
rect 23676 35077 23704 35108
rect 23661 35071 23719 35077
rect 23661 35037 23673 35071
rect 23707 35037 23719 35071
rect 23661 35031 23719 35037
rect 23937 35071 23995 35077
rect 23937 35037 23949 35071
rect 23983 35037 23995 35071
rect 23937 35031 23995 35037
rect 20073 35007 20131 35013
rect 23952 35000 23980 35031
rect 19208 34972 19838 35000
rect 20824 34972 23980 35000
rect 19208 34960 19214 34972
rect 14108 34904 14412 34932
rect 14458 34892 14464 34944
rect 14516 34932 14522 34944
rect 15105 34935 15163 34941
rect 15105 34932 15117 34935
rect 14516 34904 15117 34932
rect 14516 34892 14522 34904
rect 15105 34901 15117 34904
rect 15151 34901 15163 34935
rect 15105 34895 15163 34901
rect 16669 34935 16727 34941
rect 16669 34901 16681 34935
rect 16715 34932 16727 34935
rect 16850 34932 16856 34944
rect 16715 34904 16856 34932
rect 16715 34901 16727 34904
rect 16669 34895 16727 34901
rect 16850 34892 16856 34904
rect 16908 34892 16914 34944
rect 17954 34892 17960 34944
rect 18012 34932 18018 34944
rect 18138 34932 18144 34944
rect 18012 34904 18144 34932
rect 18012 34892 18018 34904
rect 18138 34892 18144 34904
rect 18196 34892 18202 34944
rect 19518 34892 19524 34944
rect 19576 34892 19582 34944
rect 20824 34941 20852 34972
rect 20809 34935 20867 34941
rect 20809 34901 20821 34935
rect 20855 34901 20867 34935
rect 20809 34895 20867 34901
rect 23474 34892 23480 34944
rect 23532 34892 23538 34944
rect 24121 34935 24179 34941
rect 24121 34901 24133 34935
rect 24167 34932 24179 34935
rect 25222 34932 25228 34944
rect 24167 34904 25228 34932
rect 24167 34901 24179 34904
rect 24121 34895 24179 34901
rect 25222 34892 25228 34904
rect 25280 34892 25286 34944
rect 1104 34842 25000 34864
rect 1104 34790 6884 34842
rect 6936 34790 6948 34842
rect 7000 34790 7012 34842
rect 7064 34790 7076 34842
rect 7128 34790 7140 34842
rect 7192 34790 12818 34842
rect 12870 34790 12882 34842
rect 12934 34790 12946 34842
rect 12998 34790 13010 34842
rect 13062 34790 13074 34842
rect 13126 34790 18752 34842
rect 18804 34790 18816 34842
rect 18868 34790 18880 34842
rect 18932 34790 18944 34842
rect 18996 34790 19008 34842
rect 19060 34790 24686 34842
rect 24738 34790 24750 34842
rect 24802 34790 24814 34842
rect 24866 34790 24878 34842
rect 24930 34790 24942 34842
rect 24994 34790 25000 34842
rect 1104 34768 25000 34790
rect 2130 34688 2136 34740
rect 2188 34728 2194 34740
rect 2409 34731 2467 34737
rect 2409 34728 2421 34731
rect 2188 34700 2421 34728
rect 2188 34688 2194 34700
rect 2409 34697 2421 34700
rect 2455 34697 2467 34731
rect 2409 34691 2467 34697
rect 4338 34688 4344 34740
rect 4396 34728 4402 34740
rect 4525 34731 4583 34737
rect 4525 34728 4537 34731
rect 4396 34700 4537 34728
rect 4396 34688 4402 34700
rect 4525 34697 4537 34700
rect 4571 34697 4583 34731
rect 4525 34691 4583 34697
rect 4614 34688 4620 34740
rect 4672 34728 4678 34740
rect 4982 34728 4988 34740
rect 4672 34700 4988 34728
rect 4672 34688 4678 34700
rect 4982 34688 4988 34700
rect 5040 34688 5046 34740
rect 5074 34688 5080 34740
rect 5132 34728 5138 34740
rect 8938 34728 8944 34740
rect 5132 34700 8944 34728
rect 5132 34688 5138 34700
rect 8938 34688 8944 34700
rect 8996 34688 9002 34740
rect 9030 34688 9036 34740
rect 9088 34688 9094 34740
rect 9214 34688 9220 34740
rect 9272 34728 9278 34740
rect 9858 34728 9864 34740
rect 9272 34700 9864 34728
rect 9272 34688 9278 34700
rect 9858 34688 9864 34700
rect 9916 34688 9922 34740
rect 9950 34688 9956 34740
rect 10008 34728 10014 34740
rect 10410 34728 10416 34740
rect 10008 34700 10416 34728
rect 10008 34688 10014 34700
rect 10410 34688 10416 34700
rect 10468 34688 10474 34740
rect 11054 34688 11060 34740
rect 11112 34688 11118 34740
rect 11882 34688 11888 34740
rect 11940 34728 11946 34740
rect 12618 34728 12624 34740
rect 11940 34700 12624 34728
rect 11940 34688 11946 34700
rect 12618 34688 12624 34700
rect 12676 34688 12682 34740
rect 15197 34731 15255 34737
rect 15197 34697 15209 34731
rect 15243 34728 15255 34731
rect 15286 34728 15292 34740
rect 15243 34700 15292 34728
rect 15243 34697 15255 34700
rect 15197 34691 15255 34697
rect 15286 34688 15292 34700
rect 15344 34688 15350 34740
rect 15378 34688 15384 34740
rect 15436 34728 15442 34740
rect 16945 34731 17003 34737
rect 16945 34728 16957 34731
rect 15436 34700 16957 34728
rect 15436 34688 15442 34700
rect 16945 34697 16957 34700
rect 16991 34697 17003 34731
rect 16945 34691 17003 34697
rect 18785 34731 18843 34737
rect 18785 34697 18797 34731
rect 18831 34728 18843 34731
rect 19150 34728 19156 34740
rect 18831 34700 19156 34728
rect 18831 34697 18843 34700
rect 18785 34691 18843 34697
rect 19150 34688 19156 34700
rect 19208 34688 19214 34740
rect 21453 34731 21511 34737
rect 19306 34700 21128 34728
rect 3053 34663 3111 34669
rect 3053 34629 3065 34663
rect 3099 34660 3111 34663
rect 8478 34660 8484 34672
rect 3099 34632 8484 34660
rect 3099 34629 3111 34632
rect 3053 34623 3111 34629
rect 8478 34620 8484 34632
rect 8536 34620 8542 34672
rect 9674 34660 9680 34672
rect 9324 34632 9680 34660
rect 1578 34592 1584 34604
rect 1412 34564 1584 34592
rect 1412 34536 1440 34564
rect 1578 34552 1584 34564
rect 1636 34552 1642 34604
rect 1671 34595 1729 34601
rect 1671 34561 1683 34595
rect 1717 34592 1729 34595
rect 2038 34592 2044 34604
rect 1717 34564 2044 34592
rect 1717 34561 1729 34564
rect 1671 34555 1729 34561
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 2314 34552 2320 34604
rect 2372 34552 2378 34604
rect 2774 34552 2780 34604
rect 2832 34552 2838 34604
rect 3787 34595 3845 34601
rect 3787 34561 3799 34595
rect 3833 34592 3845 34595
rect 3878 34592 3884 34604
rect 3833 34564 3884 34592
rect 3833 34561 3845 34564
rect 3787 34555 3845 34561
rect 3878 34552 3884 34564
rect 3936 34552 3942 34604
rect 4154 34552 4160 34604
rect 4212 34592 4218 34604
rect 4893 34595 4951 34601
rect 4893 34592 4905 34595
rect 4212 34564 4905 34592
rect 4212 34552 4218 34564
rect 4893 34561 4905 34564
rect 4939 34561 4951 34595
rect 4893 34555 4951 34561
rect 5074 34552 5080 34604
rect 5132 34592 5138 34604
rect 5169 34595 5227 34601
rect 5169 34592 5181 34595
rect 5132 34564 5181 34592
rect 5132 34552 5138 34564
rect 5169 34561 5181 34564
rect 5215 34561 5227 34595
rect 5169 34555 5227 34561
rect 5442 34552 5448 34604
rect 5500 34552 5506 34604
rect 5718 34552 5724 34604
rect 5776 34592 5782 34604
rect 9324 34601 9352 34632
rect 9674 34620 9680 34632
rect 9732 34620 9738 34672
rect 10042 34620 10048 34672
rect 10100 34620 10106 34672
rect 10686 34620 10692 34672
rect 10744 34660 10750 34672
rect 16482 34660 16488 34672
rect 10744 34632 16488 34660
rect 10744 34620 10750 34632
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 16850 34660 16856 34672
rect 16684 34632 16856 34660
rect 6639 34595 6697 34601
rect 6639 34592 6651 34595
rect 5776 34564 6651 34592
rect 5776 34552 5782 34564
rect 6639 34561 6651 34564
rect 6685 34592 6697 34595
rect 8757 34595 8815 34601
rect 6685 34564 7052 34592
rect 6685 34561 6697 34564
rect 6639 34555 6697 34561
rect 1394 34484 1400 34536
rect 1452 34484 1458 34536
rect 2332 34524 2360 34552
rect 3513 34527 3571 34533
rect 3513 34524 3525 34527
rect 2332 34496 3525 34524
rect 3513 34493 3525 34496
rect 3559 34493 3571 34527
rect 3513 34487 3571 34493
rect 4522 34484 4528 34536
rect 4580 34524 4586 34536
rect 5460 34524 5488 34552
rect 6178 34524 6184 34536
rect 4580 34496 6184 34524
rect 4580 34484 4586 34496
rect 6178 34484 6184 34496
rect 6236 34524 6242 34536
rect 6365 34527 6423 34533
rect 6365 34524 6377 34527
rect 6236 34496 6377 34524
rect 6236 34484 6242 34496
rect 6365 34493 6377 34496
rect 6411 34493 6423 34527
rect 6365 34487 6423 34493
rect 2222 34416 2228 34468
rect 2280 34456 2286 34468
rect 3326 34456 3332 34468
rect 2280 34428 3332 34456
rect 2280 34416 2286 34428
rect 3326 34416 3332 34428
rect 3384 34416 3390 34468
rect 4614 34416 4620 34468
rect 4672 34456 4678 34468
rect 4982 34456 4988 34468
rect 4672 34428 4988 34456
rect 4672 34416 4678 34428
rect 4982 34416 4988 34428
rect 5040 34416 5046 34468
rect 7024 34456 7052 34564
rect 8757 34561 8769 34595
rect 8803 34592 8815 34595
rect 9309 34595 9367 34601
rect 9493 34598 9551 34601
rect 9309 34592 9321 34595
rect 8803 34564 9321 34592
rect 8803 34561 8815 34564
rect 8757 34555 8815 34561
rect 9309 34561 9321 34564
rect 9355 34561 9367 34595
rect 9309 34555 9367 34561
rect 9416 34595 9551 34598
rect 9416 34570 9505 34595
rect 9033 34527 9091 34533
rect 9033 34493 9045 34527
rect 9079 34524 9091 34527
rect 9079 34496 9168 34524
rect 9079 34493 9091 34496
rect 9033 34487 9091 34493
rect 7024 34428 7512 34456
rect 7484 34400 7512 34428
rect 1210 34348 1216 34400
rect 1268 34388 1274 34400
rect 2498 34388 2504 34400
rect 1268 34360 2504 34388
rect 1268 34348 1274 34360
rect 2498 34348 2504 34360
rect 2556 34348 2562 34400
rect 3602 34348 3608 34400
rect 3660 34388 3666 34400
rect 3878 34388 3884 34400
rect 3660 34360 3884 34388
rect 3660 34348 3666 34360
rect 3878 34348 3884 34360
rect 3936 34388 3942 34400
rect 5442 34388 5448 34400
rect 3936 34360 5448 34388
rect 3936 34348 3942 34360
rect 5442 34348 5448 34360
rect 5500 34348 5506 34400
rect 7374 34348 7380 34400
rect 7432 34348 7438 34400
rect 7466 34348 7472 34400
rect 7524 34348 7530 34400
rect 7650 34348 7656 34400
rect 7708 34388 7714 34400
rect 8110 34388 8116 34400
rect 7708 34360 8116 34388
rect 7708 34348 7714 34360
rect 8110 34348 8116 34360
rect 8168 34348 8174 34400
rect 8849 34391 8907 34397
rect 8849 34357 8861 34391
rect 8895 34388 8907 34391
rect 9030 34388 9036 34400
rect 8895 34360 9036 34388
rect 8895 34357 8907 34360
rect 8849 34351 8907 34357
rect 9030 34348 9036 34360
rect 9088 34348 9094 34400
rect 9140 34388 9168 34496
rect 9214 34484 9220 34536
rect 9272 34524 9278 34536
rect 9416 34524 9444 34570
rect 9493 34561 9505 34570
rect 9539 34561 9551 34595
rect 9493 34555 9551 34561
rect 9582 34552 9588 34604
rect 9640 34552 9646 34604
rect 10060 34592 10088 34620
rect 10287 34595 10345 34601
rect 10287 34592 10299 34595
rect 10060 34564 10299 34592
rect 10287 34561 10299 34564
rect 10333 34561 10345 34595
rect 10287 34555 10345 34561
rect 10410 34552 10416 34604
rect 10468 34592 10474 34604
rect 13446 34592 13452 34604
rect 10468 34564 13452 34592
rect 10468 34552 10474 34564
rect 13446 34552 13452 34564
rect 13504 34552 13510 34604
rect 13722 34552 13728 34604
rect 13780 34592 13786 34604
rect 16684 34601 16712 34632
rect 16850 34620 16856 34632
rect 16908 34660 16914 34672
rect 16908 34632 17356 34660
rect 16908 34620 16914 34632
rect 14459 34595 14517 34601
rect 14459 34592 14471 34595
rect 13780 34564 14471 34592
rect 13780 34552 13786 34564
rect 14459 34561 14471 34564
rect 14505 34592 14517 34595
rect 16669 34595 16727 34601
rect 14505 34564 15332 34592
rect 14505 34561 14517 34564
rect 14459 34555 14517 34561
rect 9272 34496 9444 34524
rect 9272 34484 9278 34496
rect 9766 34484 9772 34536
rect 9824 34524 9830 34536
rect 10042 34524 10048 34536
rect 9824 34496 10048 34524
rect 9824 34484 9830 34496
rect 10042 34484 10048 34496
rect 10100 34484 10106 34536
rect 14090 34484 14096 34536
rect 14148 34524 14154 34536
rect 14185 34527 14243 34533
rect 14185 34524 14197 34527
rect 14148 34496 14197 34524
rect 14148 34484 14154 34496
rect 14185 34493 14197 34496
rect 14231 34493 14243 34527
rect 15304 34524 15332 34564
rect 16669 34561 16681 34595
rect 16715 34561 16727 34595
rect 16669 34555 16727 34561
rect 17034 34552 17040 34604
rect 17092 34552 17098 34604
rect 17328 34601 17356 34632
rect 17402 34620 17408 34672
rect 17460 34660 17466 34672
rect 19306 34660 19334 34700
rect 17460 34632 19334 34660
rect 17460 34620 17466 34632
rect 19518 34620 19524 34672
rect 19576 34620 19582 34672
rect 20438 34620 20444 34672
rect 20496 34660 20502 34672
rect 21100 34660 21128 34700
rect 21453 34697 21465 34731
rect 21499 34728 21511 34731
rect 21499 34700 23428 34728
rect 21499 34697 21511 34700
rect 21453 34691 21511 34697
rect 20496 34632 21036 34660
rect 21100 34632 21680 34660
rect 20496 34620 20502 34632
rect 17313 34595 17371 34601
rect 17313 34561 17325 34595
rect 17359 34561 17371 34595
rect 17313 34555 17371 34561
rect 17494 34552 17500 34604
rect 17552 34552 17558 34604
rect 18969 34595 19027 34601
rect 18969 34561 18981 34595
rect 19015 34561 19027 34595
rect 18969 34555 19027 34561
rect 19061 34595 19119 34601
rect 19061 34561 19073 34595
rect 19107 34592 19119 34595
rect 19150 34592 19156 34604
rect 19107 34564 19156 34592
rect 19107 34561 19119 34564
rect 19061 34555 19119 34561
rect 16945 34527 17003 34533
rect 15304 34496 16712 34524
rect 14185 34487 14243 34493
rect 9401 34391 9459 34397
rect 9401 34388 9413 34391
rect 9140 34360 9413 34388
rect 9401 34357 9413 34360
rect 9447 34357 9459 34391
rect 9401 34351 9459 34357
rect 9490 34348 9496 34400
rect 9548 34388 9554 34400
rect 9677 34391 9735 34397
rect 9677 34388 9689 34391
rect 9548 34360 9689 34388
rect 9548 34348 9554 34360
rect 9677 34357 9689 34360
rect 9723 34357 9735 34391
rect 9677 34351 9735 34357
rect 9858 34348 9864 34400
rect 9916 34388 9922 34400
rect 10870 34388 10876 34400
rect 9916 34360 10876 34388
rect 9916 34348 9922 34360
rect 10870 34348 10876 34360
rect 10928 34348 10934 34400
rect 16684 34388 16712 34496
rect 16945 34493 16957 34527
rect 16991 34524 17003 34527
rect 17405 34527 17463 34533
rect 17405 34524 17417 34527
rect 16991 34496 17417 34524
rect 16991 34493 17003 34496
rect 16945 34487 17003 34493
rect 17405 34493 17417 34496
rect 17451 34493 17463 34527
rect 18984 34524 19012 34555
rect 19150 34552 19156 34564
rect 19208 34552 19214 34604
rect 19334 34601 19340 34604
rect 19328 34592 19340 34601
rect 19295 34564 19340 34592
rect 19328 34555 19340 34564
rect 19334 34552 19340 34555
rect 19392 34552 19398 34604
rect 19536 34592 19564 34620
rect 21008 34601 21036 34632
rect 21652 34601 21680 34632
rect 22079 34625 22137 34631
rect 20533 34595 20591 34601
rect 20533 34592 20545 34595
rect 19536 34564 20545 34592
rect 20533 34561 20545 34564
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 21637 34595 21695 34601
rect 21637 34561 21649 34595
rect 21683 34561 21695 34595
rect 22079 34591 22091 34625
rect 22125 34622 22137 34625
rect 22125 34592 22140 34622
rect 22186 34592 22192 34604
rect 22125 34591 22192 34592
rect 22079 34585 22192 34591
rect 22112 34564 22192 34585
rect 21637 34555 21695 34561
rect 22186 34552 22192 34564
rect 22244 34552 22250 34604
rect 23400 34601 23428 34700
rect 23658 34688 23664 34740
rect 23716 34688 23722 34740
rect 23750 34688 23756 34740
rect 23808 34728 23814 34740
rect 23808 34700 24164 34728
rect 23808 34688 23814 34700
rect 23934 34620 23940 34672
rect 23992 34620 23998 34672
rect 24136 34669 24164 34700
rect 24121 34663 24179 34669
rect 24121 34629 24133 34663
rect 24167 34629 24179 34663
rect 24121 34623 24179 34629
rect 23385 34595 23443 34601
rect 23385 34561 23397 34595
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 23750 34552 23756 34604
rect 23808 34592 23814 34604
rect 23845 34595 23903 34601
rect 23845 34592 23857 34595
rect 23808 34564 23857 34592
rect 23808 34552 23814 34564
rect 23845 34561 23857 34564
rect 23891 34561 23903 34595
rect 23845 34555 23903 34561
rect 17405 34487 17463 34493
rect 17512 34496 19012 34524
rect 20625 34527 20683 34533
rect 16761 34459 16819 34465
rect 16761 34425 16773 34459
rect 16807 34456 16819 34459
rect 17129 34459 17187 34465
rect 17129 34456 17141 34459
rect 16807 34428 17141 34456
rect 16807 34425 16819 34428
rect 16761 34419 16819 34425
rect 17129 34425 17141 34428
rect 17175 34425 17187 34459
rect 17129 34419 17187 34425
rect 17512 34388 17540 34496
rect 20625 34493 20637 34527
rect 20671 34524 20683 34527
rect 21082 34524 21088 34536
rect 20671 34496 21088 34524
rect 20671 34493 20683 34496
rect 20625 34487 20683 34493
rect 21082 34484 21088 34496
rect 21140 34484 21146 34536
rect 21821 34527 21879 34533
rect 21821 34524 21833 34527
rect 21192 34496 21833 34524
rect 21192 34456 21220 34496
rect 21821 34493 21833 34496
rect 21867 34493 21879 34527
rect 23952 34524 23980 34620
rect 21821 34487 21879 34493
rect 23216 34496 23980 34524
rect 23216 34465 23244 34496
rect 24394 34484 24400 34536
rect 24452 34484 24458 34536
rect 19996 34428 21220 34456
rect 23201 34459 23259 34465
rect 19996 34400 20024 34428
rect 23201 34425 23213 34459
rect 23247 34425 23259 34459
rect 23201 34419 23259 34425
rect 16684 34360 17540 34388
rect 19978 34348 19984 34400
rect 20036 34348 20042 34400
rect 20438 34348 20444 34400
rect 20496 34348 20502 34400
rect 20809 34391 20867 34397
rect 20809 34357 20821 34391
rect 20855 34388 20867 34391
rect 21542 34388 21548 34400
rect 20855 34360 21548 34388
rect 20855 34357 20867 34360
rect 20809 34351 20867 34357
rect 21542 34348 21548 34360
rect 21600 34348 21606 34400
rect 22833 34391 22891 34397
rect 22833 34357 22845 34391
rect 22879 34388 22891 34391
rect 23106 34388 23112 34400
rect 22879 34360 23112 34388
rect 22879 34357 22891 34360
rect 22833 34351 22891 34357
rect 23106 34348 23112 34360
rect 23164 34348 23170 34400
rect 1104 34298 24840 34320
rect 1104 34246 3917 34298
rect 3969 34246 3981 34298
rect 4033 34246 4045 34298
rect 4097 34246 4109 34298
rect 4161 34246 4173 34298
rect 4225 34246 9851 34298
rect 9903 34246 9915 34298
rect 9967 34246 9979 34298
rect 10031 34246 10043 34298
rect 10095 34246 10107 34298
rect 10159 34246 15785 34298
rect 15837 34246 15849 34298
rect 15901 34246 15913 34298
rect 15965 34246 15977 34298
rect 16029 34246 16041 34298
rect 16093 34246 21719 34298
rect 21771 34246 21783 34298
rect 21835 34246 21847 34298
rect 21899 34246 21911 34298
rect 21963 34246 21975 34298
rect 22027 34246 24840 34298
rect 1104 34224 24840 34246
rect 2406 34144 2412 34196
rect 2464 34184 2470 34196
rect 3050 34184 3056 34196
rect 2464 34156 3056 34184
rect 2464 34144 2470 34156
rect 3050 34144 3056 34156
rect 3108 34144 3114 34196
rect 5718 34184 5724 34196
rect 4264 34156 5724 34184
rect 2590 34076 2596 34128
rect 2648 34116 2654 34128
rect 3970 34116 3976 34128
rect 2648 34088 3976 34116
rect 2648 34076 2654 34088
rect 3970 34076 3976 34088
rect 4028 34076 4034 34128
rect 2958 34048 2964 34060
rect 2700 34020 2964 34048
rect 842 33940 848 33992
rect 900 33980 906 33992
rect 1394 33980 1400 33992
rect 900 33952 1400 33980
rect 900 33940 906 33952
rect 1394 33940 1400 33952
rect 1452 33940 1458 33992
rect 1671 33983 1729 33989
rect 1671 33949 1683 33983
rect 1717 33980 1729 33983
rect 2700 33980 2728 34020
rect 2958 34008 2964 34020
rect 3016 34008 3022 34060
rect 3053 34051 3111 34057
rect 3053 34017 3065 34051
rect 3099 34048 3111 34051
rect 4264 34048 4292 34156
rect 5718 34144 5724 34156
rect 5776 34144 5782 34196
rect 6288 34156 9628 34184
rect 3099 34020 4292 34048
rect 3099 34017 3111 34020
rect 3053 34011 3111 34017
rect 4522 34008 4528 34060
rect 4580 34008 4586 34060
rect 1717 33952 2728 33980
rect 1717 33949 1729 33952
rect 1671 33943 1729 33949
rect 2774 33940 2780 33992
rect 2832 33940 2838 33992
rect 3789 33983 3847 33989
rect 3789 33980 3801 33983
rect 2976 33952 3801 33980
rect 1210 33872 1216 33924
rect 1268 33912 1274 33924
rect 2976 33912 3004 33952
rect 3789 33949 3801 33952
rect 3835 33949 3847 33983
rect 4767 33983 4825 33989
rect 4767 33980 4779 33983
rect 3789 33943 3847 33949
rect 3988 33952 4779 33980
rect 1268 33884 3004 33912
rect 1268 33872 1274 33884
rect 3326 33872 3332 33924
rect 3384 33912 3390 33924
rect 3988 33912 4016 33952
rect 4767 33949 4779 33952
rect 4813 33980 4825 33983
rect 6288 33980 6316 34156
rect 7374 34076 7380 34128
rect 7432 34116 7438 34128
rect 7469 34119 7527 34125
rect 7469 34116 7481 34119
rect 7432 34088 7481 34116
rect 7432 34076 7438 34088
rect 7469 34085 7481 34088
rect 7515 34085 7527 34119
rect 7469 34079 7527 34085
rect 6362 34008 6368 34060
rect 6420 34048 6426 34060
rect 7883 34051 7941 34057
rect 6420 34020 7788 34048
rect 6420 34008 6426 34020
rect 4813 33952 6316 33980
rect 4813 33949 4825 33952
rect 4767 33943 4825 33949
rect 6730 33940 6736 33992
rect 6788 33980 6794 33992
rect 7760 33989 7788 34020
rect 7883 34017 7895 34051
rect 7929 34048 7941 34051
rect 8754 34048 8760 34060
rect 7929 34020 8760 34048
rect 7929 34017 7941 34020
rect 7883 34011 7941 34017
rect 8754 34008 8760 34020
rect 8812 34008 8818 34060
rect 6825 33983 6883 33989
rect 6825 33980 6837 33983
rect 6788 33952 6837 33980
rect 6788 33940 6794 33952
rect 6825 33949 6837 33952
rect 6871 33949 6883 33983
rect 6825 33943 6883 33949
rect 7009 33983 7067 33989
rect 7009 33949 7021 33983
rect 7055 33949 7067 33983
rect 7009 33943 7067 33949
rect 7745 33983 7803 33989
rect 7745 33949 7757 33983
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 3384 33884 4016 33912
rect 4065 33915 4123 33921
rect 3384 33872 3390 33884
rect 4065 33881 4077 33915
rect 4111 33912 4123 33915
rect 6270 33912 6276 33924
rect 4111 33884 6276 33912
rect 4111 33881 4123 33884
rect 4065 33875 4123 33881
rect 6270 33872 6276 33884
rect 6328 33872 6334 33924
rect 2130 33804 2136 33856
rect 2188 33844 2194 33856
rect 2409 33847 2467 33853
rect 2409 33844 2421 33847
rect 2188 33816 2421 33844
rect 2188 33804 2194 33816
rect 2409 33813 2421 33816
rect 2455 33813 2467 33847
rect 2409 33807 2467 33813
rect 5534 33804 5540 33856
rect 5592 33804 5598 33856
rect 7024 33844 7052 33943
rect 8018 33940 8024 33992
rect 8076 33940 8082 33992
rect 8938 33940 8944 33992
rect 8996 33940 9002 33992
rect 9183 33983 9241 33989
rect 9183 33980 9195 33983
rect 9048 33952 9195 33980
rect 9048 33912 9076 33952
rect 9183 33949 9195 33952
rect 9229 33949 9241 33983
rect 9183 33943 9241 33949
rect 8496 33884 9076 33912
rect 9600 33912 9628 34156
rect 9674 34144 9680 34196
rect 9732 34184 9738 34196
rect 9953 34187 10011 34193
rect 9953 34184 9965 34187
rect 9732 34156 9965 34184
rect 9732 34144 9738 34156
rect 9953 34153 9965 34156
rect 9999 34153 10011 34187
rect 9953 34147 10011 34153
rect 14366 34144 14372 34196
rect 14424 34184 14430 34196
rect 17313 34187 17371 34193
rect 14424 34156 17264 34184
rect 14424 34144 14430 34156
rect 10962 34116 10968 34128
rect 9692 34088 10968 34116
rect 9692 34060 9720 34088
rect 10962 34076 10968 34088
rect 11020 34076 11026 34128
rect 13538 34076 13544 34128
rect 13596 34076 13602 34128
rect 17236 34116 17264 34156
rect 17313 34153 17325 34187
rect 17359 34184 17371 34187
rect 17494 34184 17500 34196
rect 17359 34156 17500 34184
rect 17359 34153 17371 34156
rect 17313 34147 17371 34153
rect 17494 34144 17500 34156
rect 17552 34144 17558 34196
rect 17586 34144 17592 34196
rect 17644 34184 17650 34196
rect 19886 34184 19892 34196
rect 17644 34156 19892 34184
rect 17644 34144 17650 34156
rect 17236 34088 19334 34116
rect 9674 34008 9680 34060
rect 9732 34008 9738 34060
rect 13998 34008 14004 34060
rect 14056 34008 14062 34060
rect 15194 34008 15200 34060
rect 15252 34048 15258 34060
rect 15933 34051 15991 34057
rect 15933 34048 15945 34051
rect 15252 34020 15945 34048
rect 15252 34008 15258 34020
rect 15933 34017 15945 34020
rect 15979 34017 15991 34051
rect 15933 34011 15991 34017
rect 17696 34020 18184 34048
rect 10226 33940 10232 33992
rect 10284 33980 10290 33992
rect 11882 33980 11888 33992
rect 10284 33952 11888 33980
rect 10284 33940 10290 33952
rect 11882 33940 11888 33952
rect 11940 33980 11946 33992
rect 12529 33983 12587 33989
rect 12529 33980 12541 33983
rect 11940 33952 12541 33980
rect 11940 33940 11946 33952
rect 12529 33949 12541 33952
rect 12575 33949 12587 33983
rect 12529 33943 12587 33949
rect 12803 33983 12861 33989
rect 12803 33949 12815 33983
rect 12849 33980 12861 33983
rect 13630 33980 13636 33992
rect 12849 33952 13636 33980
rect 12849 33949 12861 33952
rect 12803 33943 12861 33949
rect 13630 33940 13636 33952
rect 13688 33940 13694 33992
rect 14016 33980 14044 34008
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 14016 33952 14105 33980
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 14335 33983 14393 33989
rect 14335 33980 14347 33983
rect 14093 33943 14151 33949
rect 14200 33952 14347 33980
rect 14200 33912 14228 33952
rect 14335 33949 14347 33952
rect 14381 33980 14393 33983
rect 14381 33952 14780 33980
rect 14381 33949 14393 33952
rect 14335 33943 14393 33949
rect 9600 33884 14228 33912
rect 14752 33912 14780 33952
rect 14826 33940 14832 33992
rect 14884 33980 14890 33992
rect 15102 33980 15108 33992
rect 14884 33952 15108 33980
rect 14884 33940 14890 33952
rect 15102 33940 15108 33952
rect 15160 33940 15166 33992
rect 16175 33983 16233 33989
rect 16175 33980 16187 33983
rect 15396 33952 16187 33980
rect 15396 33924 15424 33952
rect 16175 33949 16187 33952
rect 16221 33980 16233 33983
rect 16758 33980 16764 33992
rect 16221 33952 16764 33980
rect 16221 33949 16233 33952
rect 16175 33943 16233 33949
rect 16758 33940 16764 33952
rect 16816 33940 16822 33992
rect 17494 33940 17500 33992
rect 17552 33940 17558 33992
rect 14752 33884 15332 33912
rect 8496 33856 8524 33884
rect 7834 33844 7840 33856
rect 7024 33816 7840 33844
rect 7834 33804 7840 33816
rect 7892 33804 7898 33856
rect 8478 33804 8484 33856
rect 8536 33804 8542 33856
rect 8662 33804 8668 33856
rect 8720 33804 8726 33856
rect 8938 33804 8944 33856
rect 8996 33844 9002 33856
rect 12434 33844 12440 33856
rect 8996 33816 12440 33844
rect 8996 33804 9002 33816
rect 12434 33804 12440 33816
rect 12492 33804 12498 33856
rect 13170 33804 13176 33856
rect 13228 33844 13234 33856
rect 14366 33844 14372 33856
rect 13228 33816 14372 33844
rect 13228 33804 13234 33816
rect 14366 33804 14372 33816
rect 14424 33804 14430 33856
rect 14918 33804 14924 33856
rect 14976 33844 14982 33856
rect 15105 33847 15163 33853
rect 15105 33844 15117 33847
rect 14976 33816 15117 33844
rect 14976 33804 14982 33816
rect 15105 33813 15117 33816
rect 15151 33813 15163 33847
rect 15304 33844 15332 33884
rect 15378 33872 15384 33924
rect 15436 33872 15442 33924
rect 17402 33912 17408 33924
rect 16868 33884 17408 33912
rect 16868 33844 16896 33884
rect 17402 33872 17408 33884
rect 17460 33872 17466 33924
rect 15304 33816 16896 33844
rect 15105 33807 15163 33813
rect 16942 33804 16948 33856
rect 17000 33804 17006 33856
rect 17696 33853 17724 34020
rect 18156 33989 18184 34020
rect 17865 33983 17923 33989
rect 17865 33980 17877 33983
rect 17788 33952 17877 33980
rect 17788 33856 17816 33952
rect 17865 33949 17877 33952
rect 17911 33949 17923 33983
rect 17865 33943 17923 33949
rect 18141 33983 18199 33989
rect 18141 33949 18153 33983
rect 18187 33949 18199 33983
rect 19306 33980 19334 34088
rect 19628 34057 19656 34156
rect 19886 34144 19892 34156
rect 19944 34144 19950 34196
rect 21082 34144 21088 34196
rect 21140 34144 21146 34196
rect 22373 34187 22431 34193
rect 22373 34153 22385 34187
rect 22419 34184 22431 34187
rect 23382 34184 23388 34196
rect 22419 34156 23388 34184
rect 22419 34153 22431 34156
rect 22373 34147 22431 34153
rect 23382 34144 23388 34156
rect 23440 34144 23446 34196
rect 20625 34119 20683 34125
rect 20625 34085 20637 34119
rect 20671 34085 20683 34119
rect 20625 34079 20683 34085
rect 23109 34119 23167 34125
rect 23109 34085 23121 34119
rect 23155 34085 23167 34119
rect 23109 34079 23167 34085
rect 19613 34051 19671 34057
rect 19613 34017 19625 34051
rect 19659 34017 19671 34051
rect 19613 34011 19671 34017
rect 19887 33983 19945 33989
rect 19887 33980 19899 33983
rect 19306 33952 19899 33980
rect 18141 33943 18199 33949
rect 19887 33949 19899 33952
rect 19933 33980 19945 33983
rect 20254 33980 20260 33992
rect 19933 33952 20260 33980
rect 19933 33949 19945 33952
rect 19887 33943 19945 33949
rect 20254 33940 20260 33952
rect 20312 33940 20318 33992
rect 20640 33980 20668 34079
rect 21269 34051 21327 34057
rect 21269 34017 21281 34051
rect 21315 34048 21327 34051
rect 21453 34051 21511 34057
rect 21453 34048 21465 34051
rect 21315 34020 21465 34048
rect 21315 34017 21327 34020
rect 21269 34011 21327 34017
rect 21453 34017 21465 34020
rect 21499 34017 21511 34051
rect 23124 34048 23152 34079
rect 23124 34020 23980 34048
rect 21453 34011 21511 34017
rect 20993 33983 21051 33989
rect 20993 33980 21005 33983
rect 20640 33952 21005 33980
rect 20993 33949 21005 33952
rect 21039 33980 21051 33983
rect 21361 33983 21419 33989
rect 21361 33980 21373 33983
rect 21039 33952 21373 33980
rect 21039 33949 21051 33952
rect 20993 33943 21051 33949
rect 21361 33949 21373 33952
rect 21407 33949 21419 33983
rect 21361 33943 21419 33949
rect 21542 33940 21548 33992
rect 21600 33940 21606 33992
rect 22554 33940 22560 33992
rect 22612 33940 22618 33992
rect 22830 33940 22836 33992
rect 22888 33940 22894 33992
rect 23293 33983 23351 33989
rect 23293 33949 23305 33983
rect 23339 33980 23351 33983
rect 23339 33952 23428 33980
rect 23339 33949 23351 33952
rect 23293 33943 23351 33949
rect 17681 33847 17739 33853
rect 17681 33813 17693 33847
rect 17727 33813 17739 33847
rect 17681 33807 17739 33813
rect 17770 33804 17776 33856
rect 17828 33804 17834 33856
rect 18230 33804 18236 33856
rect 18288 33804 18294 33856
rect 21269 33847 21327 33853
rect 21269 33813 21281 33847
rect 21315 33844 21327 33847
rect 21634 33844 21640 33856
rect 21315 33816 21640 33844
rect 21315 33813 21327 33816
rect 21269 33807 21327 33813
rect 21634 33804 21640 33816
rect 21692 33804 21698 33856
rect 22646 33804 22652 33856
rect 22704 33804 22710 33856
rect 23400 33853 23428 33952
rect 23474 33940 23480 33992
rect 23532 33980 23538 33992
rect 23952 33989 23980 34020
rect 23569 33983 23627 33989
rect 23569 33980 23581 33983
rect 23532 33952 23581 33980
rect 23532 33940 23538 33952
rect 23569 33949 23581 33952
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23845 33983 23903 33989
rect 23845 33949 23857 33983
rect 23891 33949 23903 33983
rect 23845 33943 23903 33949
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 23860 33912 23888 33943
rect 23492 33884 23888 33912
rect 23492 33856 23520 33884
rect 23385 33847 23443 33853
rect 23385 33813 23397 33847
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 23474 33804 23480 33856
rect 23532 33804 23538 33856
rect 23658 33804 23664 33856
rect 23716 33804 23722 33856
rect 24121 33847 24179 33853
rect 24121 33813 24133 33847
rect 24167 33844 24179 33847
rect 25222 33844 25228 33856
rect 24167 33816 25228 33844
rect 24167 33813 24179 33816
rect 24121 33807 24179 33813
rect 25222 33804 25228 33816
rect 25280 33804 25286 33856
rect 1104 33754 25000 33776
rect 1104 33702 6884 33754
rect 6936 33702 6948 33754
rect 7000 33702 7012 33754
rect 7064 33702 7076 33754
rect 7128 33702 7140 33754
rect 7192 33702 12818 33754
rect 12870 33702 12882 33754
rect 12934 33702 12946 33754
rect 12998 33702 13010 33754
rect 13062 33702 13074 33754
rect 13126 33702 18752 33754
rect 18804 33702 18816 33754
rect 18868 33702 18880 33754
rect 18932 33702 18944 33754
rect 18996 33702 19008 33754
rect 19060 33702 24686 33754
rect 24738 33702 24750 33754
rect 24802 33702 24814 33754
rect 24866 33702 24878 33754
rect 24930 33702 24942 33754
rect 24994 33702 25000 33754
rect 1104 33680 25000 33702
rect 1946 33600 1952 33652
rect 2004 33640 2010 33652
rect 3053 33643 3111 33649
rect 2004 33612 3004 33640
rect 2004 33600 2010 33612
rect 1118 33532 1124 33584
rect 1176 33532 1182 33584
rect 2976 33572 3004 33612
rect 3053 33609 3065 33643
rect 3099 33640 3111 33643
rect 3234 33640 3240 33652
rect 3099 33612 3240 33640
rect 3099 33609 3111 33612
rect 3053 33603 3111 33609
rect 3234 33600 3240 33612
rect 3292 33600 3298 33652
rect 3786 33600 3792 33652
rect 3844 33600 3850 33652
rect 4341 33643 4399 33649
rect 4341 33609 4353 33643
rect 4387 33640 4399 33643
rect 8202 33640 8208 33652
rect 4387 33612 8208 33640
rect 4387 33609 4399 33612
rect 4341 33603 4399 33609
rect 8202 33600 8208 33612
rect 8260 33600 8266 33652
rect 8662 33600 8668 33652
rect 8720 33600 8726 33652
rect 8849 33643 8907 33649
rect 8849 33609 8861 33643
rect 8895 33609 8907 33643
rect 8849 33603 8907 33609
rect 9125 33643 9183 33649
rect 9125 33609 9137 33643
rect 9171 33640 9183 33643
rect 9490 33640 9496 33652
rect 9171 33612 9496 33640
rect 9171 33609 9183 33612
rect 9125 33603 9183 33609
rect 3142 33572 3148 33584
rect 2976 33544 3148 33572
rect 3142 33532 3148 33544
rect 3200 33532 3206 33584
rect 3329 33575 3387 33581
rect 3329 33541 3341 33575
rect 3375 33572 3387 33575
rect 3804 33572 3832 33600
rect 3375 33544 3832 33572
rect 3375 33541 3387 33544
rect 3329 33535 3387 33541
rect 3970 33532 3976 33584
rect 4028 33532 4034 33584
rect 4157 33575 4215 33581
rect 4157 33541 4169 33575
rect 4203 33572 4215 33575
rect 4614 33572 4620 33584
rect 4203 33544 4620 33572
rect 4203 33541 4215 33544
rect 4157 33535 4215 33541
rect 4614 33532 4620 33544
rect 4672 33532 4678 33584
rect 4890 33532 4896 33584
rect 4948 33572 4954 33584
rect 4948 33544 5396 33572
rect 4948 33532 4954 33544
rect 1136 33504 1164 33532
rect 1731 33507 1789 33513
rect 1731 33504 1743 33507
rect 1136 33476 1743 33504
rect 1731 33473 1743 33476
rect 1777 33504 1789 33507
rect 2222 33504 2228 33516
rect 1777 33476 2228 33504
rect 1777 33473 1789 33476
rect 1731 33467 1789 33473
rect 2222 33464 2228 33476
rect 2280 33464 2286 33516
rect 3418 33464 3424 33516
rect 3476 33464 3482 33516
rect 3789 33507 3847 33513
rect 3789 33473 3801 33507
rect 3835 33504 3847 33507
rect 3988 33504 4016 33532
rect 5135 33507 5193 33513
rect 5135 33504 5147 33507
rect 3835 33476 4016 33504
rect 4816 33476 5147 33504
rect 3835 33473 3847 33476
rect 3789 33467 3847 33473
rect 1394 33396 1400 33448
rect 1452 33436 1458 33448
rect 1489 33439 1547 33445
rect 1489 33436 1501 33439
rect 1452 33408 1501 33436
rect 1452 33396 1458 33408
rect 1489 33405 1501 33408
rect 1535 33405 1547 33439
rect 1489 33399 1547 33405
rect 2516 33408 2898 33436
rect 2516 33377 2544 33408
rect 4338 33396 4344 33448
rect 4396 33436 4402 33448
rect 4816 33436 4844 33476
rect 5135 33473 5147 33476
rect 5181 33473 5193 33507
rect 5368 33504 5396 33544
rect 6546 33532 6552 33584
rect 6604 33572 6610 33584
rect 6730 33572 6736 33584
rect 6604 33544 6736 33572
rect 6604 33532 6610 33544
rect 6730 33532 6736 33544
rect 6788 33532 6794 33584
rect 5902 33504 5908 33516
rect 5368 33476 5908 33504
rect 5135 33467 5193 33473
rect 5902 33464 5908 33476
rect 5960 33464 5966 33516
rect 7024 33476 7328 33504
rect 7024 33448 7052 33476
rect 4396 33408 4844 33436
rect 4893 33439 4951 33445
rect 4396 33396 4402 33408
rect 4893 33405 4905 33439
rect 4939 33405 4951 33439
rect 4893 33399 4951 33405
rect 2501 33371 2559 33377
rect 2501 33337 2513 33371
rect 2547 33337 2559 33371
rect 2501 33331 2559 33337
rect 4522 33328 4528 33380
rect 4580 33368 4586 33380
rect 4908 33368 4936 33399
rect 6638 33396 6644 33448
rect 6696 33436 6702 33448
rect 6917 33439 6975 33445
rect 6917 33436 6929 33439
rect 6696 33408 6929 33436
rect 6696 33396 6702 33408
rect 6917 33405 6929 33408
rect 6963 33405 6975 33439
rect 6917 33399 6975 33405
rect 7006 33396 7012 33448
rect 7064 33396 7070 33448
rect 7101 33439 7159 33445
rect 7101 33405 7113 33439
rect 7147 33436 7159 33439
rect 7190 33436 7196 33448
rect 7147 33408 7196 33436
rect 7147 33405 7159 33408
rect 7101 33399 7159 33405
rect 7190 33396 7196 33408
rect 7248 33396 7254 33448
rect 7300 33436 7328 33476
rect 8110 33464 8116 33516
rect 8168 33464 8174 33516
rect 8680 33504 8708 33600
rect 8864 33572 8892 33603
rect 9490 33600 9496 33612
rect 9548 33600 9554 33652
rect 9674 33640 9680 33652
rect 9646 33600 9680 33640
rect 9732 33600 9738 33652
rect 10686 33640 10692 33652
rect 9782 33612 10692 33640
rect 9214 33572 9220 33584
rect 8864 33544 9220 33572
rect 9214 33532 9220 33544
rect 9272 33532 9278 33584
rect 9033 33507 9091 33513
rect 9033 33504 9045 33507
rect 8680 33476 9045 33504
rect 9033 33473 9045 33476
rect 9079 33473 9091 33507
rect 9033 33467 9091 33473
rect 9309 33507 9367 33513
rect 9309 33473 9321 33507
rect 9355 33473 9367 33507
rect 9646 33504 9674 33600
rect 9782 33513 9810 33612
rect 10686 33600 10692 33612
rect 10744 33600 10750 33652
rect 15378 33640 15384 33652
rect 11072 33612 15384 33640
rect 11072 33584 11100 33612
rect 15378 33600 15384 33612
rect 15436 33600 15442 33652
rect 16945 33643 17003 33649
rect 16945 33609 16957 33643
rect 16991 33640 17003 33643
rect 17034 33640 17040 33652
rect 16991 33612 17040 33640
rect 16991 33609 17003 33612
rect 16945 33603 17003 33609
rect 17034 33600 17040 33612
rect 17092 33600 17098 33652
rect 18874 33640 18880 33652
rect 17144 33612 18880 33640
rect 11054 33532 11060 33584
rect 11112 33532 11118 33584
rect 13633 33575 13691 33581
rect 13633 33541 13645 33575
rect 13679 33572 13691 33575
rect 17144 33572 17172 33612
rect 18874 33600 18880 33612
rect 18932 33600 18938 33652
rect 19058 33600 19064 33652
rect 19116 33640 19122 33652
rect 20990 33640 20996 33652
rect 19116 33612 20996 33640
rect 19116 33600 19122 33612
rect 20990 33600 20996 33612
rect 21048 33600 21054 33652
rect 22646 33600 22652 33652
rect 22704 33600 22710 33652
rect 22830 33600 22836 33652
rect 22888 33640 22894 33652
rect 23201 33643 23259 33649
rect 23201 33640 23213 33643
rect 22888 33612 23213 33640
rect 22888 33600 22894 33612
rect 23201 33609 23213 33612
rect 23247 33609 23259 33643
rect 23201 33603 23259 33609
rect 23658 33600 23664 33652
rect 23716 33600 23722 33652
rect 17678 33572 17684 33584
rect 13679 33544 17172 33572
rect 17236 33544 17684 33572
rect 13679 33541 13691 33544
rect 13633 33535 13691 33541
rect 9309 33467 9367 33473
rect 9416 33476 9674 33504
rect 9767 33507 9825 33513
rect 7837 33439 7895 33445
rect 7837 33436 7849 33439
rect 7300 33408 7849 33436
rect 7837 33405 7849 33408
rect 7883 33405 7895 33439
rect 7837 33399 7895 33405
rect 7975 33439 8033 33445
rect 7975 33405 7987 33439
rect 8021 33436 8033 33439
rect 8757 33439 8815 33445
rect 8021 33408 8524 33436
rect 8021 33405 8033 33408
rect 7975 33399 8033 33405
rect 4580 33340 4936 33368
rect 4580 33328 4586 33340
rect 7374 33328 7380 33380
rect 7432 33368 7438 33380
rect 7561 33371 7619 33377
rect 7561 33368 7573 33371
rect 7432 33340 7573 33368
rect 7432 33328 7438 33340
rect 7561 33337 7573 33340
rect 7607 33337 7619 33371
rect 7561 33331 7619 33337
rect 8496 33368 8524 33408
rect 8757 33405 8769 33439
rect 8803 33436 8815 33439
rect 9324 33436 9352 33467
rect 8803 33408 9352 33436
rect 8803 33405 8815 33408
rect 8757 33399 8815 33405
rect 9416 33368 9444 33476
rect 9767 33473 9779 33507
rect 9813 33473 9825 33507
rect 9767 33467 9825 33473
rect 9858 33464 9864 33516
rect 9916 33504 9922 33516
rect 9916 33476 10640 33504
rect 9916 33464 9922 33476
rect 9493 33439 9551 33445
rect 9493 33405 9505 33439
rect 9539 33405 9551 33439
rect 10612 33436 10640 33476
rect 10686 33464 10692 33516
rect 10744 33504 10750 33516
rect 11793 33507 11851 33513
rect 11793 33504 11805 33507
rect 10744 33476 11805 33504
rect 10744 33464 10750 33476
rect 11793 33473 11805 33476
rect 11839 33473 11851 33507
rect 11793 33467 11851 33473
rect 11974 33464 11980 33516
rect 12032 33464 12038 33516
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 15439 33507 15497 33513
rect 15439 33504 15451 33507
rect 14056 33476 15451 33504
rect 14056 33464 14062 33476
rect 15439 33473 15451 33476
rect 15485 33504 15497 33507
rect 16574 33504 16580 33516
rect 15485 33476 16580 33504
rect 15485 33473 15497 33476
rect 15439 33467 15497 33473
rect 16574 33464 16580 33476
rect 16632 33464 16638 33516
rect 17126 33464 17132 33516
rect 17184 33464 17190 33516
rect 17236 33513 17264 33544
rect 17678 33532 17684 33544
rect 17736 33572 17742 33584
rect 19150 33572 19156 33584
rect 17736 33544 19156 33572
rect 17736 33532 17742 33544
rect 19150 33532 19156 33544
rect 19208 33572 19214 33584
rect 19208 33544 21864 33572
rect 19208 33532 19214 33544
rect 17221 33507 17279 33513
rect 17221 33473 17233 33507
rect 17267 33473 17279 33507
rect 17477 33507 17535 33513
rect 17477 33504 17489 33507
rect 17221 33467 17279 33473
rect 17328 33476 17489 33504
rect 11992 33436 12020 33464
rect 12526 33436 12532 33448
rect 10612 33408 12020 33436
rect 12084 33408 12532 33436
rect 9493 33399 9551 33405
rect 8496 33340 9444 33368
rect 5902 33260 5908 33312
rect 5960 33260 5966 33312
rect 6546 33260 6552 33312
rect 6604 33300 6610 33312
rect 8496 33300 8524 33340
rect 6604 33272 8524 33300
rect 9508 33300 9536 33399
rect 10428 33340 10824 33368
rect 9766 33300 9772 33312
rect 9508 33272 9772 33300
rect 6604 33260 6610 33272
rect 9766 33260 9772 33272
rect 9824 33300 9830 33312
rect 10428 33300 10456 33340
rect 10796 33312 10824 33340
rect 11698 33328 11704 33380
rect 11756 33368 11762 33380
rect 12084 33368 12112 33408
rect 12526 33396 12532 33408
rect 12584 33436 12590 33448
rect 12713 33439 12771 33445
rect 12713 33436 12725 33439
rect 12584 33408 12725 33436
rect 12584 33396 12590 33408
rect 12713 33405 12725 33408
rect 12759 33405 12771 33439
rect 12713 33399 12771 33405
rect 12802 33396 12808 33448
rect 12860 33445 12866 33448
rect 12860 33439 12888 33445
rect 12876 33405 12888 33439
rect 12860 33399 12888 33405
rect 12989 33439 13047 33445
rect 12989 33405 13001 33439
rect 13035 33436 13047 33439
rect 13630 33436 13636 33448
rect 13035 33408 13636 33436
rect 13035 33405 13047 33408
rect 12989 33399 13047 33405
rect 12860 33396 12866 33399
rect 13630 33396 13636 33408
rect 13688 33396 13694 33448
rect 15194 33396 15200 33448
rect 15252 33396 15258 33448
rect 17328 33436 17356 33476
rect 17477 33473 17489 33476
rect 17523 33504 17535 33507
rect 17770 33504 17776 33516
rect 17523 33476 17776 33504
rect 17523 33473 17535 33476
rect 17477 33467 17535 33473
rect 17770 33464 17776 33476
rect 17828 33464 17834 33516
rect 18230 33464 18236 33516
rect 18288 33464 18294 33516
rect 18598 33464 18604 33516
rect 18656 33504 18662 33516
rect 18693 33507 18751 33513
rect 18693 33504 18705 33507
rect 18656 33476 18705 33504
rect 18656 33464 18662 33476
rect 18693 33473 18705 33476
rect 18739 33504 18751 33507
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 18739 33476 19073 33504
rect 18739 33473 18751 33476
rect 18693 33467 18751 33473
rect 19061 33473 19073 33476
rect 19107 33473 19119 33507
rect 19061 33467 19119 33473
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33504 19303 33507
rect 19521 33507 19579 33513
rect 19291 33476 19380 33504
rect 19291 33473 19303 33476
rect 19245 33467 19303 33473
rect 17236 33408 17356 33436
rect 18248 33436 18276 33464
rect 18785 33439 18843 33445
rect 18785 33436 18797 33439
rect 18248 33408 18797 33436
rect 11756 33340 12112 33368
rect 12437 33371 12495 33377
rect 11756 33328 11762 33340
rect 12437 33337 12449 33371
rect 12483 33337 12495 33371
rect 12437 33331 12495 33337
rect 9824 33272 10456 33300
rect 9824 33260 9830 33272
rect 10502 33260 10508 33312
rect 10560 33260 10566 33312
rect 10778 33260 10784 33312
rect 10836 33260 10842 33312
rect 12452 33300 12480 33331
rect 13814 33328 13820 33380
rect 13872 33368 13878 33380
rect 15212 33368 15240 33396
rect 17236 33368 17264 33408
rect 18785 33405 18797 33408
rect 18831 33405 18843 33439
rect 18785 33399 18843 33405
rect 18969 33439 19027 33445
rect 18969 33405 18981 33439
rect 19015 33436 19027 33439
rect 19153 33439 19211 33445
rect 19153 33436 19165 33439
rect 19015 33408 19165 33436
rect 19015 33405 19027 33408
rect 18969 33399 19027 33405
rect 19153 33405 19165 33408
rect 19199 33405 19211 33439
rect 19153 33399 19211 33405
rect 19352 33377 19380 33476
rect 19521 33473 19533 33507
rect 19567 33473 19579 33507
rect 19521 33467 19579 33473
rect 13872 33340 15240 33368
rect 16132 33340 17264 33368
rect 18601 33371 18659 33377
rect 13872 33328 13878 33340
rect 12894 33300 12900 33312
rect 12452 33272 12900 33300
rect 12894 33260 12900 33272
rect 12952 33260 12958 33312
rect 14182 33260 14188 33312
rect 14240 33300 14246 33312
rect 16132 33300 16160 33340
rect 18601 33337 18613 33371
rect 18647 33368 18659 33371
rect 19337 33371 19395 33377
rect 18647 33340 19288 33368
rect 18647 33337 18659 33340
rect 18601 33331 18659 33337
rect 14240 33272 16160 33300
rect 14240 33260 14246 33272
rect 16206 33260 16212 33312
rect 16264 33260 16270 33312
rect 18874 33260 18880 33312
rect 18932 33260 18938 33312
rect 19260 33300 19288 33340
rect 19337 33337 19349 33371
rect 19383 33337 19395 33371
rect 19337 33331 19395 33337
rect 19536 33300 19564 33467
rect 20990 33464 20996 33516
rect 21048 33504 21054 33516
rect 21836 33513 21864 33544
rect 21637 33507 21695 33513
rect 21637 33504 21649 33507
rect 21048 33476 21649 33504
rect 21048 33464 21054 33476
rect 21637 33473 21649 33476
rect 21683 33473 21695 33507
rect 21637 33467 21695 33473
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 22077 33507 22135 33513
rect 22077 33504 22089 33507
rect 21821 33467 21879 33473
rect 21928 33476 22089 33504
rect 21652 33436 21680 33467
rect 21928 33436 21956 33476
rect 22077 33473 22089 33476
rect 22123 33473 22135 33507
rect 22664 33504 22692 33600
rect 23676 33572 23704 33600
rect 24121 33575 24179 33581
rect 24121 33572 24133 33575
rect 23676 33544 24133 33572
rect 24121 33541 24133 33544
rect 24167 33541 24179 33575
rect 24121 33535 24179 33541
rect 22664 33476 23060 33504
rect 22077 33467 22135 33473
rect 21652 33408 21956 33436
rect 23032 33368 23060 33476
rect 23106 33464 23112 33516
rect 23164 33504 23170 33516
rect 23293 33507 23351 33513
rect 23293 33504 23305 33507
rect 23164 33476 23305 33504
rect 23164 33464 23170 33476
rect 23293 33473 23305 33476
rect 23339 33504 23351 33507
rect 23661 33507 23719 33513
rect 23661 33504 23673 33507
rect 23339 33476 23673 33504
rect 23339 33473 23351 33476
rect 23293 33467 23351 33473
rect 23661 33473 23673 33476
rect 23707 33473 23719 33507
rect 23661 33467 23719 33473
rect 23845 33507 23903 33513
rect 23845 33473 23857 33507
rect 23891 33473 23903 33507
rect 23845 33467 23903 33473
rect 23569 33439 23627 33445
rect 23569 33405 23581 33439
rect 23615 33436 23627 33439
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 23615 33408 23765 33436
rect 23615 33405 23627 33408
rect 23569 33399 23627 33405
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 23860 33368 23888 33467
rect 23032 33340 23888 33368
rect 19260 33272 19564 33300
rect 21453 33303 21511 33309
rect 21453 33269 21465 33303
rect 21499 33300 21511 33303
rect 22186 33300 22192 33312
rect 21499 33272 22192 33300
rect 21499 33269 21511 33272
rect 21453 33263 21511 33269
rect 22186 33260 22192 33272
rect 22244 33260 22250 33312
rect 23382 33260 23388 33312
rect 23440 33260 23446 33312
rect 23474 33260 23480 33312
rect 23532 33260 23538 33312
rect 24394 33260 24400 33312
rect 24452 33260 24458 33312
rect 1104 33210 24840 33232
rect 1104 33158 3917 33210
rect 3969 33158 3981 33210
rect 4033 33158 4045 33210
rect 4097 33158 4109 33210
rect 4161 33158 4173 33210
rect 4225 33158 9851 33210
rect 9903 33158 9915 33210
rect 9967 33158 9979 33210
rect 10031 33158 10043 33210
rect 10095 33158 10107 33210
rect 10159 33158 15785 33210
rect 15837 33158 15849 33210
rect 15901 33158 15913 33210
rect 15965 33158 15977 33210
rect 16029 33158 16041 33210
rect 16093 33158 21719 33210
rect 21771 33158 21783 33210
rect 21835 33158 21847 33210
rect 21899 33158 21911 33210
rect 21963 33158 21975 33210
rect 22027 33158 24840 33210
rect 1104 33136 24840 33158
rect 1394 33056 1400 33108
rect 1452 33056 1458 33108
rect 2590 33056 2596 33108
rect 2648 33096 2654 33108
rect 3234 33096 3240 33108
rect 2648 33068 3240 33096
rect 2648 33056 2654 33068
rect 3234 33056 3240 33068
rect 3292 33056 3298 33108
rect 3329 33099 3387 33105
rect 3329 33065 3341 33099
rect 3375 33096 3387 33099
rect 3418 33096 3424 33108
rect 3375 33068 3424 33096
rect 3375 33065 3387 33068
rect 3329 33059 3387 33065
rect 3418 33056 3424 33068
rect 3476 33056 3482 33108
rect 3786 33056 3792 33108
rect 3844 33096 3850 33108
rect 4525 33099 4583 33105
rect 4525 33096 4537 33099
rect 3844 33068 4537 33096
rect 3844 33056 3850 33068
rect 4525 33065 4537 33068
rect 4571 33065 4583 33099
rect 4525 33059 4583 33065
rect 8110 33056 8116 33108
rect 8168 33096 8174 33108
rect 8205 33099 8263 33105
rect 8205 33096 8217 33099
rect 8168 33068 8217 33096
rect 8168 33056 8174 33068
rect 8205 33065 8217 33068
rect 8251 33065 8263 33099
rect 8205 33059 8263 33065
rect 9674 33056 9680 33108
rect 9732 33096 9738 33108
rect 9732 33068 12848 33096
rect 9732 33056 9738 33068
rect 1412 32960 1440 33056
rect 4890 33028 4896 33040
rect 3160 33000 4896 33028
rect 2314 32960 2320 32972
rect 1412 32932 2320 32960
rect 2314 32920 2320 32932
rect 2372 32920 2378 32972
rect 3160 32904 3188 33000
rect 3326 32920 3332 32972
rect 3384 32960 3390 32972
rect 3988 32969 4016 33000
rect 4890 32988 4896 33000
rect 4948 32988 4954 33040
rect 10502 32988 10508 33040
rect 10560 33028 10566 33040
rect 10597 33031 10655 33037
rect 10597 33028 10609 33031
rect 10560 33000 10609 33028
rect 10560 32988 10566 33000
rect 10597 32997 10609 33000
rect 10643 32997 10655 33031
rect 10597 32991 10655 32997
rect 11606 32988 11612 33040
rect 11664 32988 11670 33040
rect 12820 33028 12848 33068
rect 12894 33056 12900 33108
rect 12952 33056 12958 33108
rect 15933 33099 15991 33105
rect 15933 33065 15945 33099
rect 15979 33096 15991 33099
rect 16114 33096 16120 33108
rect 15979 33068 16120 33096
rect 15979 33065 15991 33068
rect 15933 33059 15991 33065
rect 16114 33056 16120 33068
rect 16172 33056 16178 33108
rect 16574 33056 16580 33108
rect 16632 33096 16638 33108
rect 16632 33068 18552 33096
rect 16632 33056 16638 33068
rect 13998 33028 14004 33040
rect 12820 33000 14004 33028
rect 13998 32988 14004 33000
rect 14056 32988 14062 33040
rect 14737 33031 14795 33037
rect 14737 32997 14749 33031
rect 14783 33028 14795 33031
rect 14826 33028 14832 33040
rect 14783 33000 14832 33028
rect 14783 32997 14795 33000
rect 14737 32991 14795 32997
rect 14826 32988 14832 33000
rect 14884 32988 14890 33040
rect 18524 33028 18552 33068
rect 18598 33056 18604 33108
rect 18656 33056 18662 33108
rect 20622 33096 20628 33108
rect 19306 33068 20628 33096
rect 19306 33028 19334 33068
rect 20622 33056 20628 33068
rect 20680 33056 20686 33108
rect 22281 33099 22339 33105
rect 22281 33065 22293 33099
rect 22327 33096 22339 33099
rect 23382 33096 23388 33108
rect 22327 33068 23388 33096
rect 22327 33065 22339 33068
rect 22281 33059 22339 33065
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 23492 33068 25728 33096
rect 18524 33000 19334 33028
rect 21913 33031 21971 33037
rect 21913 32997 21925 33031
rect 21959 33028 21971 33031
rect 21959 33000 23060 33028
rect 21959 32997 21971 33000
rect 21913 32991 21971 32997
rect 3973 32963 4031 32969
rect 3384 32932 3924 32960
rect 3384 32920 3390 32932
rect 1394 32852 1400 32904
rect 1452 32852 1458 32904
rect 2591 32895 2649 32901
rect 2591 32861 2603 32895
rect 2637 32861 2649 32895
rect 2591 32855 2649 32861
rect 1670 32784 1676 32836
rect 1728 32784 1734 32836
rect 2606 32824 2634 32855
rect 3142 32852 3148 32904
rect 3200 32852 3206 32904
rect 3789 32895 3847 32901
rect 3789 32861 3801 32895
rect 3835 32861 3847 32895
rect 3896 32892 3924 32932
rect 3973 32929 3985 32963
rect 4019 32929 4031 32963
rect 3973 32923 4031 32929
rect 5534 32920 5540 32972
rect 5592 32920 5598 32972
rect 6178 32920 6184 32972
rect 6236 32960 6242 32972
rect 7193 32963 7251 32969
rect 7193 32960 7205 32963
rect 6236 32932 7205 32960
rect 6236 32920 6242 32932
rect 7193 32929 7205 32932
rect 7239 32929 7251 32963
rect 7193 32923 7251 32929
rect 9030 32920 9036 32972
rect 9088 32960 9094 32972
rect 10137 32963 10195 32969
rect 10137 32960 10149 32963
rect 9088 32932 10149 32960
rect 9088 32920 9094 32932
rect 10137 32929 10149 32932
rect 10183 32960 10195 32963
rect 10686 32960 10692 32972
rect 10183 32932 10692 32960
rect 10183 32929 10195 32932
rect 10137 32923 10195 32929
rect 10686 32920 10692 32932
rect 10744 32920 10750 32972
rect 11011 32963 11069 32969
rect 11011 32929 11023 32963
rect 11057 32960 11069 32963
rect 11330 32960 11336 32972
rect 11057 32932 11336 32960
rect 11057 32929 11069 32932
rect 11011 32923 11069 32929
rect 11330 32920 11336 32932
rect 11388 32920 11394 32972
rect 11624 32960 11652 32988
rect 11624 32932 11836 32960
rect 5261 32895 5319 32901
rect 5261 32892 5273 32895
rect 3896 32864 5273 32892
rect 3789 32855 3847 32861
rect 5261 32861 5273 32864
rect 5307 32861 5319 32895
rect 5261 32855 5319 32861
rect 5353 32895 5411 32901
rect 5353 32861 5365 32895
rect 5399 32892 5411 32895
rect 5902 32892 5908 32904
rect 5399 32864 5908 32892
rect 5399 32861 5411 32864
rect 5353 32855 5411 32861
rect 3418 32824 3424 32836
rect 2606 32796 3424 32824
rect 3418 32784 3424 32796
rect 3476 32784 3482 32836
rect 1210 32716 1216 32768
rect 1268 32756 1274 32768
rect 3804 32756 3832 32855
rect 5902 32852 5908 32864
rect 5960 32852 5966 32904
rect 6914 32852 6920 32904
rect 6972 32892 6978 32904
rect 8018 32892 8024 32904
rect 6972 32865 8024 32892
rect 6972 32864 7463 32865
rect 6972 32852 6978 32864
rect 4338 32784 4344 32836
rect 4396 32824 4402 32836
rect 5721 32827 5779 32833
rect 4396 32796 5212 32824
rect 4396 32784 4402 32796
rect 1268 32728 3832 32756
rect 1268 32716 1274 32728
rect 4706 32716 4712 32768
rect 4764 32756 4770 32768
rect 4985 32759 5043 32765
rect 4985 32756 4997 32759
rect 4764 32728 4997 32756
rect 4764 32716 4770 32728
rect 4985 32725 4997 32728
rect 5031 32725 5043 32759
rect 5184 32756 5212 32796
rect 5721 32793 5733 32827
rect 5767 32793 5779 32827
rect 7006 32824 7012 32836
rect 5721 32787 5779 32793
rect 5920 32796 7012 32824
rect 5350 32756 5356 32768
rect 5184 32728 5356 32756
rect 4985 32719 5043 32725
rect 5350 32716 5356 32728
rect 5408 32756 5414 32768
rect 5736 32756 5764 32787
rect 5920 32768 5948 32796
rect 7006 32784 7012 32796
rect 7064 32784 7070 32836
rect 7451 32831 7463 32864
rect 7497 32864 8024 32865
rect 7497 32834 7512 32864
rect 8018 32852 8024 32864
rect 8076 32852 8082 32904
rect 8754 32852 8760 32904
rect 8812 32892 8818 32904
rect 9214 32892 9220 32904
rect 8812 32864 9220 32892
rect 8812 32852 8818 32864
rect 9214 32852 9220 32864
rect 9272 32852 9278 32904
rect 9953 32895 10011 32901
rect 9953 32861 9965 32895
rect 9999 32861 10011 32895
rect 9953 32855 10011 32861
rect 7497 32831 7509 32834
rect 7451 32825 7509 32831
rect 5408 32728 5764 32756
rect 5408 32716 5414 32728
rect 5902 32716 5908 32768
rect 5960 32716 5966 32768
rect 6086 32716 6092 32768
rect 6144 32716 6150 32768
rect 6270 32716 6276 32768
rect 6328 32716 6334 32768
rect 7024 32756 7052 32784
rect 7742 32756 7748 32768
rect 7024 32728 7748 32756
rect 7742 32716 7748 32728
rect 7800 32716 7806 32768
rect 9968 32756 9996 32855
rect 10870 32852 10876 32904
rect 10928 32852 10934 32904
rect 11146 32852 11152 32904
rect 11204 32852 11210 32904
rect 11808 32892 11836 32932
rect 11882 32920 11888 32972
rect 11940 32920 11946 32972
rect 13906 32920 13912 32972
rect 13964 32960 13970 32972
rect 15151 32963 15209 32969
rect 15151 32960 15163 32963
rect 13964 32932 15163 32960
rect 13964 32920 13970 32932
rect 15151 32929 15163 32932
rect 15197 32960 15209 32963
rect 15197 32932 16160 32960
rect 15197 32929 15209 32932
rect 15151 32923 15209 32929
rect 16132 32904 16160 32932
rect 17586 32920 17592 32972
rect 17644 32920 17650 32972
rect 21266 32920 21272 32972
rect 21324 32960 21330 32972
rect 22646 32960 22652 32972
rect 21324 32932 22652 32960
rect 21324 32920 21330 32932
rect 22646 32920 22652 32932
rect 22704 32920 22710 32972
rect 12158 32901 12164 32904
rect 12127 32895 12164 32901
rect 12127 32892 12139 32895
rect 11808 32864 12139 32892
rect 12127 32861 12139 32864
rect 12127 32855 12164 32861
rect 12158 32852 12164 32855
rect 12216 32852 12222 32904
rect 12526 32852 12532 32904
rect 12584 32892 12590 32904
rect 14093 32895 14151 32901
rect 14093 32892 14105 32895
rect 12584 32864 14105 32892
rect 12584 32852 12590 32864
rect 14093 32861 14105 32864
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 14277 32895 14335 32901
rect 14277 32861 14289 32895
rect 14323 32861 14335 32895
rect 14277 32855 14335 32861
rect 11793 32827 11851 32833
rect 11793 32793 11805 32827
rect 11839 32824 11851 32827
rect 14182 32824 14188 32836
rect 11839 32796 14188 32824
rect 11839 32793 11851 32796
rect 11793 32787 11851 32793
rect 14182 32784 14188 32796
rect 14240 32784 14246 32836
rect 10410 32756 10416 32768
rect 9968 32728 10416 32756
rect 10410 32716 10416 32728
rect 10468 32756 10474 32768
rect 12802 32756 12808 32768
rect 10468 32728 12808 32756
rect 10468 32716 10474 32728
rect 12802 32716 12808 32728
rect 12860 32716 12866 32768
rect 14292 32756 14320 32855
rect 15010 32852 15016 32904
rect 15068 32852 15074 32904
rect 15286 32852 15292 32904
rect 15344 32852 15350 32904
rect 16022 32852 16028 32904
rect 16080 32852 16086 32904
rect 16114 32852 16120 32904
rect 16172 32852 16178 32904
rect 17402 32852 17408 32904
rect 17460 32892 17466 32904
rect 17770 32892 17776 32904
rect 17460 32864 17776 32892
rect 17460 32852 17466 32864
rect 17770 32852 17776 32864
rect 17828 32901 17834 32904
rect 22094 32901 22100 32904
rect 17828 32895 17889 32901
rect 17828 32861 17843 32895
rect 17877 32861 17889 32895
rect 22089 32892 22100 32901
rect 17828 32855 17889 32861
rect 19306 32864 22100 32892
rect 17828 32852 17834 32855
rect 16040 32824 16068 32852
rect 19306 32824 19334 32864
rect 22089 32855 22100 32864
rect 22094 32852 22100 32855
rect 22152 32852 22158 32904
rect 22186 32852 22192 32904
rect 22244 32894 22250 32904
rect 23032 32901 23060 33000
rect 23017 32895 23075 32901
rect 22244 32866 22287 32894
rect 22244 32852 22250 32866
rect 23017 32861 23029 32895
rect 23063 32861 23075 32895
rect 23492 32892 23520 33068
rect 23661 33031 23719 33037
rect 23661 32997 23673 33031
rect 23707 32997 23719 33031
rect 23661 32991 23719 32997
rect 23017 32855 23075 32861
rect 23124 32864 23520 32892
rect 23569 32895 23627 32901
rect 23124 32824 23152 32864
rect 23569 32861 23581 32895
rect 23615 32892 23627 32895
rect 23676 32892 23704 32991
rect 25700 32972 25728 33068
rect 25682 32920 25688 32972
rect 25740 32920 25746 32972
rect 23615 32864 23704 32892
rect 23615 32861 23627 32864
rect 23569 32855 23627 32861
rect 23750 32852 23756 32904
rect 23808 32852 23814 32904
rect 23845 32895 23903 32901
rect 23845 32861 23857 32895
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 16040 32796 19334 32824
rect 22756 32796 23152 32824
rect 15194 32756 15200 32768
rect 14292 32728 15200 32756
rect 15194 32716 15200 32728
rect 15252 32716 15258 32768
rect 15378 32716 15384 32768
rect 15436 32756 15442 32768
rect 22756 32756 22784 32796
rect 23290 32784 23296 32836
rect 23348 32784 23354 32836
rect 15436 32728 22784 32756
rect 22833 32759 22891 32765
rect 15436 32716 15442 32728
rect 22833 32725 22845 32759
rect 22879 32756 22891 32759
rect 23308 32756 23336 32784
rect 22879 32728 23336 32756
rect 23385 32759 23443 32765
rect 22879 32725 22891 32728
rect 22833 32719 22891 32725
rect 23385 32725 23397 32759
rect 23431 32756 23443 32759
rect 23768 32756 23796 32852
rect 23860 32824 23888 32855
rect 23934 32852 23940 32904
rect 23992 32852 23998 32904
rect 25038 32824 25044 32836
rect 23860 32796 25044 32824
rect 25038 32784 25044 32796
rect 25096 32784 25102 32836
rect 23431 32728 23796 32756
rect 24121 32759 24179 32765
rect 23431 32725 23443 32728
rect 23385 32719 23443 32725
rect 24121 32725 24133 32759
rect 24167 32756 24179 32759
rect 25222 32756 25228 32768
rect 24167 32728 25228 32756
rect 24167 32725 24179 32728
rect 24121 32719 24179 32725
rect 25222 32716 25228 32728
rect 25280 32716 25286 32768
rect 1104 32666 25000 32688
rect 1104 32614 6884 32666
rect 6936 32614 6948 32666
rect 7000 32614 7012 32666
rect 7064 32614 7076 32666
rect 7128 32614 7140 32666
rect 7192 32614 12818 32666
rect 12870 32614 12882 32666
rect 12934 32614 12946 32666
rect 12998 32614 13010 32666
rect 13062 32614 13074 32666
rect 13126 32614 18752 32666
rect 18804 32614 18816 32666
rect 18868 32614 18880 32666
rect 18932 32614 18944 32666
rect 18996 32614 19008 32666
rect 19060 32614 24686 32666
rect 24738 32614 24750 32666
rect 24802 32614 24814 32666
rect 24866 32614 24878 32666
rect 24930 32614 24942 32666
rect 24994 32614 25000 32666
rect 1104 32592 25000 32614
rect 1118 32512 1124 32564
rect 1176 32552 1182 32564
rect 1176 32524 3096 32552
rect 1176 32512 1182 32524
rect 3068 32484 3096 32524
rect 4614 32512 4620 32564
rect 4672 32552 4678 32564
rect 4982 32552 4988 32564
rect 4672 32524 4988 32552
rect 4672 32512 4678 32524
rect 4982 32512 4988 32524
rect 5040 32552 5046 32564
rect 6086 32552 6092 32564
rect 5040 32524 6092 32552
rect 5040 32512 5046 32524
rect 6086 32512 6092 32524
rect 6144 32512 6150 32564
rect 6270 32512 6276 32564
rect 6328 32512 6334 32564
rect 7558 32512 7564 32564
rect 7616 32552 7622 32564
rect 7742 32552 7748 32564
rect 7616 32524 7748 32552
rect 7616 32512 7622 32524
rect 7742 32512 7748 32524
rect 7800 32552 7806 32564
rect 11057 32555 11115 32561
rect 7800 32524 10330 32552
rect 7800 32512 7806 32524
rect 3881 32487 3939 32493
rect 3881 32484 3893 32487
rect 3068 32456 3893 32484
rect 3881 32453 3893 32456
rect 3927 32453 3939 32487
rect 3881 32447 3939 32453
rect 5718 32444 5724 32496
rect 5776 32444 5782 32496
rect 6288 32484 6316 32512
rect 10134 32484 10140 32496
rect 6288 32456 10140 32484
rect 10134 32444 10140 32456
rect 10192 32444 10198 32496
rect 10302 32455 10330 32524
rect 11057 32521 11069 32555
rect 11103 32552 11115 32555
rect 11146 32552 11152 32564
rect 11103 32524 11152 32552
rect 11103 32521 11115 32524
rect 11057 32515 11115 32521
rect 11146 32512 11152 32524
rect 11204 32512 11210 32564
rect 13906 32512 13912 32564
rect 13964 32552 13970 32564
rect 14093 32555 14151 32561
rect 14093 32552 14105 32555
rect 13964 32524 14105 32552
rect 13964 32512 13970 32524
rect 14093 32521 14105 32524
rect 14139 32521 14151 32555
rect 14093 32515 14151 32521
rect 15194 32512 15200 32564
rect 15252 32512 15258 32564
rect 15378 32512 15384 32564
rect 15436 32512 15442 32564
rect 16758 32512 16764 32564
rect 16816 32552 16822 32564
rect 22649 32555 22707 32561
rect 16816 32524 22048 32552
rect 16816 32512 16822 32524
rect 10302 32449 10361 32455
rect 2406 32376 2412 32428
rect 2464 32425 2470 32428
rect 2464 32419 2492 32425
rect 2480 32385 2492 32419
rect 2464 32379 2492 32385
rect 3329 32419 3387 32425
rect 3329 32385 3341 32419
rect 3375 32385 3387 32419
rect 5736 32416 5764 32444
rect 6086 32416 6092 32428
rect 5736 32388 6092 32416
rect 3329 32379 3387 32385
rect 2464 32376 2470 32379
rect 1397 32351 1455 32357
rect 1397 32317 1409 32351
rect 1443 32348 1455 32351
rect 1486 32348 1492 32360
rect 1443 32320 1492 32348
rect 1443 32317 1455 32320
rect 1397 32311 1455 32317
rect 1486 32308 1492 32320
rect 1544 32308 1550 32360
rect 1578 32308 1584 32360
rect 1636 32308 1642 32360
rect 2041 32351 2099 32357
rect 2041 32317 2053 32351
rect 2087 32348 2099 32351
rect 2130 32348 2136 32360
rect 2087 32320 2136 32348
rect 2087 32317 2099 32320
rect 2041 32311 2099 32317
rect 2130 32308 2136 32320
rect 2188 32308 2194 32360
rect 2314 32308 2320 32360
rect 2372 32308 2378 32360
rect 2590 32308 2596 32360
rect 2648 32308 2654 32360
rect 2958 32308 2964 32360
rect 3016 32348 3022 32360
rect 3237 32351 3295 32357
rect 3237 32348 3249 32351
rect 3016 32320 3249 32348
rect 3016 32308 3022 32320
rect 3237 32317 3249 32320
rect 3283 32317 3295 32351
rect 3237 32311 3295 32317
rect 1210 32172 1216 32224
rect 1268 32212 1274 32224
rect 3344 32212 3372 32379
rect 6086 32376 6092 32388
rect 6144 32376 6150 32428
rect 8295 32419 8353 32425
rect 8295 32385 8307 32419
rect 8341 32416 8353 32419
rect 8341 32388 8708 32416
rect 8341 32385 8353 32388
rect 8295 32379 8353 32385
rect 3418 32308 3424 32360
rect 3476 32348 3482 32360
rect 3605 32351 3663 32357
rect 3605 32348 3617 32351
rect 3476 32320 3617 32348
rect 3476 32308 3482 32320
rect 3605 32317 3617 32320
rect 3651 32348 3663 32351
rect 3786 32348 3792 32360
rect 3651 32320 3792 32348
rect 3651 32317 3663 32320
rect 3605 32311 3663 32317
rect 3786 32308 3792 32320
rect 3844 32348 3850 32360
rect 4246 32348 4252 32360
rect 3844 32320 4252 32348
rect 3844 32308 3850 32320
rect 4246 32308 4252 32320
rect 4304 32308 4310 32360
rect 4614 32308 4620 32360
rect 4672 32308 4678 32360
rect 8021 32351 8079 32357
rect 8021 32317 8033 32351
rect 8067 32317 8079 32351
rect 8680 32348 8708 32388
rect 8754 32376 8760 32428
rect 8812 32416 8818 32428
rect 9766 32416 9772 32428
rect 8812 32388 9772 32416
rect 8812 32376 8818 32388
rect 9766 32376 9772 32388
rect 9824 32416 9830 32428
rect 10045 32419 10103 32425
rect 10045 32416 10057 32419
rect 9824 32388 10057 32416
rect 9824 32376 9830 32388
rect 10045 32385 10057 32388
rect 10091 32385 10103 32419
rect 10302 32418 10315 32449
rect 10303 32415 10315 32418
rect 10349 32415 10361 32449
rect 10594 32444 10600 32496
rect 10652 32484 10658 32496
rect 13722 32484 13728 32496
rect 10652 32456 13728 32484
rect 10652 32444 10658 32456
rect 13722 32444 13728 32456
rect 13780 32484 13786 32496
rect 13780 32456 14136 32484
rect 13780 32444 13786 32456
rect 10303 32409 10361 32415
rect 10045 32379 10103 32385
rect 9306 32348 9312 32360
rect 8680 32320 9312 32348
rect 8021 32311 8079 32317
rect 4632 32280 4660 32308
rect 5626 32280 5632 32292
rect 4632 32252 5632 32280
rect 5626 32240 5632 32252
rect 5684 32240 5690 32292
rect 1268 32184 3372 32212
rect 1268 32172 1274 32184
rect 5350 32172 5356 32224
rect 5408 32212 5414 32224
rect 6730 32212 6736 32224
rect 5408 32184 6736 32212
rect 5408 32172 5414 32184
rect 6730 32172 6736 32184
rect 6788 32172 6794 32224
rect 8036 32212 8064 32311
rect 9306 32308 9312 32320
rect 9364 32308 9370 32360
rect 8386 32212 8392 32224
rect 8036 32184 8392 32212
rect 8386 32172 8392 32184
rect 8444 32172 8450 32224
rect 9030 32172 9036 32224
rect 9088 32172 9094 32224
rect 10060 32212 10088 32379
rect 10870 32376 10876 32428
rect 10928 32416 10934 32428
rect 11974 32416 11980 32428
rect 10928 32388 11980 32416
rect 10928 32376 10934 32388
rect 11974 32376 11980 32388
rect 12032 32376 12038 32428
rect 14108 32416 14136 32456
rect 14182 32444 14188 32496
rect 14240 32484 14246 32496
rect 14328 32487 14386 32493
rect 14328 32484 14340 32487
rect 14240 32456 14340 32484
rect 14240 32444 14246 32456
rect 14328 32453 14340 32456
rect 14374 32453 14386 32487
rect 14328 32447 14386 32453
rect 14458 32444 14464 32496
rect 14516 32444 14522 32496
rect 16574 32484 16580 32496
rect 14844 32456 16580 32484
rect 14844 32425 14872 32456
rect 16574 32444 16580 32456
rect 16632 32444 16638 32496
rect 19420 32487 19478 32493
rect 19420 32453 19432 32487
rect 19466 32484 19478 32487
rect 19518 32484 19524 32496
rect 19466 32456 19524 32484
rect 19466 32453 19478 32456
rect 19420 32447 19478 32453
rect 19518 32444 19524 32456
rect 19576 32444 19582 32496
rect 14829 32419 14887 32425
rect 14829 32416 14841 32419
rect 14108 32388 14841 32416
rect 14829 32385 14841 32388
rect 14875 32385 14887 32419
rect 14829 32379 14887 32385
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32416 19211 32419
rect 19242 32416 19248 32428
rect 19199 32388 19248 32416
rect 19199 32385 19211 32388
rect 19153 32379 19211 32385
rect 19242 32376 19248 32388
rect 19300 32376 19306 32428
rect 22020 32425 22048 32524
rect 22649 32521 22661 32555
rect 22695 32552 22707 32555
rect 23661 32555 23719 32561
rect 22695 32524 23612 32552
rect 22695 32521 22707 32524
rect 22649 32515 22707 32521
rect 23584 32425 23612 32524
rect 23661 32521 23673 32555
rect 23707 32552 23719 32555
rect 23934 32552 23940 32564
rect 23707 32524 23940 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 23934 32512 23940 32524
rect 23992 32512 23998 32564
rect 22005 32419 22063 32425
rect 22005 32385 22017 32419
rect 22051 32385 22063 32419
rect 22005 32379 22063 32385
rect 22557 32419 22615 32425
rect 22557 32385 22569 32419
rect 22603 32385 22615 32419
rect 22557 32379 22615 32385
rect 22833 32419 22891 32425
rect 22833 32385 22845 32419
rect 22879 32385 22891 32419
rect 23293 32419 23351 32425
rect 23293 32416 23305 32419
rect 22833 32379 22891 32385
rect 22940 32388 23305 32416
rect 15108 32360 15160 32366
rect 11330 32308 11336 32360
rect 11388 32348 11394 32360
rect 11514 32348 11520 32360
rect 11388 32320 11520 32348
rect 11388 32308 11394 32320
rect 11514 32308 11520 32320
rect 11572 32308 11578 32360
rect 15194 32308 15200 32360
rect 15252 32348 15258 32360
rect 15470 32348 15476 32360
rect 15252 32320 15476 32348
rect 15252 32308 15258 32320
rect 15470 32308 15476 32320
rect 15528 32308 15534 32360
rect 22572 32348 22600 32379
rect 22066 32320 22600 32348
rect 15108 32302 15160 32308
rect 21821 32283 21879 32289
rect 20088 32252 20668 32280
rect 11146 32212 11152 32224
rect 10060 32184 11152 32212
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 15562 32172 15568 32224
rect 15620 32212 15626 32224
rect 16298 32212 16304 32224
rect 15620 32184 16304 32212
rect 15620 32172 15626 32184
rect 16298 32172 16304 32184
rect 16356 32212 16362 32224
rect 19150 32212 19156 32224
rect 16356 32184 19156 32212
rect 16356 32172 16362 32184
rect 19150 32172 19156 32184
rect 19208 32212 19214 32224
rect 20088 32212 20116 32252
rect 19208 32184 20116 32212
rect 19208 32172 19214 32184
rect 20530 32172 20536 32224
rect 20588 32172 20594 32224
rect 20640 32212 20668 32252
rect 21821 32249 21833 32283
rect 21867 32280 21879 32283
rect 22066 32280 22094 32320
rect 22848 32280 22876 32379
rect 21867 32252 22094 32280
rect 22296 32252 22876 32280
rect 21867 32249 21879 32252
rect 21821 32243 21879 32249
rect 22296 32212 22324 32252
rect 20640 32184 22324 32212
rect 22373 32215 22431 32221
rect 22373 32181 22385 32215
rect 22419 32212 22431 32215
rect 22940 32212 22968 32388
rect 23293 32385 23305 32388
rect 23339 32385 23351 32419
rect 23293 32379 23351 32385
rect 23569 32419 23627 32425
rect 23569 32385 23581 32419
rect 23615 32385 23627 32419
rect 23569 32379 23627 32385
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 23860 32348 23888 32379
rect 24118 32376 24124 32428
rect 24176 32376 24182 32428
rect 24213 32419 24271 32425
rect 24213 32385 24225 32419
rect 24259 32385 24271 32419
rect 24213 32379 24271 32385
rect 23400 32320 23888 32348
rect 23400 32289 23428 32320
rect 23385 32283 23443 32289
rect 23385 32249 23397 32283
rect 23431 32249 23443 32283
rect 24228 32280 24256 32379
rect 23385 32243 23443 32249
rect 23860 32252 24256 32280
rect 22419 32184 22968 32212
rect 23109 32215 23167 32221
rect 22419 32181 22431 32184
rect 22373 32175 22431 32181
rect 23109 32181 23121 32215
rect 23155 32212 23167 32215
rect 23860 32212 23888 32252
rect 23155 32184 23888 32212
rect 23937 32215 23995 32221
rect 23155 32181 23167 32184
rect 23109 32175 23167 32181
rect 23937 32181 23949 32215
rect 23983 32212 23995 32215
rect 24026 32212 24032 32224
rect 23983 32184 24032 32212
rect 23983 32181 23995 32184
rect 23937 32175 23995 32181
rect 24026 32172 24032 32184
rect 24084 32172 24090 32224
rect 24394 32172 24400 32224
rect 24452 32172 24458 32224
rect 1104 32122 24840 32144
rect 1104 32070 3917 32122
rect 3969 32070 3981 32122
rect 4033 32070 4045 32122
rect 4097 32070 4109 32122
rect 4161 32070 4173 32122
rect 4225 32070 9851 32122
rect 9903 32070 9915 32122
rect 9967 32070 9979 32122
rect 10031 32070 10043 32122
rect 10095 32070 10107 32122
rect 10159 32070 15785 32122
rect 15837 32070 15849 32122
rect 15901 32070 15913 32122
rect 15965 32070 15977 32122
rect 16029 32070 16041 32122
rect 16093 32070 21719 32122
rect 21771 32070 21783 32122
rect 21835 32070 21847 32122
rect 21899 32070 21911 32122
rect 21963 32070 21975 32122
rect 22027 32070 24840 32122
rect 1104 32048 24840 32070
rect 2409 32011 2467 32017
rect 2409 31977 2421 32011
rect 2455 32008 2467 32011
rect 2590 32008 2596 32020
rect 2455 31980 2596 32008
rect 2455 31977 2467 31980
rect 2409 31971 2467 31977
rect 2590 31968 2596 31980
rect 2648 31968 2654 32020
rect 4709 32011 4767 32017
rect 4709 31977 4721 32011
rect 4755 32008 4767 32011
rect 5166 32008 5172 32020
rect 4755 31980 5172 32008
rect 4755 31977 4767 31980
rect 4709 31971 4767 31977
rect 5166 31968 5172 31980
rect 5224 31968 5230 32020
rect 9582 32008 9588 32020
rect 5920 31980 9588 32008
rect 5920 31940 5948 31980
rect 9582 31968 9588 31980
rect 9640 31968 9646 32020
rect 9692 31980 11744 32008
rect 3068 31912 5948 31940
rect 842 31832 848 31884
rect 900 31832 906 31884
rect 2406 31832 2412 31884
rect 2464 31872 2470 31884
rect 2958 31872 2964 31884
rect 2464 31844 2964 31872
rect 2464 31832 2470 31844
rect 2958 31832 2964 31844
rect 3016 31832 3022 31884
rect 3068 31881 3096 31912
rect 6730 31900 6736 31952
rect 6788 31940 6794 31952
rect 9692 31940 9720 31980
rect 6788 31912 9720 31940
rect 6788 31900 6794 31912
rect 3053 31875 3111 31881
rect 3053 31841 3065 31875
rect 3099 31841 3111 31875
rect 3053 31835 3111 31841
rect 3160 31844 5580 31872
rect 860 31804 888 31832
rect 1397 31807 1455 31813
rect 1397 31804 1409 31807
rect 860 31776 1409 31804
rect 1320 31680 1348 31776
rect 1397 31773 1409 31776
rect 1443 31773 1455 31807
rect 1397 31767 1455 31773
rect 1671 31807 1729 31813
rect 1671 31773 1683 31807
rect 1717 31804 1729 31807
rect 2682 31804 2688 31816
rect 1717 31776 2688 31804
rect 1717 31773 1729 31776
rect 1671 31767 1729 31773
rect 2682 31764 2688 31776
rect 2740 31764 2746 31816
rect 2774 31764 2780 31816
rect 2832 31764 2838 31816
rect 3160 31804 3188 31844
rect 5552 31816 5580 31844
rect 7650 31832 7656 31884
rect 7708 31872 7714 31884
rect 8110 31872 8116 31884
rect 7708 31844 8116 31872
rect 7708 31832 7714 31844
rect 8110 31832 8116 31844
rect 8168 31832 8174 31884
rect 8386 31832 8392 31884
rect 8444 31872 8450 31884
rect 9122 31872 9128 31884
rect 8444 31844 9128 31872
rect 8444 31832 8450 31844
rect 9122 31832 9128 31844
rect 9180 31832 9186 31884
rect 11716 31872 11744 31980
rect 11882 31968 11888 32020
rect 11940 32008 11946 32020
rect 14458 32008 14464 32020
rect 11940 31980 14464 32008
rect 11940 31968 11946 31980
rect 14458 31968 14464 31980
rect 14516 31968 14522 32020
rect 15102 31968 15108 32020
rect 15160 31968 15166 32020
rect 15286 31968 15292 32020
rect 15344 32008 15350 32020
rect 15562 32008 15568 32020
rect 15344 31980 15568 32008
rect 15344 31968 15350 31980
rect 15562 31968 15568 31980
rect 15620 31968 15626 32020
rect 16758 32008 16764 32020
rect 16316 31980 16764 32008
rect 16206 31900 16212 31952
rect 16264 31900 16270 31952
rect 11716 31844 13216 31872
rect 2884 31776 3188 31804
rect 2222 31696 2228 31748
rect 2280 31696 2286 31748
rect 2406 31696 2412 31748
rect 2464 31736 2470 31748
rect 2884 31736 2912 31776
rect 3786 31764 3792 31816
rect 3844 31764 3850 31816
rect 4890 31764 4896 31816
rect 4948 31764 4954 31816
rect 5534 31764 5540 31816
rect 5592 31764 5598 31816
rect 5813 31807 5871 31813
rect 5813 31773 5825 31807
rect 5859 31773 5871 31807
rect 6086 31804 6092 31816
rect 6047 31776 6092 31804
rect 5813 31767 5871 31773
rect 2464 31708 2912 31736
rect 4065 31739 4123 31745
rect 2464 31696 2470 31708
rect 4065 31705 4077 31739
rect 4111 31705 4123 31739
rect 5828 31736 5856 31767
rect 6086 31764 6092 31776
rect 6144 31764 6150 31816
rect 6178 31764 6184 31816
rect 6236 31804 6242 31816
rect 6454 31804 6460 31816
rect 6236 31776 6460 31804
rect 6236 31764 6242 31776
rect 6454 31764 6460 31776
rect 6512 31764 6518 31816
rect 8478 31764 8484 31816
rect 8536 31804 8542 31816
rect 10870 31804 10876 31816
rect 8536 31776 10876 31804
rect 8536 31764 8542 31776
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 11057 31807 11115 31813
rect 11057 31773 11069 31807
rect 11103 31773 11115 31807
rect 11057 31767 11115 31773
rect 11331 31807 11389 31813
rect 11331 31773 11343 31807
rect 11377 31804 11389 31807
rect 11716 31804 11744 31844
rect 11377 31776 11744 31804
rect 11377 31773 11389 31776
rect 11331 31767 11389 31773
rect 6270 31736 6276 31748
rect 5828 31708 6276 31736
rect 4065 31699 4123 31705
rect 1302 31628 1308 31680
rect 1360 31628 1366 31680
rect 2240 31668 2268 31696
rect 2958 31668 2964 31680
rect 2240 31640 2964 31668
rect 2958 31628 2964 31640
rect 3016 31668 3022 31680
rect 4080 31668 4108 31699
rect 6270 31696 6276 31708
rect 6328 31696 6334 31748
rect 7466 31696 7472 31748
rect 7524 31736 7530 31748
rect 11072 31736 11100 31767
rect 12342 31764 12348 31816
rect 12400 31764 12406 31816
rect 12526 31764 12532 31816
rect 12584 31804 12590 31816
rect 13081 31807 13139 31813
rect 13081 31804 13093 31807
rect 12584 31776 13093 31804
rect 12584 31764 12590 31776
rect 13081 31773 13093 31776
rect 13127 31773 13139 31807
rect 13188 31804 13216 31844
rect 13814 31832 13820 31884
rect 13872 31872 13878 31884
rect 14093 31875 14151 31881
rect 14093 31872 14105 31875
rect 13872 31844 14105 31872
rect 13872 31832 13878 31844
rect 14093 31841 14105 31844
rect 14139 31841 14151 31875
rect 14093 31835 14151 31841
rect 15470 31832 15476 31884
rect 15528 31872 15534 31884
rect 15749 31875 15807 31881
rect 15749 31872 15761 31875
rect 15528 31844 15761 31872
rect 15528 31832 15534 31844
rect 15749 31841 15761 31844
rect 15795 31841 15807 31875
rect 16316 31872 16344 31980
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 17126 31968 17132 32020
rect 17184 32008 17190 32020
rect 17405 32011 17463 32017
rect 17405 32008 17417 32011
rect 17184 31980 17417 32008
rect 17184 31968 17190 31980
rect 17405 31977 17417 31980
rect 17451 31977 17463 32011
rect 17405 31971 17463 31977
rect 18414 31968 18420 32020
rect 18472 32008 18478 32020
rect 23477 32011 23535 32017
rect 18472 31980 22508 32008
rect 18472 31968 18478 31980
rect 19521 31943 19579 31949
rect 19521 31909 19533 31943
rect 19567 31909 19579 31943
rect 19521 31903 19579 31909
rect 16485 31875 16543 31881
rect 16485 31872 16497 31875
rect 16316 31844 16497 31872
rect 15749 31835 15807 31841
rect 16485 31841 16497 31844
rect 16531 31841 16543 31875
rect 16485 31835 16543 31841
rect 16574 31832 16580 31884
rect 16632 31881 16638 31884
rect 16632 31875 16660 31881
rect 16648 31841 16660 31875
rect 16632 31835 16660 31841
rect 16761 31875 16819 31881
rect 16761 31841 16773 31875
rect 16807 31872 16819 31875
rect 16942 31872 16948 31884
rect 16807 31844 16948 31872
rect 16807 31841 16819 31844
rect 16761 31835 16819 31841
rect 16632 31832 16638 31835
rect 16942 31832 16948 31844
rect 17000 31832 17006 31884
rect 18046 31832 18052 31884
rect 18104 31872 18110 31884
rect 18414 31872 18420 31884
rect 18104 31844 18420 31872
rect 18104 31832 18110 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 19536 31872 19564 31903
rect 20530 31900 20536 31952
rect 20588 31900 20594 31952
rect 20625 31943 20683 31949
rect 20625 31909 20637 31943
rect 20671 31940 20683 31943
rect 20714 31940 20720 31952
rect 20671 31912 20720 31940
rect 20671 31909 20683 31912
rect 20625 31903 20683 31909
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31909 20959 31943
rect 20901 31903 20959 31909
rect 21177 31943 21235 31949
rect 21177 31909 21189 31943
rect 21223 31940 21235 31943
rect 21637 31943 21695 31949
rect 21223 31912 21588 31940
rect 21223 31909 21235 31912
rect 21177 31903 21235 31909
rect 19536 31844 20116 31872
rect 13188 31776 14044 31804
rect 13081 31767 13139 31773
rect 12360 31736 12388 31764
rect 7524 31708 9352 31736
rect 11072 31708 12388 31736
rect 7524 31696 7530 31708
rect 3016 31640 4108 31668
rect 3016 31628 3022 31640
rect 5810 31628 5816 31680
rect 5868 31668 5874 31680
rect 6362 31668 6368 31680
rect 5868 31640 6368 31668
rect 5868 31628 5874 31640
rect 6362 31628 6368 31640
rect 6420 31628 6426 31680
rect 6730 31628 6736 31680
rect 6788 31668 6794 31680
rect 6825 31671 6883 31677
rect 6825 31668 6837 31671
rect 6788 31640 6837 31668
rect 6788 31628 6794 31640
rect 6825 31637 6837 31640
rect 6871 31637 6883 31671
rect 6825 31631 6883 31637
rect 9030 31628 9036 31680
rect 9088 31668 9094 31680
rect 9214 31668 9220 31680
rect 9088 31640 9220 31668
rect 9088 31628 9094 31640
rect 9214 31628 9220 31640
rect 9272 31628 9278 31680
rect 9324 31668 9352 31708
rect 11238 31668 11244 31680
rect 9324 31640 11244 31668
rect 11238 31628 11244 31640
rect 11296 31628 11302 31680
rect 12066 31628 12072 31680
rect 12124 31628 12130 31680
rect 13173 31671 13231 31677
rect 13173 31637 13185 31671
rect 13219 31668 13231 31671
rect 13538 31668 13544 31680
rect 13219 31640 13544 31668
rect 13219 31637 13231 31640
rect 13173 31631 13231 31637
rect 13538 31628 13544 31640
rect 13596 31628 13602 31680
rect 14016 31668 14044 31776
rect 14274 31764 14280 31816
rect 14332 31804 14338 31816
rect 14367 31807 14425 31813
rect 14367 31804 14379 31807
rect 14332 31776 14379 31804
rect 14332 31764 14338 31776
rect 14367 31773 14379 31776
rect 14413 31773 14425 31807
rect 15286 31804 15292 31816
rect 14367 31767 14425 31773
rect 14476 31776 15292 31804
rect 14476 31668 14504 31776
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 15562 31764 15568 31816
rect 15620 31764 15626 31816
rect 20088 31813 20116 31844
rect 19705 31807 19763 31813
rect 19705 31773 19717 31807
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 20073 31807 20131 31813
rect 20073 31773 20085 31807
rect 20119 31773 20131 31807
rect 20073 31767 20131 31773
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31804 20223 31807
rect 20548 31804 20576 31900
rect 20916 31872 20944 31903
rect 20916 31844 21404 31872
rect 21376 31813 21404 31844
rect 20809 31807 20867 31813
rect 20809 31804 20821 31807
rect 20211 31776 20484 31804
rect 20548 31776 20821 31804
rect 20211 31773 20223 31776
rect 20165 31767 20223 31773
rect 19518 31696 19524 31748
rect 19576 31736 19582 31748
rect 19720 31736 19748 31767
rect 19576 31708 19748 31736
rect 19576 31696 19582 31708
rect 14016 31640 14504 31668
rect 16114 31628 16120 31680
rect 16172 31668 16178 31680
rect 16574 31668 16580 31680
rect 16172 31640 16580 31668
rect 16172 31628 16178 31640
rect 16574 31628 16580 31640
rect 16632 31628 16638 31680
rect 20456 31668 20484 31776
rect 20809 31773 20821 31776
rect 20855 31773 20867 31807
rect 20809 31767 20867 31773
rect 21085 31807 21143 31813
rect 21085 31773 21097 31807
rect 21131 31773 21143 31807
rect 21085 31767 21143 31773
rect 21361 31807 21419 31813
rect 21361 31773 21373 31807
rect 21407 31773 21419 31807
rect 21560 31804 21588 31912
rect 21637 31909 21649 31943
rect 21683 31940 21695 31943
rect 22480 31940 22508 31980
rect 23477 31977 23489 32011
rect 23523 32008 23535 32011
rect 24118 32008 24124 32020
rect 23523 31980 24124 32008
rect 23523 31977 23535 31980
rect 23477 31971 23535 31977
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 23750 31940 23756 31952
rect 21683 31912 22094 31940
rect 22480 31912 23756 31940
rect 21683 31909 21695 31912
rect 21637 31903 21695 31909
rect 21726 31832 21732 31884
rect 21784 31872 21790 31884
rect 22066 31872 22094 31912
rect 23750 31900 23756 31912
rect 23808 31900 23814 31952
rect 21784 31844 21956 31872
rect 22066 31844 23888 31872
rect 21784 31832 21790 31844
rect 21821 31807 21879 31813
rect 21821 31804 21833 31807
rect 21560 31776 21833 31804
rect 21361 31767 21419 31773
rect 21821 31773 21833 31776
rect 21867 31773 21879 31807
rect 21928 31804 21956 31844
rect 23474 31804 23480 31816
rect 21928 31776 23480 31804
rect 21821 31767 21879 31773
rect 21100 31736 21128 31767
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 23860 31813 23888 31844
rect 23952 31844 25544 31872
rect 23661 31807 23719 31813
rect 23661 31773 23673 31807
rect 23707 31804 23719 31807
rect 23845 31807 23903 31813
rect 23707 31776 23796 31804
rect 23707 31773 23719 31776
rect 23661 31767 23719 31773
rect 20732 31708 21128 31736
rect 23768 31736 23796 31776
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 23952 31736 23980 31844
rect 25516 31816 25544 31844
rect 24213 31807 24271 31813
rect 24213 31773 24225 31807
rect 24259 31804 24271 31807
rect 25130 31804 25136 31816
rect 24259 31776 25136 31804
rect 24259 31773 24271 31776
rect 24213 31767 24271 31773
rect 25130 31764 25136 31776
rect 25188 31764 25194 31816
rect 25498 31764 25504 31816
rect 25556 31764 25562 31816
rect 23768 31708 23980 31736
rect 20530 31668 20536 31680
rect 20456 31640 20536 31668
rect 20530 31628 20536 31640
rect 20588 31628 20594 31680
rect 20622 31628 20628 31680
rect 20680 31668 20686 31680
rect 20732 31668 20760 31708
rect 20680 31640 20760 31668
rect 20680 31628 20686 31640
rect 21174 31628 21180 31680
rect 21232 31668 21238 31680
rect 24302 31668 24308 31680
rect 21232 31640 24308 31668
rect 21232 31628 21238 31640
rect 24302 31628 24308 31640
rect 24360 31628 24366 31680
rect 1104 31578 25000 31600
rect 1104 31526 6884 31578
rect 6936 31526 6948 31578
rect 7000 31526 7012 31578
rect 7064 31526 7076 31578
rect 7128 31526 7140 31578
rect 7192 31526 12818 31578
rect 12870 31526 12882 31578
rect 12934 31526 12946 31578
rect 12998 31526 13010 31578
rect 13062 31526 13074 31578
rect 13126 31526 18752 31578
rect 18804 31526 18816 31578
rect 18868 31526 18880 31578
rect 18932 31526 18944 31578
rect 18996 31526 19008 31578
rect 19060 31526 24686 31578
rect 24738 31526 24750 31578
rect 24802 31526 24814 31578
rect 24866 31526 24878 31578
rect 24930 31526 24942 31578
rect 24994 31526 25000 31578
rect 1104 31504 25000 31526
rect 1762 31464 1768 31476
rect 1686 31436 1768 31464
rect 1686 31347 1714 31436
rect 1762 31424 1768 31436
rect 1820 31464 1826 31476
rect 1946 31464 1952 31476
rect 1820 31436 1952 31464
rect 1820 31424 1826 31436
rect 1946 31424 1952 31436
rect 2004 31424 2010 31476
rect 3694 31424 3700 31476
rect 3752 31464 3758 31476
rect 3881 31467 3939 31473
rect 3881 31464 3893 31467
rect 3752 31436 3893 31464
rect 3752 31424 3758 31436
rect 3881 31433 3893 31436
rect 3927 31433 3939 31467
rect 7190 31464 7196 31476
rect 3881 31427 3939 31433
rect 4080 31436 6316 31464
rect 4080 31396 4108 31436
rect 3068 31368 4108 31396
rect 4157 31399 4215 31405
rect 1671 31341 1729 31347
rect 1671 31307 1683 31341
rect 1717 31307 1729 31341
rect 3068 31337 3096 31368
rect 4157 31365 4169 31399
rect 4203 31396 4215 31399
rect 4338 31396 4344 31408
rect 4203 31368 4344 31396
rect 4203 31365 4215 31368
rect 4157 31359 4215 31365
rect 4338 31356 4344 31368
rect 4396 31356 4402 31408
rect 4430 31356 4436 31408
rect 4488 31356 4494 31408
rect 4522 31356 4528 31408
rect 4580 31356 4586 31408
rect 5261 31399 5319 31405
rect 5261 31396 5273 31399
rect 4816 31368 5273 31396
rect 1671 31301 1729 31307
rect 3053 31331 3111 31337
rect 3053 31297 3065 31331
rect 3099 31297 3111 31331
rect 3053 31291 3111 31297
rect 3697 31331 3755 31337
rect 3697 31297 3709 31331
rect 3743 31328 3755 31331
rect 4816 31328 4844 31368
rect 5261 31365 5273 31368
rect 5307 31396 5319 31399
rect 5442 31396 5448 31408
rect 5307 31368 5448 31396
rect 5307 31365 5319 31368
rect 5261 31359 5319 31365
rect 5442 31356 5448 31368
rect 5500 31356 5506 31408
rect 3743 31300 4844 31328
rect 4893 31331 4951 31337
rect 3743 31297 3755 31300
rect 3697 31291 3755 31297
rect 4893 31297 4905 31331
rect 4939 31328 4951 31331
rect 5534 31328 5540 31340
rect 4939 31300 5540 31328
rect 4939 31297 4951 31300
rect 4893 31291 4951 31297
rect 5534 31288 5540 31300
rect 5592 31288 5598 31340
rect 6288 31328 6316 31436
rect 6380 31436 6868 31464
rect 6380 31408 6408 31436
rect 6362 31356 6368 31408
rect 6420 31356 6426 31408
rect 6454 31356 6460 31408
rect 6512 31396 6518 31408
rect 6840 31405 6868 31436
rect 6932 31436 7196 31464
rect 6932 31405 6960 31436
rect 7190 31424 7196 31436
rect 7248 31424 7254 31476
rect 7558 31424 7564 31476
rect 7616 31464 7622 31476
rect 7834 31464 7840 31476
rect 7616 31436 7840 31464
rect 7616 31424 7622 31436
rect 7834 31424 7840 31436
rect 7892 31424 7898 31476
rect 8665 31467 8723 31473
rect 8665 31433 8677 31467
rect 8711 31464 8723 31467
rect 8711 31436 12296 31464
rect 8711 31433 8723 31436
rect 8665 31427 8723 31433
rect 6549 31399 6607 31405
rect 6549 31396 6561 31399
rect 6512 31368 6561 31396
rect 6512 31356 6518 31368
rect 6549 31365 6561 31368
rect 6595 31365 6607 31399
rect 6549 31359 6607 31365
rect 6825 31399 6883 31405
rect 6825 31365 6837 31399
rect 6871 31365 6883 31399
rect 6825 31359 6883 31365
rect 6917 31399 6975 31405
rect 6917 31365 6929 31399
rect 6963 31365 6975 31399
rect 6917 31359 6975 31365
rect 7208 31368 7420 31396
rect 7208 31328 7236 31368
rect 6288 31300 7236 31328
rect 7282 31288 7288 31340
rect 7340 31288 7346 31340
rect 7392 31328 7420 31368
rect 7466 31356 7472 31408
rect 7524 31396 7530 31408
rect 7653 31399 7711 31405
rect 7653 31396 7665 31399
rect 7524 31368 7665 31396
rect 7524 31356 7530 31368
rect 7653 31365 7665 31368
rect 7699 31365 7711 31399
rect 7653 31359 7711 31365
rect 8938 31356 8944 31408
rect 8996 31356 9002 31408
rect 9030 31356 9036 31408
rect 9088 31356 9094 31408
rect 9324 31368 9720 31396
rect 9324 31328 9352 31368
rect 7392 31300 9352 31328
rect 9398 31288 9404 31340
rect 9456 31288 9462 31340
rect 9692 31328 9720 31368
rect 9766 31356 9772 31408
rect 9824 31356 9830 31408
rect 12158 31356 12164 31408
rect 12216 31356 12222 31408
rect 12268 31405 12296 31436
rect 13630 31424 13636 31476
rect 13688 31464 13694 31476
rect 22186 31464 22192 31476
rect 13688 31436 22192 31464
rect 13688 31424 13694 31436
rect 22186 31424 22192 31436
rect 22244 31424 22250 31476
rect 12253 31399 12311 31405
rect 12253 31365 12265 31399
rect 12299 31396 12311 31399
rect 14642 31396 14648 31408
rect 12299 31368 14648 31396
rect 12299 31365 12311 31368
rect 12253 31359 12311 31365
rect 14642 31356 14648 31368
rect 14700 31356 14706 31408
rect 15102 31356 15108 31408
rect 15160 31396 15166 31408
rect 17310 31396 17316 31408
rect 15160 31368 15332 31396
rect 15160 31356 15166 31368
rect 15304 31358 15332 31368
rect 16684 31368 17316 31396
rect 15363 31361 15421 31367
rect 15363 31358 15375 31361
rect 10594 31328 10600 31340
rect 9692 31300 10600 31328
rect 10594 31288 10600 31300
rect 10652 31288 10658 31340
rect 11609 31331 11667 31337
rect 11609 31297 11621 31331
rect 11655 31328 11667 31331
rect 12176 31328 12204 31356
rect 12771 31331 12829 31337
rect 12771 31328 12783 31331
rect 11655 31300 12112 31328
rect 12176 31300 12783 31328
rect 11655 31297 11667 31300
rect 11609 31291 11667 31297
rect 1394 31220 1400 31272
rect 1452 31220 1458 31272
rect 2777 31263 2835 31269
rect 2777 31229 2789 31263
rect 2823 31229 2835 31263
rect 2777 31223 2835 31229
rect 2792 31192 2820 31223
rect 3326 31220 3332 31272
rect 3384 31260 3390 31272
rect 3384 31232 4002 31260
rect 3384 31220 3390 31232
rect 6730 31220 6736 31272
rect 6788 31220 6794 31272
rect 9214 31220 9220 31272
rect 9272 31220 9278 31272
rect 2056 31164 2820 31192
rect 1302 31084 1308 31136
rect 1360 31124 1366 31136
rect 2056 31124 2084 31164
rect 5442 31152 5448 31204
rect 5500 31192 5506 31204
rect 6178 31192 6184 31204
rect 5500 31164 6184 31192
rect 5500 31152 5506 31164
rect 6178 31152 6184 31164
rect 6236 31152 6242 31204
rect 7834 31152 7840 31204
rect 7892 31152 7898 31204
rect 9953 31195 10011 31201
rect 9953 31161 9965 31195
rect 9999 31192 10011 31195
rect 10870 31192 10876 31204
rect 9999 31164 10876 31192
rect 9999 31161 10011 31164
rect 9953 31155 10011 31161
rect 10870 31152 10876 31164
rect 10928 31152 10934 31204
rect 1360 31096 2084 31124
rect 1360 31084 1366 31096
rect 2222 31084 2228 31136
rect 2280 31124 2286 31136
rect 2409 31127 2467 31133
rect 2409 31124 2421 31127
rect 2280 31096 2421 31124
rect 2280 31084 2286 31096
rect 2409 31093 2421 31096
rect 2455 31093 2467 31127
rect 6196 31124 6224 31152
rect 6546 31124 6552 31136
rect 6196 31096 6552 31124
rect 2409 31087 2467 31093
rect 6546 31084 6552 31096
rect 6604 31084 6610 31136
rect 11698 31084 11704 31136
rect 11756 31084 11762 31136
rect 12084 31124 12112 31300
rect 12771 31297 12783 31300
rect 12817 31297 12829 31331
rect 13906 31328 13912 31340
rect 12771 31291 12829 31297
rect 13832 31300 13912 31328
rect 12342 31220 12348 31272
rect 12400 31260 12406 31272
rect 12529 31263 12587 31269
rect 12529 31260 12541 31263
rect 12400 31232 12541 31260
rect 12400 31220 12406 31232
rect 12529 31229 12541 31232
rect 12575 31229 12587 31263
rect 12529 31223 12587 31229
rect 12434 31152 12440 31204
rect 12492 31152 12498 31204
rect 13541 31195 13599 31201
rect 13541 31161 13553 31195
rect 13587 31192 13599 31195
rect 13832 31192 13860 31300
rect 13906 31288 13912 31300
rect 13964 31288 13970 31340
rect 14093 31331 14151 31337
rect 14093 31297 14105 31331
rect 14139 31326 14151 31331
rect 15304 31330 15375 31358
rect 15362 31327 15375 31330
rect 15409 31328 15421 31361
rect 16298 31328 16304 31340
rect 15409 31327 16304 31328
rect 14139 31298 14226 31326
rect 15362 31300 16304 31327
rect 14139 31297 14151 31298
rect 14093 31291 14151 31297
rect 14198 31260 14226 31298
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 16684 31337 16712 31368
rect 17310 31356 17316 31368
rect 17368 31356 17374 31408
rect 23290 31396 23296 31408
rect 17880 31368 23296 31396
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 14642 31260 14648 31272
rect 14198 31232 14648 31260
rect 14642 31220 14648 31232
rect 14700 31220 14706 31272
rect 15105 31263 15163 31269
rect 15105 31229 15117 31263
rect 15151 31229 15163 31263
rect 16684 31260 16712 31291
rect 16850 31288 16856 31340
rect 16908 31328 16914 31340
rect 16943 31331 17001 31337
rect 16943 31328 16955 31331
rect 16908 31300 16955 31328
rect 16908 31288 16914 31300
rect 16943 31297 16955 31300
rect 16989 31328 17001 31331
rect 17880 31328 17908 31368
rect 23290 31356 23296 31368
rect 23348 31356 23354 31408
rect 16989 31300 17908 31328
rect 16989 31297 17001 31300
rect 16943 31291 17001 31297
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18233 31331 18291 31337
rect 18233 31328 18245 31331
rect 18012 31300 18245 31328
rect 18012 31288 18018 31300
rect 18233 31297 18245 31300
rect 18279 31297 18291 31331
rect 18233 31291 18291 31297
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31297 18567 31331
rect 19794 31328 19800 31340
rect 19755 31300 19800 31328
rect 18509 31291 18567 31297
rect 18524 31260 18552 31291
rect 19794 31288 19800 31300
rect 19852 31288 19858 31340
rect 20162 31288 20168 31340
rect 20220 31288 20226 31340
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 20772 31300 21097 31328
rect 20772 31288 20778 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 21450 31288 21456 31340
rect 21508 31288 21514 31340
rect 22186 31288 22192 31340
rect 22244 31328 22250 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22244 31300 22477 31328
rect 22244 31288 22250 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 23109 31331 23167 31337
rect 23109 31297 23121 31331
rect 23155 31297 23167 31331
rect 23753 31331 23811 31337
rect 23753 31328 23765 31331
rect 23109 31291 23167 31297
rect 23400 31300 23765 31328
rect 15105 31223 15163 31229
rect 15764 31232 16712 31260
rect 18064 31232 18552 31260
rect 19521 31263 19579 31269
rect 14918 31192 14924 31204
rect 13587 31164 13860 31192
rect 13924 31164 14924 31192
rect 13587 31161 13599 31164
rect 13541 31155 13599 31161
rect 12158 31124 12164 31136
rect 12084 31096 12164 31124
rect 12158 31084 12164 31096
rect 12216 31124 12222 31136
rect 13924 31124 13952 31164
rect 14918 31152 14924 31164
rect 14976 31152 14982 31204
rect 12216 31096 13952 31124
rect 12216 31084 12222 31096
rect 13998 31084 14004 31136
rect 14056 31084 14062 31136
rect 14458 31084 14464 31136
rect 14516 31124 14522 31136
rect 15120 31124 15148 31223
rect 15764 31124 15792 31232
rect 18064 31201 18092 31232
rect 19521 31229 19533 31263
rect 19567 31229 19579 31263
rect 19521 31223 19579 31229
rect 18049 31195 18107 31201
rect 18049 31161 18061 31195
rect 18095 31161 18107 31195
rect 18049 31155 18107 31161
rect 14516 31096 15792 31124
rect 14516 31084 14522 31096
rect 16114 31084 16120 31136
rect 16172 31084 16178 31136
rect 17402 31084 17408 31136
rect 17460 31124 17466 31136
rect 17681 31127 17739 31133
rect 17681 31124 17693 31127
rect 17460 31096 17693 31124
rect 17460 31084 17466 31096
rect 17681 31093 17693 31096
rect 17727 31093 17739 31127
rect 17681 31087 17739 31093
rect 18598 31084 18604 31136
rect 18656 31084 18662 31136
rect 19536 31124 19564 31223
rect 20180 31124 20208 31288
rect 20901 31263 20959 31269
rect 20901 31229 20913 31263
rect 20947 31229 20959 31263
rect 23124 31260 23152 31291
rect 20901 31223 20959 31229
rect 22296 31232 23152 31260
rect 20533 31195 20591 31201
rect 20533 31161 20545 31195
rect 20579 31192 20591 31195
rect 20622 31192 20628 31204
rect 20579 31164 20628 31192
rect 20579 31161 20591 31164
rect 20533 31155 20591 31161
rect 20622 31152 20628 31164
rect 20680 31192 20686 31204
rect 20916 31192 20944 31223
rect 22296 31201 22324 31232
rect 20680 31164 20944 31192
rect 22281 31195 22339 31201
rect 20680 31152 20686 31164
rect 22281 31161 22293 31195
rect 22327 31161 22339 31195
rect 22281 31155 22339 31161
rect 22925 31195 22983 31201
rect 22925 31161 22937 31195
rect 22971 31192 22983 31195
rect 23400 31192 23428 31300
rect 23753 31297 23765 31300
rect 23799 31297 23811 31331
rect 23753 31291 23811 31297
rect 23842 31288 23848 31340
rect 23900 31328 23906 31340
rect 24121 31331 24179 31337
rect 24121 31328 24133 31331
rect 23900 31300 24133 31328
rect 23900 31288 23906 31300
rect 24121 31297 24133 31300
rect 24167 31297 24179 31331
rect 24121 31291 24179 31297
rect 24213 31331 24271 31337
rect 24213 31297 24225 31331
rect 24259 31297 24271 31331
rect 24213 31291 24271 31297
rect 24228 31260 24256 31291
rect 23584 31232 24256 31260
rect 23584 31201 23612 31232
rect 22971 31164 23428 31192
rect 23569 31195 23627 31201
rect 22971 31161 22983 31164
rect 22925 31155 22983 31161
rect 23569 31161 23581 31195
rect 23615 31161 23627 31195
rect 23569 31155 23627 31161
rect 19536 31096 20208 31124
rect 21358 31084 21364 31136
rect 21416 31084 21422 31136
rect 23934 31084 23940 31136
rect 23992 31084 23998 31136
rect 24394 31084 24400 31136
rect 24452 31084 24458 31136
rect 1104 31034 24840 31056
rect 1104 30982 3917 31034
rect 3969 30982 3981 31034
rect 4033 30982 4045 31034
rect 4097 30982 4109 31034
rect 4161 30982 4173 31034
rect 4225 30982 9851 31034
rect 9903 30982 9915 31034
rect 9967 30982 9979 31034
rect 10031 30982 10043 31034
rect 10095 30982 10107 31034
rect 10159 30982 15785 31034
rect 15837 30982 15849 31034
rect 15901 30982 15913 31034
rect 15965 30982 15977 31034
rect 16029 30982 16041 31034
rect 16093 30982 21719 31034
rect 21771 30982 21783 31034
rect 21835 30982 21847 31034
rect 21899 30982 21911 31034
rect 21963 30982 21975 31034
rect 22027 30982 24840 31034
rect 1104 30960 24840 30982
rect 1578 30880 1584 30932
rect 1636 30920 1642 30932
rect 2314 30920 2320 30932
rect 1636 30892 2320 30920
rect 1636 30880 1642 30892
rect 2314 30880 2320 30892
rect 2372 30880 2378 30932
rect 3326 30880 3332 30932
rect 3384 30880 3390 30932
rect 4522 30880 4528 30932
rect 4580 30920 4586 30932
rect 5261 30923 5319 30929
rect 5261 30920 5273 30923
rect 4580 30892 5273 30920
rect 4580 30880 4586 30892
rect 5261 30889 5273 30892
rect 5307 30889 5319 30923
rect 5261 30883 5319 30889
rect 5994 30880 6000 30932
rect 6052 30920 6058 30932
rect 6052 30892 7052 30920
rect 6052 30880 6058 30892
rect 7024 30852 7052 30892
rect 7190 30880 7196 30932
rect 7248 30920 7254 30932
rect 7377 30923 7435 30929
rect 7377 30920 7389 30923
rect 7248 30892 7389 30920
rect 7248 30880 7254 30892
rect 7377 30889 7389 30892
rect 7423 30889 7435 30923
rect 7377 30883 7435 30889
rect 9030 30880 9036 30932
rect 9088 30920 9094 30932
rect 9953 30923 10011 30929
rect 9953 30920 9965 30923
rect 9088 30892 9965 30920
rect 9088 30880 9094 30892
rect 9953 30889 9965 30892
rect 9999 30889 10011 30923
rect 9953 30883 10011 30889
rect 10134 30880 10140 30932
rect 10192 30880 10198 30932
rect 12342 30880 12348 30932
rect 12400 30880 12406 30932
rect 12526 30880 12532 30932
rect 12584 30880 12590 30932
rect 12805 30923 12863 30929
rect 12805 30889 12817 30923
rect 12851 30920 12863 30923
rect 12851 30892 13952 30920
rect 12851 30889 12863 30892
rect 12805 30883 12863 30889
rect 8386 30852 8392 30864
rect 7024 30824 8392 30852
rect 8386 30812 8392 30824
rect 8444 30812 8450 30864
rect 10152 30852 10180 30880
rect 11054 30852 11060 30864
rect 10152 30824 11060 30852
rect 11054 30812 11060 30824
rect 11112 30812 11118 30864
rect 6270 30744 6276 30796
rect 6328 30784 6334 30796
rect 6365 30787 6423 30793
rect 6365 30784 6377 30787
rect 6328 30756 6377 30784
rect 6328 30744 6334 30756
rect 6365 30753 6377 30756
rect 6411 30753 6423 30787
rect 6365 30747 6423 30753
rect 8294 30744 8300 30796
rect 8352 30784 8358 30796
rect 8938 30784 8944 30796
rect 8352 30756 8944 30784
rect 8352 30744 8358 30756
rect 8938 30744 8944 30756
rect 8996 30744 9002 30796
rect 10410 30744 10416 30796
rect 10468 30784 10474 30796
rect 10505 30787 10563 30793
rect 10505 30784 10517 30787
rect 10468 30756 10517 30784
rect 10468 30744 10474 30756
rect 10505 30753 10517 30756
rect 10551 30753 10563 30787
rect 10505 30747 10563 30753
rect 10778 30744 10784 30796
rect 10836 30744 10842 30796
rect 11146 30744 11152 30796
rect 11204 30744 11210 30796
rect 11422 30744 11428 30796
rect 11480 30744 11486 30796
rect 11514 30744 11520 30796
rect 11572 30793 11578 30796
rect 11572 30787 11600 30793
rect 11588 30753 11600 30787
rect 11572 30747 11600 30753
rect 11701 30787 11759 30793
rect 11701 30753 11713 30787
rect 11747 30784 11759 30787
rect 11882 30784 11888 30796
rect 11747 30756 11888 30784
rect 11747 30753 11759 30756
rect 11701 30747 11759 30753
rect 11572 30744 11578 30747
rect 11882 30744 11888 30756
rect 11940 30784 11946 30796
rect 12066 30784 12072 30796
rect 11940 30756 12072 30784
rect 11940 30744 11946 30756
rect 12066 30744 12072 30756
rect 12124 30744 12130 30796
rect 12360 30784 12388 30880
rect 13924 30852 13952 30892
rect 14642 30880 14648 30932
rect 14700 30880 14706 30932
rect 16114 30880 16120 30932
rect 16172 30920 16178 30932
rect 16172 30892 16436 30920
rect 16172 30880 16178 30892
rect 14660 30852 14688 30880
rect 16408 30861 16436 30892
rect 17402 30880 17408 30932
rect 17460 30880 17466 30932
rect 17589 30923 17647 30929
rect 17589 30889 17601 30923
rect 17635 30920 17647 30923
rect 17954 30920 17960 30932
rect 17635 30892 17960 30920
rect 17635 30889 17647 30892
rect 17589 30883 17647 30889
rect 13924 30824 14688 30852
rect 16393 30855 16451 30861
rect 16393 30821 16405 30855
rect 16439 30821 16451 30855
rect 16393 30815 16451 30821
rect 12526 30784 12532 30796
rect 12360 30756 12532 30784
rect 12526 30744 12532 30756
rect 12584 30744 12590 30796
rect 13906 30744 13912 30796
rect 13964 30744 13970 30796
rect 13998 30744 14004 30796
rect 14056 30784 14062 30796
rect 14056 30756 14964 30784
rect 14056 30744 14062 30756
rect 2130 30676 2136 30728
rect 2188 30716 2194 30728
rect 2317 30719 2375 30725
rect 2317 30716 2329 30719
rect 2188 30688 2329 30716
rect 2188 30676 2194 30688
rect 2317 30685 2329 30688
rect 2363 30685 2375 30719
rect 2590 30716 2596 30728
rect 2551 30688 2596 30716
rect 2317 30679 2375 30685
rect 1486 30608 1492 30660
rect 1544 30608 1550 30660
rect 1670 30608 1676 30660
rect 1728 30608 1734 30660
rect 2332 30648 2360 30679
rect 2590 30676 2596 30688
rect 2648 30676 2654 30728
rect 3786 30676 3792 30728
rect 3844 30676 3850 30728
rect 4154 30676 4160 30728
rect 4212 30716 4218 30728
rect 4249 30719 4307 30725
rect 4249 30716 4261 30719
rect 4212 30688 4261 30716
rect 4212 30676 4218 30688
rect 4249 30685 4261 30688
rect 4295 30685 4307 30719
rect 4249 30679 4307 30685
rect 4430 30676 4436 30728
rect 4488 30716 4494 30728
rect 4523 30719 4581 30725
rect 4523 30716 4535 30719
rect 4488 30688 4535 30716
rect 4488 30676 4494 30688
rect 4523 30685 4535 30688
rect 4569 30716 4581 30719
rect 5350 30716 5356 30728
rect 4569 30688 5356 30716
rect 4569 30685 4581 30688
rect 4523 30679 4581 30685
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 6639 30719 6697 30725
rect 6639 30685 6651 30719
rect 6685 30716 6697 30719
rect 6685 30688 6868 30716
rect 6685 30685 6697 30688
rect 6639 30679 6697 30685
rect 4172 30648 4200 30676
rect 6840 30660 6868 30688
rect 9122 30676 9128 30728
rect 9180 30716 9186 30728
rect 9215 30719 9273 30725
rect 9215 30716 9227 30719
rect 9180 30688 9227 30716
rect 9180 30676 9186 30688
rect 9215 30685 9227 30688
rect 9261 30685 9273 30719
rect 9215 30679 9273 30685
rect 10594 30676 10600 30728
rect 10652 30716 10658 30728
rect 10689 30719 10747 30725
rect 10689 30716 10701 30719
rect 10652 30688 10701 30716
rect 10652 30676 10658 30688
rect 10689 30685 10701 30688
rect 10735 30716 10747 30719
rect 10796 30716 10824 30744
rect 10735 30688 10824 30716
rect 12345 30719 12403 30725
rect 10735 30685 10747 30688
rect 10689 30679 10747 30685
rect 12345 30685 12357 30719
rect 12391 30716 12403 30719
rect 12713 30719 12771 30725
rect 12713 30716 12725 30719
rect 12391 30688 12725 30716
rect 12391 30685 12403 30688
rect 12345 30679 12403 30685
rect 12713 30685 12725 30688
rect 12759 30685 12771 30719
rect 12713 30679 12771 30685
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30685 13047 30719
rect 13924 30716 13952 30744
rect 14936 30725 14964 30756
rect 15102 30744 15108 30796
rect 15160 30744 15166 30796
rect 15562 30744 15568 30796
rect 15620 30784 15626 30796
rect 15620 30756 15976 30784
rect 15620 30744 15626 30756
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13924 30688 14105 30716
rect 12989 30679 13047 30685
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14093 30679 14151 30685
rect 14461 30719 14519 30725
rect 14461 30685 14473 30719
rect 14507 30685 14519 30719
rect 14461 30679 14519 30685
rect 14921 30719 14979 30725
rect 14921 30685 14933 30719
rect 14967 30685 14979 30719
rect 14921 30679 14979 30685
rect 2332 30620 4200 30648
rect 4338 30608 4344 30660
rect 4396 30608 4402 30660
rect 6822 30608 6828 30660
rect 6880 30608 6886 30660
rect 10318 30608 10324 30660
rect 10376 30648 10382 30660
rect 10502 30648 10508 30660
rect 10376 30620 10508 30648
rect 10376 30608 10382 30620
rect 10502 30608 10508 30620
rect 10560 30608 10566 30660
rect 934 30540 940 30592
rect 992 30580 998 30592
rect 1210 30580 1216 30592
rect 992 30552 1216 30580
rect 992 30540 998 30552
rect 1210 30540 1216 30552
rect 1268 30540 1274 30592
rect 3973 30583 4031 30589
rect 3973 30549 3985 30583
rect 4019 30580 4031 30583
rect 4246 30580 4252 30592
rect 4019 30552 4252 30580
rect 4019 30549 4031 30552
rect 3973 30543 4031 30549
rect 4246 30540 4252 30552
rect 4304 30540 4310 30592
rect 4356 30580 4384 30608
rect 12158 30580 12164 30592
rect 4356 30552 12164 30580
rect 12158 30540 12164 30552
rect 12216 30540 12222 30592
rect 12342 30540 12348 30592
rect 12400 30580 12406 30592
rect 13004 30580 13032 30679
rect 13538 30608 13544 30660
rect 13596 30648 13602 30660
rect 14476 30648 14504 30679
rect 15286 30676 15292 30728
rect 15344 30716 15350 30728
rect 15948 30725 15976 30756
rect 16758 30744 16764 30796
rect 16816 30793 16822 30796
rect 16816 30787 16844 30793
rect 16832 30753 16844 30787
rect 16816 30747 16844 30753
rect 16945 30787 17003 30793
rect 16945 30753 16957 30787
rect 16991 30784 17003 30787
rect 17420 30784 17448 30880
rect 16991 30756 17448 30784
rect 16991 30753 17003 30756
rect 16945 30747 17003 30753
rect 16816 30744 16822 30747
rect 15749 30719 15807 30725
rect 15749 30716 15761 30719
rect 15344 30688 15761 30716
rect 15344 30676 15350 30688
rect 15749 30685 15761 30688
rect 15795 30685 15807 30719
rect 15749 30679 15807 30685
rect 15933 30719 15991 30725
rect 15933 30685 15945 30719
rect 15979 30716 15991 30719
rect 16114 30716 16120 30728
rect 15979 30688 16120 30716
rect 15979 30685 15991 30688
rect 15933 30679 15991 30685
rect 16114 30676 16120 30688
rect 16172 30676 16178 30728
rect 16666 30676 16672 30728
rect 16724 30676 16730 30728
rect 17604 30716 17632 30883
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 18598 30880 18604 30932
rect 18656 30920 18662 30932
rect 19337 30923 19395 30929
rect 19337 30920 19349 30923
rect 18656 30892 19349 30920
rect 18656 30880 18662 30892
rect 19337 30889 19349 30892
rect 19383 30889 19395 30923
rect 19337 30883 19395 30889
rect 19812 30892 20116 30920
rect 19061 30855 19119 30861
rect 19061 30821 19073 30855
rect 19107 30852 19119 30855
rect 19812 30852 19840 30892
rect 19107 30824 19840 30852
rect 19889 30855 19947 30861
rect 19107 30821 19119 30824
rect 19061 30815 19119 30821
rect 19889 30821 19901 30855
rect 19935 30821 19947 30855
rect 19889 30815 19947 30821
rect 17678 30744 17684 30796
rect 17736 30744 17742 30796
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30784 19579 30787
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19567 30756 19717 30784
rect 19567 30753 19579 30756
rect 19521 30747 19579 30753
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 17937 30719 17995 30725
rect 17937 30716 17949 30719
rect 17604 30688 17949 30716
rect 17937 30685 17949 30688
rect 17983 30685 17995 30719
rect 17937 30679 17995 30685
rect 19245 30719 19303 30725
rect 19245 30685 19257 30719
rect 19291 30716 19303 30719
rect 19613 30719 19671 30725
rect 19613 30716 19625 30719
rect 19291 30688 19625 30716
rect 19291 30685 19303 30688
rect 19245 30679 19303 30685
rect 19613 30685 19625 30688
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19797 30719 19855 30725
rect 19797 30685 19809 30719
rect 19843 30716 19855 30719
rect 19904 30716 19932 30815
rect 20088 30725 20116 30892
rect 20622 30880 20628 30932
rect 20680 30880 20686 30932
rect 20717 30923 20775 30929
rect 20717 30889 20729 30923
rect 20763 30920 20775 30923
rect 21450 30920 21456 30932
rect 20763 30892 21456 30920
rect 20763 30889 20775 30892
rect 20717 30883 20775 30889
rect 21450 30880 21456 30892
rect 21508 30880 21514 30932
rect 23109 30923 23167 30929
rect 23109 30889 23121 30923
rect 23155 30920 23167 30923
rect 23155 30892 23704 30920
rect 23155 30889 23167 30892
rect 23109 30883 23167 30889
rect 20640 30725 20668 30880
rect 22833 30855 22891 30861
rect 22833 30821 22845 30855
rect 22879 30821 22891 30855
rect 22833 30815 22891 30821
rect 23477 30855 23535 30861
rect 23477 30821 23489 30855
rect 23523 30821 23535 30855
rect 23477 30815 23535 30821
rect 19843 30688 19932 30716
rect 20073 30719 20131 30725
rect 19843 30685 19855 30688
rect 19797 30679 19855 30685
rect 20073 30685 20085 30719
rect 20119 30685 20131 30719
rect 20073 30679 20131 30685
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30685 20683 30719
rect 20625 30679 20683 30685
rect 13596 30620 14504 30648
rect 13596 30608 13602 30620
rect 19260 30592 19288 30679
rect 20806 30676 20812 30728
rect 20864 30676 20870 30728
rect 22278 30676 22284 30728
rect 22336 30676 22342 30728
rect 19521 30651 19579 30657
rect 19521 30617 19533 30651
rect 19567 30648 19579 30651
rect 22848 30648 22876 30815
rect 23492 30784 23520 30815
rect 23032 30756 23520 30784
rect 23032 30725 23060 30756
rect 23017 30719 23075 30725
rect 23017 30685 23029 30719
rect 23063 30685 23075 30719
rect 23017 30679 23075 30685
rect 23290 30676 23296 30728
rect 23348 30676 23354 30728
rect 23676 30725 23704 30892
rect 23661 30719 23719 30725
rect 23661 30685 23673 30719
rect 23707 30685 23719 30719
rect 23661 30679 23719 30685
rect 24578 30676 24584 30728
rect 24636 30716 24642 30728
rect 25866 30716 25872 30728
rect 24636 30688 25872 30716
rect 24636 30676 24642 30688
rect 25866 30676 25872 30688
rect 25924 30676 25930 30728
rect 23845 30651 23903 30657
rect 23845 30648 23857 30651
rect 19567 30620 22784 30648
rect 22848 30620 23857 30648
rect 19567 30617 19579 30620
rect 19521 30611 19579 30617
rect 12400 30552 13032 30580
rect 12400 30540 12406 30552
rect 13446 30540 13452 30592
rect 13504 30580 13510 30592
rect 14458 30580 14464 30592
rect 13504 30552 14464 30580
rect 13504 30540 13510 30552
rect 14458 30540 14464 30552
rect 14516 30540 14522 30592
rect 16298 30540 16304 30592
rect 16356 30580 16362 30592
rect 18598 30580 18604 30592
rect 16356 30552 18604 30580
rect 16356 30540 16362 30552
rect 18598 30540 18604 30552
rect 18656 30540 18662 30592
rect 19242 30540 19248 30592
rect 19300 30540 19306 30592
rect 22097 30583 22155 30589
rect 22097 30549 22109 30583
rect 22143 30580 22155 30583
rect 22554 30580 22560 30592
rect 22143 30552 22560 30580
rect 22143 30549 22155 30552
rect 22097 30543 22155 30549
rect 22554 30540 22560 30552
rect 22612 30540 22618 30592
rect 22756 30580 22784 30620
rect 23845 30617 23857 30620
rect 23891 30617 23903 30651
rect 23845 30611 23903 30617
rect 24213 30651 24271 30657
rect 24213 30617 24225 30651
rect 24259 30648 24271 30651
rect 25130 30648 25136 30660
rect 24259 30620 25136 30648
rect 24259 30617 24271 30620
rect 24213 30611 24271 30617
rect 25130 30608 25136 30620
rect 25188 30608 25194 30660
rect 23290 30580 23296 30592
rect 22756 30552 23296 30580
rect 23290 30540 23296 30552
rect 23348 30540 23354 30592
rect 23566 30540 23572 30592
rect 23624 30580 23630 30592
rect 24578 30580 24584 30592
rect 23624 30552 24584 30580
rect 23624 30540 23630 30552
rect 24578 30540 24584 30552
rect 24636 30540 24642 30592
rect 1104 30490 25000 30512
rect 1104 30438 6884 30490
rect 6936 30438 6948 30490
rect 7000 30438 7012 30490
rect 7064 30438 7076 30490
rect 7128 30438 7140 30490
rect 7192 30438 12818 30490
rect 12870 30438 12882 30490
rect 12934 30438 12946 30490
rect 12998 30438 13010 30490
rect 13062 30438 13074 30490
rect 13126 30438 18752 30490
rect 18804 30438 18816 30490
rect 18868 30438 18880 30490
rect 18932 30438 18944 30490
rect 18996 30438 19008 30490
rect 19060 30438 24686 30490
rect 24738 30438 24750 30490
rect 24802 30438 24814 30490
rect 24866 30438 24878 30490
rect 24930 30438 24942 30490
rect 24994 30438 25000 30490
rect 1104 30416 25000 30438
rect 3881 30379 3939 30385
rect 1688 30348 3188 30376
rect 1302 30268 1308 30320
rect 1360 30308 1366 30320
rect 1688 30308 1716 30348
rect 1360 30280 1716 30308
rect 3160 30308 3188 30348
rect 3881 30345 3893 30379
rect 3927 30345 3939 30379
rect 3881 30339 3939 30345
rect 3329 30311 3387 30317
rect 3329 30308 3341 30311
rect 3160 30280 3341 30308
rect 1360 30268 1366 30280
rect 3329 30277 3341 30280
rect 3375 30277 3387 30311
rect 3896 30308 3924 30339
rect 3970 30336 3976 30388
rect 4028 30376 4034 30388
rect 4430 30376 4436 30388
rect 4028 30348 4436 30376
rect 4028 30336 4034 30348
rect 4430 30336 4436 30348
rect 4488 30336 4494 30388
rect 4706 30336 4712 30388
rect 4764 30376 4770 30388
rect 10965 30379 11023 30385
rect 4764 30348 10916 30376
rect 4764 30336 4770 30348
rect 6454 30308 6460 30320
rect 3896 30280 6460 30308
rect 3329 30271 3387 30277
rect 6454 30268 6460 30280
rect 6512 30268 6518 30320
rect 9398 30308 9404 30320
rect 6564 30280 9404 30308
rect 2406 30200 2412 30252
rect 2464 30200 2470 30252
rect 2682 30200 2688 30252
rect 2740 30200 2746 30252
rect 3418 30200 3424 30252
rect 3476 30200 3482 30252
rect 3694 30200 3700 30252
rect 3752 30200 3758 30252
rect 3878 30200 3884 30252
rect 3936 30240 3942 30252
rect 4431 30243 4489 30249
rect 4431 30240 4443 30243
rect 3936 30212 4443 30240
rect 3936 30200 3942 30212
rect 4431 30209 4443 30212
rect 4477 30209 4489 30243
rect 4431 30203 4489 30209
rect 4522 30200 4528 30252
rect 4580 30240 4586 30252
rect 6564 30240 6592 30280
rect 9398 30268 9404 30280
rect 9456 30268 9462 30320
rect 10888 30308 10916 30348
rect 10965 30345 10977 30379
rect 11011 30376 11023 30379
rect 11146 30376 11152 30388
rect 11011 30348 11152 30376
rect 11011 30345 11023 30348
rect 10965 30339 11023 30345
rect 11146 30336 11152 30348
rect 11204 30336 11210 30388
rect 11514 30336 11520 30388
rect 11572 30336 11578 30388
rect 11698 30336 11704 30388
rect 11756 30376 11762 30388
rect 23566 30376 23572 30388
rect 11756 30348 23572 30376
rect 11756 30336 11762 30348
rect 23566 30336 23572 30348
rect 23624 30336 23630 30388
rect 23753 30379 23811 30385
rect 23753 30345 23765 30379
rect 23799 30376 23811 30379
rect 23842 30376 23848 30388
rect 23799 30348 23848 30376
rect 23799 30345 23811 30348
rect 23753 30339 23811 30345
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 23992 30348 24164 30376
rect 23992 30336 23998 30348
rect 11532 30308 11560 30336
rect 9968 30280 10362 30308
rect 10888 30280 11560 30308
rect 4580 30212 6592 30240
rect 7099 30243 7157 30249
rect 4580 30200 4586 30212
rect 7099 30209 7111 30243
rect 7145 30240 7157 30243
rect 7190 30240 7196 30252
rect 7145 30212 7196 30240
rect 7145 30209 7157 30212
rect 7099 30203 7157 30209
rect 7190 30200 7196 30212
rect 7248 30240 7254 30252
rect 8110 30240 8116 30252
rect 7248 30212 8116 30240
rect 7248 30200 7254 30212
rect 8110 30200 8116 30212
rect 8168 30200 8174 30252
rect 9968 30249 9996 30280
rect 9953 30243 10011 30249
rect 9953 30209 9965 30243
rect 9999 30209 10011 30243
rect 9953 30203 10011 30209
rect 10134 30200 10140 30252
rect 10192 30240 10198 30252
rect 10227 30243 10285 30249
rect 10227 30240 10239 30243
rect 10192 30212 10239 30240
rect 10192 30200 10198 30212
rect 10227 30209 10239 30212
rect 10273 30209 10285 30243
rect 10334 30240 10362 30280
rect 18230 30279 18236 30320
rect 18215 30273 18236 30279
rect 12526 30240 12532 30252
rect 10334 30212 12532 30240
rect 10227 30203 10285 30209
rect 12526 30200 12532 30212
rect 12584 30200 12590 30252
rect 13814 30200 13820 30252
rect 13872 30240 13878 30252
rect 13909 30243 13967 30249
rect 13909 30240 13921 30243
rect 13872 30212 13921 30240
rect 13872 30200 13878 30212
rect 13909 30209 13921 30212
rect 13955 30209 13967 30243
rect 13909 30203 13967 30209
rect 14090 30200 14096 30252
rect 14148 30240 14154 30252
rect 14183 30243 14241 30249
rect 14183 30240 14195 30243
rect 14148 30212 14195 30240
rect 14148 30200 14154 30212
rect 14183 30209 14195 30212
rect 14229 30240 14241 30243
rect 14229 30212 15976 30240
rect 14229 30209 14241 30212
rect 14183 30203 14241 30209
rect 1489 30175 1547 30181
rect 1489 30141 1501 30175
rect 1535 30172 1547 30175
rect 1578 30172 1584 30184
rect 1535 30144 1584 30172
rect 1535 30141 1547 30144
rect 1489 30135 1547 30141
rect 1578 30132 1584 30144
rect 1636 30132 1642 30184
rect 1670 30132 1676 30184
rect 1728 30132 1734 30184
rect 2133 30175 2191 30181
rect 2133 30141 2145 30175
rect 2179 30172 2191 30175
rect 2222 30172 2228 30184
rect 2179 30144 2228 30172
rect 2179 30141 2191 30144
rect 2133 30135 2191 30141
rect 2222 30132 2228 30144
rect 2280 30132 2286 30184
rect 2547 30175 2605 30181
rect 2547 30141 2559 30175
rect 2593 30172 2605 30175
rect 3786 30172 3792 30184
rect 2593 30144 3792 30172
rect 2593 30141 2605 30144
rect 2547 30135 2605 30141
rect 3786 30132 3792 30144
rect 3844 30132 3850 30184
rect 4154 30132 4160 30184
rect 4212 30132 4218 30184
rect 6454 30132 6460 30184
rect 6512 30172 6518 30184
rect 6825 30175 6883 30181
rect 6825 30172 6837 30175
rect 6512 30144 6837 30172
rect 6512 30132 6518 30144
rect 6825 30141 6837 30144
rect 6871 30141 6883 30175
rect 6825 30135 6883 30141
rect 7650 30132 7656 30184
rect 7708 30172 7714 30184
rect 7926 30172 7932 30184
rect 7708 30144 7932 30172
rect 7708 30132 7714 30144
rect 7926 30132 7932 30144
rect 7984 30132 7990 30184
rect 10686 30132 10692 30184
rect 10744 30172 10750 30184
rect 10962 30172 10968 30184
rect 10744 30144 10968 30172
rect 10744 30132 10750 30144
rect 10962 30132 10968 30144
rect 11020 30132 11026 30184
rect 12158 30132 12164 30184
rect 12216 30172 12222 30184
rect 13832 30172 13860 30200
rect 12216 30144 13860 30172
rect 15948 30172 15976 30212
rect 17586 30200 17592 30252
rect 17644 30240 17650 30252
rect 17862 30240 17868 30252
rect 17644 30212 17868 30240
rect 17644 30200 17650 30212
rect 17862 30200 17868 30212
rect 17920 30240 17926 30252
rect 17957 30243 18015 30249
rect 17957 30240 17969 30243
rect 17920 30212 17969 30240
rect 17920 30200 17926 30212
rect 17957 30209 17969 30212
rect 18003 30209 18015 30243
rect 18215 30239 18227 30273
rect 18288 30268 18294 30320
rect 18414 30268 18420 30320
rect 18472 30308 18478 30320
rect 19334 30308 19340 30320
rect 18472 30280 19340 30308
rect 18472 30268 18478 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 24136 30317 24164 30348
rect 24121 30311 24179 30317
rect 19444 30280 23704 30308
rect 18261 30242 18274 30268
rect 18261 30239 18273 30242
rect 18215 30233 18273 30239
rect 17957 30203 18015 30209
rect 18598 30200 18604 30252
rect 18656 30240 18662 30252
rect 19444 30240 19472 30280
rect 20530 30249 20536 30252
rect 18656 30212 19472 30240
rect 20513 30243 20536 30249
rect 18656 30200 18662 30212
rect 20513 30209 20525 30243
rect 20513 30203 20536 30209
rect 20530 30200 20536 30203
rect 20588 30200 20594 30252
rect 22095 30243 22153 30249
rect 22095 30209 22107 30243
rect 22141 30240 22153 30243
rect 22186 30240 22192 30252
rect 22141 30212 22192 30240
rect 22141 30209 22153 30212
rect 22095 30203 22153 30209
rect 22186 30200 22192 30212
rect 22244 30200 22250 30252
rect 22738 30200 22744 30252
rect 22796 30240 22802 30252
rect 23676 30249 23704 30280
rect 24121 30277 24133 30311
rect 24167 30277 24179 30311
rect 24121 30271 24179 30277
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 22796 30212 23397 30240
rect 22796 30200 22802 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 23385 30203 23443 30209
rect 23661 30243 23719 30249
rect 23661 30209 23673 30243
rect 23707 30209 23719 30243
rect 23661 30203 23719 30209
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 15948 30144 17632 30172
rect 12216 30132 12222 30144
rect 3050 29996 3056 30048
rect 3108 30036 3114 30048
rect 3605 30039 3663 30045
rect 3605 30036 3617 30039
rect 3108 30008 3617 30036
rect 3108 29996 3114 30008
rect 3605 30005 3617 30008
rect 3651 30005 3663 30039
rect 4172 30036 4200 30132
rect 8754 30104 8760 30116
rect 7760 30076 8760 30104
rect 4890 30036 4896 30048
rect 4172 30008 4896 30036
rect 3605 29999 3663 30005
rect 4890 29996 4896 30008
rect 4948 29996 4954 30048
rect 5166 29996 5172 30048
rect 5224 29996 5230 30048
rect 6270 29996 6276 30048
rect 6328 30036 6334 30048
rect 7760 30036 7788 30076
rect 8754 30064 8760 30076
rect 8812 30064 8818 30116
rect 9646 30076 10088 30104
rect 6328 30008 7788 30036
rect 6328 29996 6334 30008
rect 7834 29996 7840 30048
rect 7892 29996 7898 30048
rect 7926 29996 7932 30048
rect 7984 30036 7990 30048
rect 9646 30036 9674 30076
rect 7984 30008 9674 30036
rect 10060 30036 10088 30076
rect 11238 30064 11244 30116
rect 11296 30104 11302 30116
rect 12618 30104 12624 30116
rect 11296 30076 12624 30104
rect 11296 30064 11302 30076
rect 12618 30064 12624 30076
rect 12676 30064 12682 30116
rect 17604 30048 17632 30144
rect 19426 30132 19432 30184
rect 19484 30172 19490 30184
rect 20257 30175 20315 30181
rect 20257 30172 20269 30175
rect 19484 30144 20269 30172
rect 19484 30132 19490 30144
rect 20257 30141 20269 30144
rect 20303 30141 20315 30175
rect 21821 30175 21879 30181
rect 21821 30172 21833 30175
rect 20257 30135 20315 30141
rect 21284 30144 21833 30172
rect 18969 30107 19027 30113
rect 18969 30073 18981 30107
rect 19015 30104 19027 30107
rect 19242 30104 19248 30116
rect 19015 30076 19248 30104
rect 19015 30073 19027 30076
rect 18969 30067 19027 30073
rect 19242 30064 19248 30076
rect 19300 30064 19306 30116
rect 14734 30036 14740 30048
rect 10060 30008 14740 30036
rect 7984 29996 7990 30008
rect 14734 29996 14740 30008
rect 14792 29996 14798 30048
rect 14918 29996 14924 30048
rect 14976 29996 14982 30048
rect 17586 29996 17592 30048
rect 17644 29996 17650 30048
rect 19978 29996 19984 30048
rect 20036 30036 20042 30048
rect 21284 30036 21312 30144
rect 21821 30141 21833 30144
rect 21867 30141 21879 30175
rect 23952 30172 23980 30203
rect 21821 30135 21879 30141
rect 23492 30144 23980 30172
rect 23492 30113 23520 30144
rect 23477 30107 23535 30113
rect 23477 30073 23489 30107
rect 23523 30073 23535 30107
rect 23477 30067 23535 30073
rect 20036 30008 21312 30036
rect 21637 30039 21695 30045
rect 20036 29996 20042 30008
rect 21637 30005 21649 30039
rect 21683 30036 21695 30039
rect 22278 30036 22284 30048
rect 21683 30008 22284 30036
rect 21683 30005 21695 30008
rect 21637 29999 21695 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 22830 29996 22836 30048
rect 22888 29996 22894 30048
rect 23198 29996 23204 30048
rect 23256 29996 23262 30048
rect 24394 29996 24400 30048
rect 24452 29996 24458 30048
rect 1104 29946 24840 29968
rect 1104 29894 3917 29946
rect 3969 29894 3981 29946
rect 4033 29894 4045 29946
rect 4097 29894 4109 29946
rect 4161 29894 4173 29946
rect 4225 29894 9851 29946
rect 9903 29894 9915 29946
rect 9967 29894 9979 29946
rect 10031 29894 10043 29946
rect 10095 29894 10107 29946
rect 10159 29894 15785 29946
rect 15837 29894 15849 29946
rect 15901 29894 15913 29946
rect 15965 29894 15977 29946
rect 16029 29894 16041 29946
rect 16093 29894 21719 29946
rect 21771 29894 21783 29946
rect 21835 29894 21847 29946
rect 21899 29894 21911 29946
rect 21963 29894 21975 29946
rect 22027 29894 24840 29946
rect 1104 29872 24840 29894
rect 1578 29792 1584 29844
rect 1636 29832 1642 29844
rect 1636 29804 2360 29832
rect 1636 29792 1642 29804
rect 2332 29696 2360 29804
rect 2682 29792 2688 29844
rect 2740 29792 2746 29844
rect 2774 29792 2780 29844
rect 2832 29832 2838 29844
rect 3234 29832 3240 29844
rect 2832 29804 3240 29832
rect 2832 29792 2838 29804
rect 3234 29792 3240 29804
rect 3292 29792 3298 29844
rect 3602 29792 3608 29844
rect 3660 29792 3666 29844
rect 4706 29792 4712 29844
rect 4764 29792 4770 29844
rect 7834 29832 7840 29844
rect 7576 29804 7840 29832
rect 2958 29724 2964 29776
rect 3016 29764 3022 29776
rect 3694 29764 3700 29776
rect 3016 29736 3700 29764
rect 3016 29724 3022 29736
rect 3694 29724 3700 29736
rect 3752 29724 3758 29776
rect 3786 29724 3792 29776
rect 3844 29764 3850 29776
rect 3844 29736 4108 29764
rect 3844 29724 3850 29736
rect 2406 29696 2412 29708
rect 2332 29668 2412 29696
rect 2406 29656 2412 29668
rect 2464 29656 2470 29708
rect 4080 29705 4108 29736
rect 4065 29699 4123 29705
rect 2746 29668 3832 29696
rect 1578 29588 1584 29640
rect 1636 29628 1642 29640
rect 1673 29631 1731 29637
rect 1673 29628 1685 29631
rect 1636 29600 1685 29628
rect 1636 29588 1642 29600
rect 1673 29597 1685 29600
rect 1719 29597 1731 29631
rect 1673 29591 1731 29597
rect 1947 29631 2005 29637
rect 1947 29597 1959 29631
rect 1993 29628 2005 29631
rect 2038 29628 2044 29640
rect 1993 29600 2044 29628
rect 1993 29597 2005 29600
rect 1947 29591 2005 29597
rect 2038 29588 2044 29600
rect 2096 29628 2102 29640
rect 2590 29628 2596 29640
rect 2096 29600 2596 29628
rect 2096 29588 2102 29600
rect 2590 29588 2596 29600
rect 2648 29588 2654 29640
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 2746 29560 2774 29668
rect 3804 29637 3832 29668
rect 4065 29665 4077 29699
rect 4111 29696 4123 29699
rect 4724 29696 4752 29792
rect 7576 29773 7604 29804
rect 7834 29792 7840 29804
rect 7892 29792 7898 29844
rect 8110 29792 8116 29844
rect 8168 29832 8174 29844
rect 8757 29835 8815 29841
rect 8168 29804 8524 29832
rect 8168 29792 8174 29804
rect 7561 29767 7619 29773
rect 7561 29733 7573 29767
rect 7607 29733 7619 29767
rect 8496 29764 8524 29804
rect 8757 29801 8769 29835
rect 8803 29832 8815 29835
rect 8846 29832 8852 29844
rect 8803 29804 8852 29832
rect 8803 29801 8815 29804
rect 8757 29795 8815 29801
rect 8846 29792 8852 29804
rect 8904 29792 8910 29844
rect 9030 29792 9036 29844
rect 9088 29832 9094 29844
rect 10870 29832 10876 29844
rect 9088 29804 10876 29832
rect 9088 29792 9094 29804
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 11072 29804 12112 29832
rect 11072 29764 11100 29804
rect 8496 29736 11100 29764
rect 7561 29727 7619 29733
rect 11146 29724 11152 29776
rect 11204 29724 11210 29776
rect 4111 29668 4752 29696
rect 4111 29665 4123 29668
rect 4065 29659 4123 29665
rect 5166 29656 5172 29708
rect 5224 29656 5230 29708
rect 7650 29696 7656 29708
rect 6840 29668 7656 29696
rect 3421 29631 3479 29637
rect 3421 29628 3433 29631
rect 3252 29600 3433 29628
rect 1360 29532 2774 29560
rect 1360 29520 1366 29532
rect 3142 29520 3148 29572
rect 3200 29520 3206 29572
rect 3252 29560 3280 29600
rect 3421 29597 3433 29600
rect 3467 29597 3479 29631
rect 3421 29591 3479 29597
rect 3789 29631 3847 29637
rect 3789 29597 3801 29631
rect 3835 29597 3847 29631
rect 3789 29591 3847 29597
rect 5261 29631 5319 29637
rect 5261 29597 5273 29631
rect 5307 29628 5319 29631
rect 6840 29628 6868 29668
rect 7650 29656 7656 29668
rect 7708 29656 7714 29708
rect 7834 29656 7840 29708
rect 7892 29656 7898 29708
rect 7975 29699 8033 29705
rect 7975 29665 7987 29699
rect 8021 29696 8033 29699
rect 8294 29696 8300 29708
rect 8021 29668 8300 29696
rect 8021 29665 8033 29668
rect 7975 29659 8033 29665
rect 8294 29656 8300 29668
rect 8352 29656 8358 29708
rect 9398 29656 9404 29708
rect 9456 29696 9462 29708
rect 10686 29696 10692 29708
rect 9456 29668 10692 29696
rect 9456 29656 9462 29668
rect 10686 29656 10692 29668
rect 10744 29656 10750 29708
rect 11054 29656 11060 29708
rect 11112 29696 11118 29708
rect 11606 29705 11612 29708
rect 11425 29699 11483 29705
rect 11425 29696 11437 29699
rect 11112 29668 11437 29696
rect 11112 29656 11118 29668
rect 11425 29665 11437 29668
rect 11471 29665 11483 29699
rect 11425 29659 11483 29665
rect 11563 29699 11612 29705
rect 11563 29665 11575 29699
rect 11609 29665 11612 29699
rect 11563 29659 11612 29665
rect 11606 29656 11612 29659
rect 11664 29656 11670 29708
rect 11701 29699 11759 29705
rect 11701 29665 11713 29699
rect 11747 29696 11759 29699
rect 11882 29696 11888 29708
rect 11747 29668 11888 29696
rect 11747 29665 11759 29668
rect 11701 29659 11759 29665
rect 11882 29656 11888 29668
rect 11940 29656 11946 29708
rect 12084 29696 12112 29804
rect 12342 29792 12348 29844
rect 12400 29792 12406 29844
rect 17405 29835 17463 29841
rect 17405 29801 17417 29835
rect 17451 29832 17463 29835
rect 17494 29832 17500 29844
rect 17451 29804 17500 29832
rect 17451 29801 17463 29804
rect 17405 29795 17463 29801
rect 17494 29792 17500 29804
rect 17552 29792 17558 29844
rect 17586 29792 17592 29844
rect 17644 29832 17650 29844
rect 20714 29832 20720 29844
rect 17644 29804 20720 29832
rect 17644 29792 17650 29804
rect 20714 29792 20720 29804
rect 20772 29792 20778 29844
rect 22830 29832 22836 29844
rect 22204 29804 22836 29832
rect 13449 29767 13507 29773
rect 13449 29733 13461 29767
rect 13495 29764 13507 29767
rect 13630 29764 13636 29776
rect 13495 29736 13636 29764
rect 13495 29733 13507 29736
rect 13449 29727 13507 29733
rect 13630 29724 13636 29736
rect 13688 29724 13694 29776
rect 16206 29724 16212 29776
rect 16264 29724 16270 29776
rect 12084 29668 12296 29696
rect 5307 29600 6868 29628
rect 6917 29631 6975 29637
rect 5307 29597 5319 29600
rect 5261 29591 5319 29597
rect 6917 29597 6929 29631
rect 6963 29597 6975 29631
rect 6917 29591 6975 29597
rect 5353 29563 5411 29569
rect 3252 29532 5120 29560
rect 3252 29504 3280 29532
rect 1670 29452 1676 29504
rect 1728 29492 1734 29504
rect 2222 29492 2228 29504
rect 1728 29464 2228 29492
rect 1728 29452 1734 29464
rect 2222 29452 2228 29464
rect 2280 29452 2286 29504
rect 2406 29452 2412 29504
rect 2464 29492 2470 29504
rect 2682 29492 2688 29504
rect 2464 29464 2688 29492
rect 2464 29452 2470 29464
rect 2682 29452 2688 29464
rect 2740 29452 2746 29504
rect 3234 29452 3240 29504
rect 3292 29452 3298 29504
rect 4982 29452 4988 29504
rect 5040 29452 5046 29504
rect 5092 29492 5120 29532
rect 5353 29529 5365 29563
rect 5399 29560 5411 29563
rect 5626 29560 5632 29572
rect 5399 29532 5632 29560
rect 5399 29529 5411 29532
rect 5353 29523 5411 29529
rect 5626 29520 5632 29532
rect 5684 29520 5690 29572
rect 5718 29520 5724 29572
rect 5776 29520 5782 29572
rect 5810 29520 5816 29572
rect 5868 29560 5874 29572
rect 5868 29532 6316 29560
rect 5868 29520 5874 29532
rect 6288 29501 6316 29532
rect 6089 29495 6147 29501
rect 6089 29492 6101 29495
rect 5092 29464 6101 29492
rect 6089 29461 6101 29464
rect 6135 29461 6147 29495
rect 6089 29455 6147 29461
rect 6273 29495 6331 29501
rect 6273 29461 6285 29495
rect 6319 29461 6331 29495
rect 6932 29492 6960 29591
rect 7098 29588 7104 29640
rect 7156 29588 7162 29640
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 10502 29588 10508 29640
rect 10560 29588 10566 29640
rect 9766 29560 9772 29572
rect 8588 29532 9772 29560
rect 7926 29492 7932 29504
rect 6932 29464 7932 29492
rect 6273 29455 6331 29461
rect 7926 29452 7932 29464
rect 7984 29452 7990 29504
rect 8386 29452 8392 29504
rect 8444 29492 8450 29504
rect 8588 29492 8616 29532
rect 9766 29520 9772 29532
rect 9824 29520 9830 29572
rect 8444 29464 8616 29492
rect 8444 29452 8450 29464
rect 8754 29452 8760 29504
rect 8812 29492 8818 29504
rect 12158 29492 12164 29504
rect 8812 29464 12164 29492
rect 8812 29452 8818 29464
rect 12158 29452 12164 29464
rect 12216 29452 12222 29504
rect 12268 29492 12296 29668
rect 13814 29656 13820 29708
rect 13872 29696 13878 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 13872 29668 14197 29696
rect 13872 29656 13878 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 14844 29668 15700 29696
rect 12342 29588 12348 29640
rect 12400 29618 12406 29640
rect 12437 29631 12495 29637
rect 12437 29618 12449 29631
rect 12400 29597 12449 29618
rect 12483 29597 12495 29631
rect 12710 29628 12716 29640
rect 12671 29600 12716 29628
rect 12400 29591 12495 29597
rect 12400 29590 12480 29591
rect 12400 29588 12406 29590
rect 12452 29560 12480 29590
rect 12710 29588 12716 29600
rect 12768 29588 12774 29640
rect 14427 29631 14485 29637
rect 14427 29628 14439 29631
rect 14200 29600 14439 29628
rect 14200 29572 14228 29600
rect 14427 29597 14439 29600
rect 14473 29597 14485 29631
rect 14844 29628 14872 29668
rect 14427 29591 14485 29597
rect 14752 29600 14872 29628
rect 15565 29631 15623 29637
rect 14752 29572 14780 29600
rect 15565 29597 15577 29631
rect 15611 29597 15623 29631
rect 15672 29628 15700 29668
rect 15746 29656 15752 29708
rect 15804 29656 15810 29708
rect 16485 29699 16543 29705
rect 16485 29696 16497 29699
rect 15856 29668 16497 29696
rect 15856 29628 15884 29668
rect 16485 29665 16497 29668
rect 16531 29665 16543 29699
rect 16485 29659 16543 29665
rect 16761 29699 16819 29705
rect 16761 29665 16773 29699
rect 16807 29696 16819 29699
rect 16942 29696 16948 29708
rect 16807 29668 16948 29696
rect 16807 29665 16819 29668
rect 16761 29659 16819 29665
rect 16942 29656 16948 29668
rect 17000 29656 17006 29708
rect 21729 29699 21787 29705
rect 21729 29665 21741 29699
rect 21775 29696 21787 29699
rect 22097 29699 22155 29705
rect 22097 29696 22109 29699
rect 21775 29668 22109 29696
rect 21775 29665 21787 29668
rect 21729 29659 21787 29665
rect 22097 29665 22109 29668
rect 22143 29665 22155 29699
rect 22097 29659 22155 29665
rect 15672 29600 15884 29628
rect 15565 29591 15623 29597
rect 12618 29560 12624 29572
rect 12452 29532 12624 29560
rect 12618 29520 12624 29532
rect 12676 29520 12682 29572
rect 13538 29520 13544 29572
rect 13596 29560 13602 29572
rect 14182 29560 14188 29572
rect 13596 29532 14188 29560
rect 13596 29520 13602 29532
rect 14182 29520 14188 29532
rect 14240 29520 14246 29572
rect 14734 29520 14740 29572
rect 14792 29520 14798 29572
rect 15102 29492 15108 29504
rect 12268 29464 15108 29492
rect 15102 29452 15108 29464
rect 15160 29452 15166 29504
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 15580 29492 15608 29591
rect 16574 29588 16580 29640
rect 16632 29637 16638 29640
rect 16632 29631 16660 29637
rect 16648 29597 16660 29631
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 16632 29591 16660 29597
rect 20916 29600 21189 29628
rect 16632 29588 16638 29591
rect 19242 29520 19248 29572
rect 19300 29560 19306 29572
rect 20530 29560 20536 29572
rect 19300 29532 20536 29560
rect 19300 29520 19306 29532
rect 20530 29520 20536 29532
rect 20588 29560 20594 29572
rect 20916 29560 20944 29600
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21637 29631 21695 29637
rect 21637 29597 21649 29631
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 22005 29631 22063 29637
rect 22005 29597 22017 29631
rect 22051 29628 22063 29631
rect 22204 29628 22232 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 23198 29792 23204 29844
rect 23256 29832 23262 29844
rect 23256 29804 23704 29832
rect 23256 29792 23262 29804
rect 23293 29767 23351 29773
rect 23293 29733 23305 29767
rect 23339 29733 23351 29767
rect 23293 29727 23351 29733
rect 23569 29767 23627 29773
rect 23569 29733 23581 29767
rect 23615 29733 23627 29767
rect 23569 29727 23627 29733
rect 22281 29699 22339 29705
rect 22281 29665 22293 29699
rect 22327 29696 22339 29699
rect 22465 29699 22523 29705
rect 22465 29696 22477 29699
rect 22327 29668 22477 29696
rect 22327 29665 22339 29668
rect 22281 29659 22339 29665
rect 22465 29665 22477 29668
rect 22511 29665 22523 29699
rect 22465 29659 22523 29665
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22051 29600 22385 29628
rect 22051 29597 22063 29600
rect 22005 29591 22063 29597
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 21652 29560 21680 29591
rect 22554 29588 22560 29640
rect 22612 29588 22618 29640
rect 20588 29532 20944 29560
rect 21008 29532 21680 29560
rect 22281 29563 22339 29569
rect 20588 29520 20594 29532
rect 16666 29492 16672 29504
rect 15580 29464 16672 29492
rect 16666 29452 16672 29464
rect 16724 29492 16730 29504
rect 17034 29492 17040 29504
rect 16724 29464 17040 29492
rect 16724 29452 16730 29464
rect 17034 29452 17040 29464
rect 17092 29452 17098 29504
rect 17862 29452 17868 29504
rect 17920 29492 17926 29504
rect 19978 29492 19984 29504
rect 17920 29464 19984 29492
rect 17920 29452 17926 29464
rect 19978 29452 19984 29464
rect 20036 29452 20042 29504
rect 21008 29501 21036 29532
rect 22281 29529 22293 29563
rect 22327 29529 22339 29563
rect 23308 29560 23336 29727
rect 23477 29631 23535 29637
rect 23477 29597 23489 29631
rect 23523 29628 23535 29631
rect 23584 29628 23612 29727
rect 23523 29600 23612 29628
rect 23676 29628 23704 29804
rect 23753 29631 23811 29637
rect 23753 29628 23765 29631
rect 23676 29600 23765 29628
rect 23523 29597 23535 29600
rect 23477 29591 23535 29597
rect 23753 29597 23765 29600
rect 23799 29597 23811 29631
rect 23753 29591 23811 29597
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29597 23995 29631
rect 23937 29591 23995 29597
rect 23952 29560 23980 29591
rect 24210 29560 24216 29572
rect 23308 29532 23980 29560
rect 24044 29532 24216 29560
rect 22281 29523 22339 29529
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29461 21051 29495
rect 22296 29492 22324 29523
rect 24044 29492 24072 29532
rect 24210 29520 24216 29532
rect 24268 29520 24274 29572
rect 22296 29464 24072 29492
rect 24121 29495 24179 29501
rect 20993 29455 21051 29461
rect 24121 29461 24133 29495
rect 24167 29492 24179 29495
rect 25130 29492 25136 29504
rect 24167 29464 25136 29492
rect 24167 29461 24179 29464
rect 24121 29455 24179 29461
rect 25130 29452 25136 29464
rect 25188 29452 25194 29504
rect 198 29384 204 29436
rect 256 29424 262 29436
rect 566 29424 572 29436
rect 256 29396 572 29424
rect 256 29384 262 29396
rect 566 29384 572 29396
rect 624 29384 630 29436
rect 1104 29402 25000 29424
rect 1104 29350 6884 29402
rect 6936 29350 6948 29402
rect 7000 29350 7012 29402
rect 7064 29350 7076 29402
rect 7128 29350 7140 29402
rect 7192 29350 12818 29402
rect 12870 29350 12882 29402
rect 12934 29350 12946 29402
rect 12998 29350 13010 29402
rect 13062 29350 13074 29402
rect 13126 29350 18752 29402
rect 18804 29350 18816 29402
rect 18868 29350 18880 29402
rect 18932 29350 18944 29402
rect 18996 29350 19008 29402
rect 19060 29350 24686 29402
rect 24738 29350 24750 29402
rect 24802 29350 24814 29402
rect 24866 29350 24878 29402
rect 24930 29350 24942 29402
rect 24994 29350 25000 29402
rect 1104 29328 25000 29350
rect 658 29248 664 29300
rect 716 29288 722 29300
rect 4522 29288 4528 29300
rect 716 29260 4528 29288
rect 716 29248 722 29260
rect 4522 29248 4528 29260
rect 4580 29248 4586 29300
rect 5000 29260 5580 29288
rect 5000 29232 5028 29260
rect 934 29180 940 29232
rect 992 29220 998 29232
rect 1857 29223 1915 29229
rect 1857 29220 1869 29223
rect 992 29192 1869 29220
rect 992 29180 998 29192
rect 1857 29189 1869 29192
rect 1903 29189 1915 29223
rect 1857 29183 1915 29189
rect 1946 29180 1952 29232
rect 2004 29180 2010 29232
rect 2041 29223 2099 29229
rect 2041 29189 2053 29223
rect 2087 29220 2099 29223
rect 2087 29192 4936 29220
rect 2087 29189 2099 29192
rect 2041 29183 2099 29189
rect 1486 29112 1492 29164
rect 1544 29112 1550 29164
rect 1964 29152 1992 29180
rect 2467 29155 2525 29161
rect 2467 29152 2479 29155
rect 1964 29124 2479 29152
rect 2467 29121 2479 29124
rect 2513 29152 2525 29155
rect 2866 29152 2872 29164
rect 2513 29124 2872 29152
rect 2513 29121 2525 29124
rect 2467 29115 2525 29121
rect 2866 29112 2872 29124
rect 2924 29112 2930 29164
rect 3602 29112 3608 29164
rect 3660 29112 3666 29164
rect 4908 29152 4936 29192
rect 4982 29180 4988 29232
rect 5040 29180 5046 29232
rect 5552 29220 5580 29260
rect 5626 29248 5632 29300
rect 5684 29288 5690 29300
rect 5905 29291 5963 29297
rect 5905 29288 5917 29291
rect 5684 29260 5917 29288
rect 5684 29248 5690 29260
rect 5905 29257 5917 29260
rect 5951 29257 5963 29291
rect 5905 29251 5963 29257
rect 8110 29248 8116 29300
rect 8168 29288 8174 29300
rect 8389 29291 8447 29297
rect 8389 29288 8401 29291
rect 8168 29260 8401 29288
rect 8168 29248 8174 29260
rect 8389 29257 8401 29260
rect 8435 29257 8447 29291
rect 8389 29251 8447 29257
rect 8570 29248 8576 29300
rect 8628 29288 8634 29300
rect 8846 29288 8852 29300
rect 8628 29260 8852 29288
rect 8628 29248 8634 29260
rect 8846 29248 8852 29260
rect 8904 29248 8910 29300
rect 9382 29260 9674 29288
rect 9382 29220 9410 29260
rect 5092 29192 5488 29220
rect 5552 29192 9410 29220
rect 9646 29220 9674 29260
rect 10686 29248 10692 29300
rect 10744 29288 10750 29300
rect 10873 29291 10931 29297
rect 10873 29288 10885 29291
rect 10744 29260 10885 29288
rect 10744 29248 10750 29260
rect 10873 29257 10885 29260
rect 10919 29257 10931 29291
rect 10873 29251 10931 29257
rect 11238 29248 11244 29300
rect 11296 29288 11302 29300
rect 11701 29291 11759 29297
rect 11701 29288 11713 29291
rect 11296 29260 11713 29288
rect 11296 29248 11302 29260
rect 11701 29257 11713 29260
rect 11747 29257 11759 29291
rect 11701 29251 11759 29257
rect 13722 29248 13728 29300
rect 13780 29288 13786 29300
rect 14277 29291 14335 29297
rect 14277 29288 14289 29291
rect 13780 29260 14289 29288
rect 13780 29248 13786 29260
rect 14277 29257 14289 29260
rect 14323 29257 14335 29291
rect 23109 29291 23167 29297
rect 14277 29251 14335 29257
rect 14366 29260 22094 29288
rect 11609 29223 11667 29229
rect 11609 29220 11621 29223
rect 9646 29192 11621 29220
rect 5092 29152 5120 29192
rect 4908 29124 5120 29152
rect 5166 29112 5172 29164
rect 5224 29152 5230 29164
rect 5460 29152 5488 29192
rect 11609 29189 11621 29192
rect 11655 29220 11667 29223
rect 13354 29220 13360 29232
rect 11655 29192 13360 29220
rect 11655 29189 11667 29192
rect 11609 29183 11667 29189
rect 13354 29180 13360 29192
rect 13412 29180 13418 29232
rect 9459 29165 9517 29171
rect 9459 29164 9471 29165
rect 5224 29124 5267 29152
rect 5460 29124 6408 29152
rect 5224 29112 5230 29124
rect 1673 29087 1731 29093
rect 1673 29053 1685 29087
rect 1719 29084 1731 29087
rect 1719 29056 1992 29084
rect 1719 29053 1731 29056
rect 1673 29047 1731 29053
rect 1964 29028 1992 29056
rect 2130 29044 2136 29096
rect 2188 29084 2194 29096
rect 2225 29087 2283 29093
rect 2225 29084 2237 29087
rect 2188 29056 2237 29084
rect 2188 29044 2194 29056
rect 2225 29053 2237 29056
rect 2271 29053 2283 29087
rect 2225 29047 2283 29053
rect 4890 29044 4896 29096
rect 4948 29044 4954 29096
rect 6380 29084 6408 29124
rect 6454 29112 6460 29164
rect 6512 29152 6518 29164
rect 7190 29152 7196 29164
rect 6512 29124 7196 29152
rect 6512 29112 6518 29124
rect 7190 29112 7196 29124
rect 7248 29156 7254 29164
rect 7377 29156 7435 29161
rect 7248 29155 7435 29156
rect 7248 29128 7389 29155
rect 7248 29112 7254 29128
rect 7377 29121 7389 29128
rect 7423 29121 7435 29155
rect 7650 29152 7656 29164
rect 7611 29124 7656 29152
rect 7377 29115 7435 29121
rect 7650 29112 7656 29124
rect 7708 29112 7714 29164
rect 8754 29112 8760 29164
rect 8812 29152 8818 29164
rect 9398 29162 9404 29164
rect 9217 29155 9275 29161
rect 9217 29152 9229 29155
rect 8812 29124 9229 29152
rect 8812 29112 8818 29124
rect 9217 29121 9229 29124
rect 9263 29121 9275 29155
rect 9382 29124 9404 29162
rect 9217 29115 9275 29121
rect 9398 29112 9404 29124
rect 9456 29131 9471 29164
rect 9505 29131 9517 29165
rect 9456 29125 9517 29131
rect 10597 29155 10655 29161
rect 9456 29112 9462 29125
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 11330 29152 11336 29164
rect 10643 29124 11336 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 6380 29056 7420 29084
rect 1946 28976 1952 29028
rect 2004 28976 2010 29028
rect 3234 28976 3240 29028
rect 3292 28976 3298 29028
rect 3789 29019 3847 29025
rect 3789 28985 3801 29019
rect 3835 29016 3847 29019
rect 7098 29016 7104 29028
rect 3835 28988 5028 29016
rect 3835 28985 3847 28988
rect 3789 28979 3847 28985
rect 5000 28948 5028 28988
rect 5552 28988 7104 29016
rect 5552 28948 5580 28988
rect 7098 28976 7104 28988
rect 7156 28976 7162 29028
rect 7392 29016 7420 29056
rect 8570 29044 8576 29096
rect 8628 29044 8634 29096
rect 8588 29016 8616 29044
rect 7392 28988 7512 29016
rect 5000 28920 5580 28948
rect 7484 28948 7512 28988
rect 8036 28988 8616 29016
rect 10229 29019 10287 29025
rect 8036 28948 8064 28988
rect 10229 28985 10241 29019
rect 10275 29016 10287 29019
rect 10612 29016 10640 29115
rect 11330 29112 11336 29124
rect 11388 29112 11394 29164
rect 12066 29112 12072 29164
rect 12124 29152 12130 29164
rect 12803 29155 12861 29161
rect 12803 29152 12815 29155
rect 12124 29124 12815 29152
rect 12124 29112 12130 29124
rect 12803 29121 12815 29124
rect 12849 29152 12861 29155
rect 14366 29152 14394 29260
rect 14645 29223 14703 29229
rect 14645 29189 14657 29223
rect 14691 29220 14703 29223
rect 15194 29220 15200 29232
rect 14691 29192 15200 29220
rect 14691 29189 14703 29192
rect 14645 29183 14703 29189
rect 15194 29180 15200 29192
rect 15252 29180 15258 29232
rect 15381 29223 15439 29229
rect 15381 29189 15393 29223
rect 15427 29189 15439 29223
rect 15381 29183 15439 29189
rect 12849 29124 14394 29152
rect 14553 29155 14611 29161
rect 12849 29121 12861 29124
rect 12803 29115 12861 29121
rect 14553 29121 14565 29155
rect 14599 29152 14611 29155
rect 14734 29152 14740 29164
rect 14599 29124 14740 29152
rect 14599 29121 14611 29124
rect 14553 29115 14611 29121
rect 14734 29112 14740 29124
rect 14792 29112 14798 29164
rect 15013 29155 15071 29161
rect 15013 29121 15025 29155
rect 15059 29152 15071 29155
rect 15102 29152 15108 29164
rect 15059 29124 15108 29152
rect 15059 29121 15071 29124
rect 15013 29115 15071 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 15396 29152 15424 29183
rect 16574 29180 16580 29232
rect 16632 29220 16638 29232
rect 17586 29220 17592 29232
rect 16632 29192 17592 29220
rect 16632 29180 16638 29192
rect 17586 29180 17592 29192
rect 17644 29180 17650 29232
rect 19150 29191 19156 29232
rect 19135 29185 19156 29191
rect 15562 29152 15568 29164
rect 15396 29124 15568 29152
rect 15562 29112 15568 29124
rect 15620 29112 15626 29164
rect 16942 29152 16948 29164
rect 16903 29124 16948 29152
rect 16942 29112 16948 29124
rect 17000 29112 17006 29164
rect 17862 29112 17868 29164
rect 17920 29152 17926 29164
rect 18877 29155 18935 29161
rect 18877 29152 18889 29155
rect 17920 29124 18889 29152
rect 17920 29112 17926 29124
rect 18877 29121 18889 29124
rect 18923 29121 18935 29155
rect 19135 29151 19147 29185
rect 19208 29180 19214 29232
rect 19518 29180 19524 29232
rect 19576 29220 19582 29232
rect 19576 29192 20484 29220
rect 19576 29180 19582 29192
rect 19181 29154 19196 29180
rect 20456 29161 20484 29192
rect 20257 29155 20315 29161
rect 19181 29151 19193 29154
rect 20257 29152 20269 29155
rect 19135 29145 19193 29151
rect 18877 29115 18935 29121
rect 19904 29124 20269 29152
rect 10873 29087 10931 29093
rect 10873 29053 10885 29087
rect 10919 29084 10931 29087
rect 10919 29056 11468 29084
rect 10919 29053 10931 29056
rect 10873 29047 10931 29053
rect 10275 28988 10640 29016
rect 10689 29019 10747 29025
rect 10275 28985 10287 28988
rect 10229 28979 10287 28985
rect 10689 28985 10701 29019
rect 10735 29016 10747 29019
rect 11146 29016 11152 29028
rect 10735 28988 11152 29016
rect 10735 28985 10747 28988
rect 10689 28979 10747 28985
rect 11146 28976 11152 28988
rect 11204 28976 11210 29028
rect 11440 28960 11468 29056
rect 12526 29044 12532 29096
rect 12584 29044 12590 29096
rect 13446 29044 13452 29096
rect 13504 29084 13510 29096
rect 13630 29084 13636 29096
rect 13504 29056 13636 29084
rect 13504 29044 13510 29056
rect 13630 29044 13636 29056
rect 13688 29044 13694 29096
rect 14918 29044 14924 29096
rect 14976 29044 14982 29096
rect 16666 29044 16672 29096
rect 16724 29044 16730 29096
rect 12544 29016 12572 29044
rect 12544 28988 12664 29016
rect 7484 28920 8064 28948
rect 8110 28908 8116 28960
rect 8168 28948 8174 28960
rect 11054 28948 11060 28960
rect 8168 28920 11060 28948
rect 8168 28908 8174 28920
rect 11054 28908 11060 28920
rect 11112 28908 11118 28960
rect 11422 28908 11428 28960
rect 11480 28908 11486 28960
rect 12636 28948 12664 28988
rect 13188 28988 14136 29016
rect 13188 28948 13216 28988
rect 14108 28960 14136 28988
rect 15470 28976 15476 29028
rect 15528 29016 15534 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 15528 28988 15577 29016
rect 15528 28976 15534 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 19794 29016 19800 29028
rect 15565 28979 15623 28985
rect 19536 28988 19800 29016
rect 12636 28920 13216 28948
rect 13541 28951 13599 28957
rect 13541 28917 13553 28951
rect 13587 28948 13599 28951
rect 13722 28948 13728 28960
rect 13587 28920 13728 28948
rect 13587 28917 13599 28920
rect 13541 28911 13599 28917
rect 13722 28908 13728 28920
rect 13780 28908 13786 28960
rect 14090 28908 14096 28960
rect 14148 28908 14154 28960
rect 17126 28908 17132 28960
rect 17184 28948 17190 28960
rect 17681 28951 17739 28957
rect 17681 28948 17693 28951
rect 17184 28920 17693 28948
rect 17184 28908 17190 28920
rect 17681 28917 17693 28920
rect 17727 28917 17739 28951
rect 17681 28911 17739 28917
rect 17862 28908 17868 28960
rect 17920 28948 17926 28960
rect 19536 28948 19564 28988
rect 19794 28976 19800 28988
rect 19852 28976 19858 29028
rect 17920 28920 19564 28948
rect 17920 28908 17926 28920
rect 19610 28908 19616 28960
rect 19668 28948 19674 28960
rect 19904 28957 19932 29124
rect 20257 29121 20269 29124
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 22066 29152 22094 29260
rect 23109 29257 23121 29291
rect 23155 29257 23167 29291
rect 23109 29251 23167 29257
rect 23124 29220 23152 29251
rect 23124 29192 23888 29220
rect 23860 29161 23888 29192
rect 23293 29155 23351 29161
rect 23293 29152 23305 29155
rect 22066 29124 23305 29152
rect 20441 29115 20499 29121
rect 23293 29121 23305 29124
rect 23339 29121 23351 29155
rect 23293 29115 23351 29121
rect 23569 29155 23627 29161
rect 23569 29121 23581 29155
rect 23615 29121 23627 29155
rect 23569 29115 23627 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29121 23903 29155
rect 23845 29115 23903 29121
rect 24121 29155 24179 29161
rect 24121 29121 24133 29155
rect 24167 29121 24179 29155
rect 24121 29115 24179 29121
rect 23385 29019 23443 29025
rect 20272 28988 20484 29016
rect 20272 28960 20300 28988
rect 19889 28951 19947 28957
rect 19889 28948 19901 28951
rect 19668 28920 19901 28948
rect 19668 28908 19674 28920
rect 19889 28917 19901 28920
rect 19935 28917 19947 28951
rect 19889 28911 19947 28917
rect 20254 28908 20260 28960
rect 20312 28908 20318 28960
rect 20346 28908 20352 28960
rect 20404 28908 20410 28960
rect 20456 28948 20484 28988
rect 23385 28985 23397 29019
rect 23431 29016 23443 29019
rect 23584 29016 23612 29115
rect 24136 29084 24164 29115
rect 23768 29056 24164 29084
rect 23661 29019 23719 29025
rect 23661 29016 23673 29019
rect 23431 28988 23520 29016
rect 23584 28988 23673 29016
rect 23431 28985 23443 28988
rect 23385 28979 23443 28985
rect 22738 28948 22744 28960
rect 20456 28920 22744 28948
rect 22738 28908 22744 28920
rect 22796 28908 22802 28960
rect 23492 28948 23520 28988
rect 23661 28985 23673 28988
rect 23707 28985 23719 29019
rect 23661 28979 23719 28985
rect 23768 28948 23796 29056
rect 23492 28920 23796 28948
rect 24394 28908 24400 28960
rect 24452 28908 24458 28960
rect 1104 28858 24840 28880
rect 1104 28806 3917 28858
rect 3969 28806 3981 28858
rect 4033 28806 4045 28858
rect 4097 28806 4109 28858
rect 4161 28806 4173 28858
rect 4225 28806 9851 28858
rect 9903 28806 9915 28858
rect 9967 28806 9979 28858
rect 10031 28806 10043 28858
rect 10095 28806 10107 28858
rect 10159 28806 15785 28858
rect 15837 28806 15849 28858
rect 15901 28806 15913 28858
rect 15965 28806 15977 28858
rect 16029 28806 16041 28858
rect 16093 28806 21719 28858
rect 21771 28806 21783 28858
rect 21835 28806 21847 28858
rect 21899 28806 21911 28858
rect 21963 28806 21975 28858
rect 22027 28806 24840 28858
rect 1104 28784 24840 28806
rect 1578 28704 1584 28756
rect 1636 28744 1642 28756
rect 1854 28744 1860 28756
rect 1636 28716 1860 28744
rect 1636 28704 1642 28716
rect 1854 28704 1860 28716
rect 1912 28704 1918 28756
rect 2225 28747 2283 28753
rect 2225 28713 2237 28747
rect 2271 28744 2283 28747
rect 2271 28716 10916 28744
rect 2271 28713 2283 28716
rect 2225 28707 2283 28713
rect 10505 28679 10563 28685
rect 10505 28645 10517 28679
rect 10551 28645 10563 28679
rect 10505 28639 10563 28645
rect 10781 28679 10839 28685
rect 10781 28645 10793 28679
rect 10827 28645 10839 28679
rect 10888 28676 10916 28716
rect 11146 28704 11152 28756
rect 11204 28704 11210 28756
rect 11422 28704 11428 28756
rect 11480 28704 11486 28756
rect 11606 28704 11612 28756
rect 11664 28704 11670 28756
rect 18877 28747 18935 28753
rect 16408 28716 18552 28744
rect 11624 28676 11652 28704
rect 10888 28648 11652 28676
rect 10781 28639 10839 28645
rect 2130 28568 2136 28620
rect 2188 28608 2194 28620
rect 2317 28611 2375 28617
rect 2317 28608 2329 28611
rect 2188 28580 2329 28608
rect 2188 28568 2194 28580
rect 2317 28577 2329 28580
rect 2363 28577 2375 28611
rect 8110 28608 8116 28620
rect 2317 28571 2375 28577
rect 4540 28580 8116 28608
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 2038 28500 2044 28552
rect 2096 28500 2102 28552
rect 2590 28540 2596 28552
rect 2551 28512 2596 28540
rect 2590 28500 2596 28512
rect 2648 28500 2654 28552
rect 3786 28500 3792 28552
rect 3844 28540 3850 28552
rect 3881 28543 3939 28549
rect 3881 28540 3893 28543
rect 3844 28512 3893 28540
rect 3844 28500 3850 28512
rect 3881 28509 3893 28512
rect 3927 28509 3939 28543
rect 4154 28540 4160 28552
rect 4115 28512 4160 28540
rect 3881 28503 3939 28509
rect 4154 28500 4160 28512
rect 4212 28500 4218 28552
rect 750 28432 756 28484
rect 808 28472 814 28484
rect 1489 28475 1547 28481
rect 1489 28472 1501 28475
rect 808 28444 1501 28472
rect 808 28432 814 28444
rect 1489 28441 1501 28444
rect 1535 28441 1547 28475
rect 1489 28435 1547 28441
rect 1670 28432 1676 28484
rect 1728 28472 1734 28484
rect 4540 28472 4568 28580
rect 8110 28568 8116 28580
rect 8168 28568 8174 28620
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 7742 28540 7748 28552
rect 7248 28512 7748 28540
rect 7248 28500 7254 28512
rect 7742 28500 7748 28512
rect 7800 28540 7806 28552
rect 8941 28543 8999 28549
rect 8941 28540 8953 28543
rect 7800 28512 8953 28540
rect 7800 28500 7806 28512
rect 8941 28509 8953 28512
rect 8987 28509 8999 28543
rect 9214 28540 9220 28552
rect 9175 28512 9220 28540
rect 8941 28503 8999 28509
rect 9214 28500 9220 28512
rect 9272 28540 9278 28552
rect 9582 28540 9588 28552
rect 9272 28512 9588 28540
rect 9272 28500 9278 28512
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 1728 28444 4568 28472
rect 1728 28432 1734 28444
rect 5258 28432 5264 28484
rect 5316 28472 5322 28484
rect 10410 28472 10416 28484
rect 5316 28444 10416 28472
rect 5316 28432 5322 28444
rect 10410 28432 10416 28444
rect 10468 28432 10474 28484
rect 10520 28472 10548 28639
rect 10796 28608 10824 28639
rect 16408 28608 16436 28716
rect 18417 28679 18475 28685
rect 18417 28645 18429 28679
rect 18463 28645 18475 28679
rect 18524 28676 18552 28716
rect 18877 28713 18889 28747
rect 18923 28744 18935 28747
rect 19518 28744 19524 28756
rect 18923 28716 19524 28744
rect 18923 28713 18935 28716
rect 18877 28707 18935 28713
rect 19518 28704 19524 28716
rect 19576 28704 19582 28756
rect 20346 28744 20352 28756
rect 19996 28716 20352 28744
rect 19426 28676 19432 28688
rect 18524 28648 19432 28676
rect 18417 28639 18475 28645
rect 10796 28580 11560 28608
rect 10686 28500 10692 28552
rect 10744 28500 10750 28552
rect 10962 28500 10968 28552
rect 11020 28500 11026 28552
rect 11057 28543 11115 28549
rect 11057 28509 11069 28543
rect 11103 28509 11115 28543
rect 11057 28503 11115 28509
rect 11072 28472 11100 28503
rect 11330 28500 11336 28552
rect 11388 28500 11394 28552
rect 11532 28549 11560 28580
rect 15212 28580 16436 28608
rect 11517 28543 11575 28549
rect 11517 28509 11529 28543
rect 11563 28509 11575 28543
rect 11517 28503 11575 28509
rect 11698 28500 11704 28552
rect 11756 28500 11762 28552
rect 11882 28500 11888 28552
rect 11940 28540 11946 28552
rect 11975 28543 12033 28549
rect 11975 28540 11987 28543
rect 11940 28512 11987 28540
rect 11940 28500 11946 28512
rect 11975 28509 11987 28512
rect 12021 28540 12033 28543
rect 13814 28540 13820 28552
rect 12021 28512 13820 28540
rect 12021 28509 12033 28512
rect 11975 28503 12033 28509
rect 13814 28500 13820 28512
rect 13872 28500 13878 28552
rect 14090 28500 14096 28552
rect 14148 28500 14154 28552
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 15212 28540 15240 28580
rect 16666 28568 16672 28620
rect 16724 28568 16730 28620
rect 16942 28568 16948 28620
rect 17000 28568 17006 28620
rect 17218 28568 17224 28620
rect 17276 28568 17282 28620
rect 18432 28608 18460 28639
rect 19426 28636 19432 28648
rect 19484 28636 19490 28688
rect 19337 28611 19395 28617
rect 18432 28580 19288 28608
rect 14424 28512 15240 28540
rect 14424 28500 14430 28512
rect 15286 28500 15292 28552
rect 15344 28540 15350 28552
rect 16025 28543 16083 28549
rect 16025 28540 16037 28543
rect 15344 28512 16037 28540
rect 15344 28500 15350 28512
rect 16025 28509 16037 28512
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 16114 28500 16120 28552
rect 16172 28540 16178 28552
rect 16209 28543 16267 28549
rect 16209 28540 16221 28543
rect 16172 28512 16221 28540
rect 16172 28500 16178 28512
rect 16209 28509 16221 28512
rect 16255 28509 16267 28543
rect 16209 28503 16267 28509
rect 17034 28500 17040 28552
rect 17092 28549 17098 28552
rect 17092 28543 17120 28549
rect 17108 28509 17120 28543
rect 17092 28503 17120 28509
rect 17865 28543 17923 28549
rect 17865 28509 17877 28543
rect 17911 28540 17923 28543
rect 17954 28540 17960 28552
rect 17911 28512 17960 28540
rect 17911 28509 17923 28512
rect 17865 28503 17923 28509
rect 17092 28500 17098 28503
rect 17954 28500 17960 28512
rect 18012 28540 18018 28552
rect 18601 28543 18659 28549
rect 18601 28540 18613 28543
rect 18012 28512 18613 28540
rect 18012 28500 18018 28512
rect 18601 28509 18613 28512
rect 18647 28509 18659 28543
rect 18601 28503 18659 28509
rect 18690 28500 18696 28552
rect 18748 28540 18754 28552
rect 19260 28549 19288 28580
rect 19337 28577 19349 28611
rect 19383 28608 19395 28611
rect 19705 28611 19763 28617
rect 19705 28608 19717 28611
rect 19383 28580 19717 28608
rect 19383 28577 19395 28580
rect 19337 28571 19395 28577
rect 19705 28577 19717 28580
rect 19751 28577 19763 28611
rect 19705 28571 19763 28577
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28608 19947 28611
rect 19996 28608 20024 28716
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 23477 28747 23535 28753
rect 23477 28744 23489 28747
rect 23124 28716 23489 28744
rect 19935 28580 20024 28608
rect 19935 28577 19947 28580
rect 19889 28571 19947 28577
rect 19061 28543 19119 28549
rect 19061 28540 19073 28543
rect 18748 28512 19073 28540
rect 18748 28500 18754 28512
rect 19061 28509 19073 28512
rect 19107 28509 19119 28543
rect 19061 28503 19119 28509
rect 19245 28543 19303 28549
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 19610 28500 19616 28552
rect 19668 28500 19674 28552
rect 19978 28500 19984 28552
rect 20036 28500 20042 28552
rect 20255 28543 20313 28549
rect 20255 28509 20267 28543
rect 20301 28540 20313 28543
rect 20346 28540 20352 28552
rect 20301 28512 20352 28540
rect 20301 28509 20313 28512
rect 20255 28503 20313 28509
rect 20346 28500 20352 28512
rect 20404 28500 20410 28552
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 22066 28512 22845 28540
rect 22066 28472 22094 28512
rect 22833 28509 22845 28512
rect 22879 28509 22891 28543
rect 23124 28540 23152 28716
rect 23477 28713 23489 28716
rect 23523 28713 23535 28747
rect 23477 28707 23535 28713
rect 23201 28679 23259 28685
rect 23201 28645 23213 28679
rect 23247 28645 23259 28679
rect 23201 28639 23259 28645
rect 23216 28608 23244 28639
rect 23216 28580 23980 28608
rect 23952 28549 23980 28580
rect 23385 28543 23443 28549
rect 23385 28540 23397 28543
rect 23124 28512 23397 28540
rect 22833 28503 22891 28509
rect 23385 28509 23397 28512
rect 23431 28509 23443 28543
rect 23385 28503 23443 28509
rect 23661 28543 23719 28549
rect 23661 28509 23673 28543
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28509 23995 28543
rect 23937 28503 23995 28509
rect 23676 28472 23704 28503
rect 10520 28444 11100 28472
rect 11164 28444 15238 28472
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 1946 28364 1952 28416
rect 2004 28364 2010 28416
rect 3326 28364 3332 28416
rect 3384 28364 3390 28416
rect 4893 28407 4951 28413
rect 4893 28373 4905 28407
rect 4939 28404 4951 28407
rect 4982 28404 4988 28416
rect 4939 28376 4988 28404
rect 4939 28373 4951 28376
rect 4893 28367 4951 28373
rect 4982 28364 4988 28376
rect 5040 28364 5046 28416
rect 5166 28364 5172 28416
rect 5224 28404 5230 28416
rect 5442 28404 5448 28416
rect 5224 28376 5448 28404
rect 5224 28364 5230 28376
rect 5442 28364 5448 28376
rect 5500 28364 5506 28416
rect 6546 28364 6552 28416
rect 6604 28404 6610 28416
rect 7282 28404 7288 28416
rect 6604 28376 7288 28404
rect 6604 28364 6610 28376
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 9030 28364 9036 28416
rect 9088 28404 9094 28416
rect 9214 28404 9220 28416
rect 9088 28376 9220 28404
rect 9088 28364 9094 28376
rect 9214 28364 9220 28376
rect 9272 28364 9278 28416
rect 9674 28364 9680 28416
rect 9732 28404 9738 28416
rect 9953 28407 10011 28413
rect 9953 28404 9965 28407
rect 9732 28376 9965 28404
rect 9732 28364 9738 28376
rect 9953 28373 9965 28376
rect 9999 28373 10011 28407
rect 9953 28367 10011 28373
rect 10042 28364 10048 28416
rect 10100 28404 10106 28416
rect 11164 28404 11192 28444
rect 10100 28376 11192 28404
rect 10100 28364 10106 28376
rect 11882 28364 11888 28416
rect 11940 28404 11946 28416
rect 12713 28407 12771 28413
rect 12713 28404 12725 28407
rect 11940 28376 12725 28404
rect 11940 28364 11946 28376
rect 12713 28373 12725 28376
rect 12759 28373 12771 28407
rect 12713 28367 12771 28373
rect 13170 28364 13176 28416
rect 13228 28404 13234 28416
rect 13906 28404 13912 28416
rect 13228 28376 13912 28404
rect 13228 28364 13234 28376
rect 13906 28364 13912 28376
rect 13964 28364 13970 28416
rect 13998 28364 14004 28416
rect 14056 28404 14062 28416
rect 14274 28404 14280 28416
rect 14056 28376 14280 28404
rect 14056 28364 14062 28376
rect 14274 28364 14280 28376
rect 14332 28404 14338 28416
rect 15105 28407 15163 28413
rect 15105 28404 15117 28407
rect 14332 28376 15117 28404
rect 14332 28364 14338 28376
rect 15105 28373 15117 28376
rect 15151 28373 15163 28407
rect 15210 28404 15238 28444
rect 19306 28444 22094 28472
rect 22664 28444 23704 28472
rect 19306 28404 19334 28444
rect 15210 28376 19334 28404
rect 19889 28407 19947 28413
rect 15105 28367 15163 28373
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 20530 28404 20536 28416
rect 19935 28376 20536 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 20530 28364 20536 28376
rect 20588 28364 20594 28416
rect 20990 28364 20996 28416
rect 21048 28364 21054 28416
rect 22664 28413 22692 28444
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28373 22707 28407
rect 22649 28367 22707 28373
rect 24121 28407 24179 28413
rect 24121 28373 24133 28407
rect 24167 28404 24179 28407
rect 25130 28404 25136 28416
rect 24167 28376 25136 28404
rect 24167 28373 24179 28376
rect 24121 28367 24179 28373
rect 25130 28364 25136 28376
rect 25188 28364 25194 28416
rect 1104 28314 25000 28336
rect 1104 28262 6884 28314
rect 6936 28262 6948 28314
rect 7000 28262 7012 28314
rect 7064 28262 7076 28314
rect 7128 28262 7140 28314
rect 7192 28262 12818 28314
rect 12870 28262 12882 28314
rect 12934 28262 12946 28314
rect 12998 28262 13010 28314
rect 13062 28262 13074 28314
rect 13126 28262 18752 28314
rect 18804 28262 18816 28314
rect 18868 28262 18880 28314
rect 18932 28262 18944 28314
rect 18996 28262 19008 28314
rect 19060 28262 24686 28314
rect 24738 28262 24750 28314
rect 24802 28262 24814 28314
rect 24866 28262 24878 28314
rect 24930 28262 24942 28314
rect 24994 28262 25000 28314
rect 1104 28240 25000 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 1670 28200 1676 28212
rect 1627 28172 1676 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 1670 28160 1676 28172
rect 1728 28160 1734 28212
rect 2501 28203 2559 28209
rect 2501 28169 2513 28203
rect 2547 28200 2559 28203
rect 3970 28200 3976 28212
rect 2547 28172 3976 28200
rect 2547 28169 2559 28172
rect 2501 28163 2559 28169
rect 3970 28160 3976 28172
rect 4028 28160 4034 28212
rect 4065 28203 4123 28209
rect 4065 28169 4077 28203
rect 4111 28200 4123 28203
rect 5813 28203 5871 28209
rect 4111 28172 5764 28200
rect 4111 28169 4123 28172
rect 4065 28163 4123 28169
rect 2774 28132 2780 28144
rect 1688 28104 2780 28132
rect 1688 28076 1716 28104
rect 2774 28092 2780 28104
rect 2832 28092 2838 28144
rect 3145 28135 3203 28141
rect 3145 28101 3157 28135
rect 3191 28132 3203 28135
rect 3326 28132 3332 28144
rect 3191 28104 3332 28132
rect 3191 28101 3203 28104
rect 3145 28095 3203 28101
rect 3326 28092 3332 28104
rect 3384 28092 3390 28144
rect 3881 28135 3939 28141
rect 3881 28101 3893 28135
rect 3927 28132 3939 28135
rect 4154 28132 4160 28144
rect 3927 28104 4160 28132
rect 3927 28101 3939 28104
rect 3881 28095 3939 28101
rect 4154 28092 4160 28104
rect 4212 28092 4218 28144
rect 4246 28092 4252 28144
rect 4304 28132 4310 28144
rect 4522 28132 4528 28144
rect 4304 28104 4528 28132
rect 4304 28092 4310 28104
rect 4522 28092 4528 28104
rect 4580 28092 4586 28144
rect 5261 28135 5319 28141
rect 5261 28132 5273 28135
rect 4632 28104 5273 28132
rect 750 28024 756 28076
rect 808 28064 814 28076
rect 1489 28067 1547 28073
rect 1489 28064 1501 28067
rect 808 28036 1501 28064
rect 808 28024 814 28036
rect 1489 28033 1501 28036
rect 1535 28033 1547 28067
rect 1489 28027 1547 28033
rect 1670 28024 1676 28076
rect 1728 28024 1734 28076
rect 2314 28024 2320 28076
rect 2372 28024 2378 28076
rect 2958 28024 2964 28076
rect 3016 28064 3022 28076
rect 3053 28067 3111 28073
rect 3053 28064 3065 28067
rect 3016 28036 3065 28064
rect 3016 28024 3022 28036
rect 3053 28033 3065 28036
rect 3099 28033 3111 28067
rect 3053 28027 3111 28033
rect 3510 28024 3516 28076
rect 3568 28064 3574 28076
rect 4632 28064 4660 28104
rect 5261 28101 5273 28104
rect 5307 28101 5319 28135
rect 5261 28095 5319 28101
rect 5350 28092 5356 28144
rect 5408 28132 5414 28144
rect 5629 28135 5687 28141
rect 5629 28132 5641 28135
rect 5408 28104 5641 28132
rect 5408 28092 5414 28104
rect 5629 28101 5641 28104
rect 5675 28101 5687 28135
rect 5736 28132 5764 28172
rect 5813 28169 5825 28203
rect 5859 28200 5871 28203
rect 9950 28200 9956 28212
rect 5859 28172 9956 28200
rect 5859 28169 5871 28172
rect 5813 28163 5871 28169
rect 9950 28160 9956 28172
rect 10008 28160 10014 28212
rect 14918 28200 14924 28212
rect 10244 28172 14924 28200
rect 5736 28104 10088 28132
rect 5629 28095 5687 28101
rect 3568 28036 4660 28064
rect 3568 28024 3574 28036
rect 4798 28024 4804 28076
rect 4856 28024 4862 28076
rect 4893 28067 4951 28073
rect 4893 28033 4905 28067
rect 4939 28064 4951 28067
rect 5442 28064 5448 28076
rect 4939 28036 5448 28064
rect 4939 28033 4951 28036
rect 4893 28027 4951 28033
rect 5442 28024 5448 28036
rect 5500 28024 5506 28076
rect 5644 28008 5672 28095
rect 10060 28094 10088 28104
rect 6639 28067 6697 28073
rect 6639 28033 6651 28067
rect 6685 28064 6697 28067
rect 7650 28064 7656 28076
rect 6685 28036 7656 28064
rect 6685 28033 6697 28036
rect 6639 28027 6697 28033
rect 7650 28024 7656 28036
rect 7708 28024 7714 28076
rect 9582 28024 9588 28076
rect 9640 28064 9646 28076
rect 9784 28064 9994 28074
rect 10060 28066 10180 28094
rect 9640 28046 9994 28064
rect 9640 28036 9812 28046
rect 9640 28024 9646 28036
rect 3234 27956 3240 28008
rect 3292 27956 3298 28008
rect 4982 27956 4988 28008
rect 5040 27956 5046 28008
rect 5626 27956 5632 28008
rect 5684 27956 5690 28008
rect 6270 27956 6276 28008
rect 6328 27996 6334 28008
rect 6365 27999 6423 28005
rect 6365 27996 6377 27999
rect 6328 27968 6377 27996
rect 6328 27956 6334 27968
rect 6365 27965 6377 27968
rect 6411 27965 6423 27999
rect 6365 27959 6423 27965
rect 7190 27956 7196 28008
rect 7248 27996 7254 28008
rect 9858 27996 9864 28008
rect 7248 27968 9864 27996
rect 7248 27956 7254 27968
rect 9858 27956 9864 27968
rect 9916 27956 9922 28008
rect 9966 27996 9994 28046
rect 10152 28064 10180 28066
rect 10244 28064 10272 28172
rect 14918 28160 14924 28172
rect 14976 28160 14982 28212
rect 16209 28203 16267 28209
rect 16209 28169 16221 28203
rect 16255 28200 16267 28203
rect 16666 28200 16672 28212
rect 16255 28172 16672 28200
rect 16255 28169 16267 28172
rect 16209 28163 16267 28169
rect 16666 28160 16672 28172
rect 16724 28160 16730 28212
rect 16776 28172 19472 28200
rect 11146 28092 11152 28144
rect 11204 28132 11210 28144
rect 11698 28132 11704 28144
rect 11204 28104 11704 28132
rect 11204 28092 11210 28104
rect 11698 28092 11704 28104
rect 11756 28092 11762 28144
rect 14734 28092 14740 28144
rect 14792 28132 14798 28144
rect 16776 28132 16804 28172
rect 19444 28144 19472 28172
rect 19610 28160 19616 28212
rect 19668 28200 19674 28212
rect 19668 28172 19748 28200
rect 19668 28160 19674 28172
rect 14792 28104 16804 28132
rect 14792 28092 14798 28104
rect 17310 28092 17316 28144
rect 17368 28132 17374 28144
rect 17770 28132 17776 28144
rect 17368 28104 17776 28132
rect 17368 28092 17374 28104
rect 17770 28092 17776 28104
rect 17828 28092 17834 28144
rect 19334 28132 19340 28144
rect 17880 28104 19340 28132
rect 10152 28036 10272 28064
rect 10319 28077 10377 28083
rect 10319 28043 10331 28077
rect 10365 28074 10377 28077
rect 10410 28074 10416 28076
rect 10365 28046 10416 28074
rect 10365 28043 10377 28046
rect 10319 28037 10377 28043
rect 10410 28024 10416 28046
rect 10468 28024 10474 28076
rect 11054 28024 11060 28076
rect 11112 28064 11118 28076
rect 11330 28064 11336 28076
rect 11112 28036 11336 28064
rect 11112 28024 11118 28036
rect 11330 28024 11336 28036
rect 11388 28024 11394 28076
rect 13170 28064 13176 28076
rect 12406 28036 13176 28064
rect 10045 27999 10103 28005
rect 10045 27996 10057 27999
rect 9966 27968 10057 27996
rect 10045 27965 10057 27968
rect 10091 27965 10103 27999
rect 12406 27996 12434 28036
rect 13170 28024 13176 28036
rect 13228 28024 13234 28076
rect 13998 28024 14004 28076
rect 14056 28024 14062 28076
rect 15439 28067 15497 28073
rect 15439 28064 15451 28067
rect 14936 28036 15451 28064
rect 10045 27959 10103 27965
rect 10704 27968 12434 27996
rect 7282 27888 7288 27940
rect 7340 27928 7346 27940
rect 7340 27900 9674 27928
rect 7340 27888 7346 27900
rect 6822 27820 6828 27872
rect 6880 27860 6886 27872
rect 7377 27863 7435 27869
rect 7377 27860 7389 27863
rect 6880 27832 7389 27860
rect 6880 27820 6886 27832
rect 7377 27829 7389 27832
rect 7423 27829 7435 27863
rect 9646 27860 9674 27900
rect 10704 27860 10732 27968
rect 12618 27956 12624 28008
rect 12676 27996 12682 28008
rect 12805 27999 12863 28005
rect 12805 27996 12817 27999
rect 12676 27968 12817 27996
rect 12676 27956 12682 27968
rect 12805 27965 12817 27968
rect 12851 27965 12863 27999
rect 12805 27959 12863 27965
rect 12986 27956 12992 28008
rect 13044 27956 13050 28008
rect 13725 27999 13783 28005
rect 13725 27996 13737 27999
rect 13096 27968 13737 27996
rect 11698 27888 11704 27940
rect 11756 27928 11762 27940
rect 13096 27928 13124 27968
rect 13725 27965 13737 27968
rect 13771 27965 13783 27999
rect 13725 27959 13783 27965
rect 13814 27956 13820 28008
rect 13872 28005 13878 28008
rect 13872 27999 13900 28005
rect 13888 27965 13900 27999
rect 13872 27959 13900 27965
rect 13872 27956 13878 27959
rect 14366 27956 14372 28008
rect 14424 27996 14430 28008
rect 14642 27996 14648 28008
rect 14424 27968 14648 27996
rect 14424 27956 14430 27968
rect 14642 27956 14648 27968
rect 14700 27956 14706 28008
rect 11756 27900 13124 27928
rect 13449 27931 13507 27937
rect 11756 27888 11762 27900
rect 13449 27897 13461 27931
rect 13495 27897 13507 27931
rect 14936 27928 14964 28036
rect 15439 28033 15451 28036
rect 15485 28033 15497 28067
rect 15439 28027 15497 28033
rect 17678 28024 17684 28076
rect 17736 28064 17742 28076
rect 17880 28073 17908 28104
rect 19334 28092 19340 28104
rect 19392 28092 19398 28144
rect 19426 28092 19432 28144
rect 19484 28092 19490 28144
rect 19720 28141 19748 28172
rect 20990 28160 20996 28212
rect 21048 28160 21054 28212
rect 21082 28160 21088 28212
rect 21140 28200 21146 28212
rect 23477 28203 23535 28209
rect 21140 28172 22048 28200
rect 21140 28160 21146 28172
rect 19696 28135 19754 28141
rect 19696 28101 19708 28135
rect 19742 28101 19754 28135
rect 19696 28095 19754 28101
rect 21008 28132 21036 28160
rect 21008 28104 21864 28132
rect 17865 28067 17923 28073
rect 17865 28064 17877 28067
rect 17736 28036 17877 28064
rect 17736 28024 17742 28036
rect 17865 28033 17877 28036
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 17954 28024 17960 28076
rect 18012 28064 18018 28076
rect 18121 28067 18179 28073
rect 18121 28064 18133 28067
rect 18012 28036 18133 28064
rect 18012 28024 18018 28036
rect 18121 28033 18133 28036
rect 18167 28033 18179 28067
rect 18121 28027 18179 28033
rect 18598 28024 18604 28076
rect 18656 28064 18662 28076
rect 20901 28067 20959 28073
rect 18656 28036 19288 28064
rect 18656 28024 18662 28036
rect 15194 27956 15200 28008
rect 15252 27956 15258 28008
rect 19260 27937 19288 28036
rect 20901 28033 20913 28067
rect 20947 28064 20959 28067
rect 21008 28064 21036 28104
rect 21836 28073 21864 28104
rect 22020 28073 22048 28172
rect 23477 28169 23489 28203
rect 23523 28169 23535 28203
rect 23477 28163 23535 28169
rect 22186 28092 22192 28144
rect 22244 28132 22250 28144
rect 22922 28132 22928 28144
rect 22244 28104 22928 28132
rect 22244 28092 22250 28104
rect 22922 28092 22928 28104
rect 22980 28132 22986 28144
rect 23492 28132 23520 28163
rect 22980 28104 23152 28132
rect 22980 28092 22986 28104
rect 21269 28067 21327 28073
rect 21269 28064 21281 28067
rect 20947 28036 21036 28064
rect 21100 28036 21281 28064
rect 20947 28033 20959 28036
rect 20901 28027 20959 28033
rect 19426 27956 19432 28008
rect 19484 27956 19490 28008
rect 20714 27956 20720 28008
rect 20772 27996 20778 28008
rect 21100 27996 21128 28036
rect 21269 28033 21281 28036
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 21821 28067 21879 28073
rect 21821 28033 21833 28067
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22281 28067 22339 28073
rect 22281 28064 22293 28067
rect 22152 28036 22293 28064
rect 22152 28024 22158 28036
rect 22281 28033 22293 28036
rect 22327 28033 22339 28067
rect 22281 28027 22339 28033
rect 22830 28024 22836 28076
rect 22888 28024 22894 28076
rect 23124 28073 23152 28104
rect 23490 28104 23520 28132
rect 23109 28067 23167 28073
rect 23109 28033 23121 28067
rect 23155 28033 23167 28067
rect 23109 28027 23167 28033
rect 23385 28067 23443 28073
rect 23385 28033 23397 28067
rect 23431 28062 23443 28067
rect 23490 28062 23518 28104
rect 23431 28034 23518 28062
rect 23661 28067 23719 28073
rect 23431 28033 23443 28034
rect 23385 28027 23443 28033
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 20772 27968 21128 27996
rect 21177 27999 21235 28005
rect 20772 27956 20778 27968
rect 21177 27965 21189 27999
rect 21223 27996 21235 27999
rect 21913 27999 21971 28005
rect 21913 27996 21925 27999
rect 21223 27968 21925 27996
rect 21223 27965 21235 27968
rect 21177 27959 21235 27965
rect 21913 27965 21925 27968
rect 21959 27965 21971 27999
rect 23676 27996 23704 28027
rect 23934 28024 23940 28076
rect 23992 28024 23998 28076
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28033 24179 28067
rect 24121 28027 24179 28033
rect 21913 27959 21971 27965
rect 22940 27968 23704 27996
rect 13449 27891 13507 27897
rect 14384 27900 14964 27928
rect 19245 27931 19303 27937
rect 9646 27832 10732 27860
rect 7377 27823 7435 27829
rect 11054 27820 11060 27872
rect 11112 27820 11118 27872
rect 11422 27820 11428 27872
rect 11480 27860 11486 27872
rect 11974 27860 11980 27872
rect 11480 27832 11980 27860
rect 11480 27820 11486 27832
rect 11974 27820 11980 27832
rect 12032 27860 12038 27872
rect 12986 27860 12992 27872
rect 12032 27832 12992 27860
rect 12032 27820 12038 27832
rect 12986 27820 12992 27832
rect 13044 27820 13050 27872
rect 13464 27860 13492 27891
rect 13722 27860 13728 27872
rect 13464 27832 13728 27860
rect 13722 27820 13728 27832
rect 13780 27820 13786 27872
rect 13906 27820 13912 27872
rect 13964 27860 13970 27872
rect 14384 27860 14412 27900
rect 14752 27872 14780 27900
rect 19245 27897 19257 27931
rect 19291 27897 19303 27931
rect 19245 27891 19303 27897
rect 20993 27931 21051 27937
rect 20993 27897 21005 27931
rect 21039 27928 21051 27931
rect 21361 27931 21419 27937
rect 21361 27928 21373 27931
rect 21039 27900 21373 27928
rect 21039 27897 21051 27900
rect 20993 27891 21051 27897
rect 21361 27897 21373 27900
rect 21407 27897 21419 27931
rect 22554 27928 22560 27940
rect 21361 27891 21419 27897
rect 22020 27900 22560 27928
rect 13964 27832 14412 27860
rect 13964 27820 13970 27832
rect 14642 27820 14648 27872
rect 14700 27820 14706 27872
rect 14734 27820 14740 27872
rect 14792 27820 14798 27872
rect 14918 27820 14924 27872
rect 14976 27860 14982 27872
rect 19610 27860 19616 27872
rect 14976 27832 19616 27860
rect 14976 27820 14982 27832
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 20806 27820 20812 27872
rect 20864 27820 20870 27872
rect 21085 27863 21143 27869
rect 21085 27829 21097 27863
rect 21131 27860 21143 27863
rect 22020 27860 22048 27900
rect 22554 27888 22560 27900
rect 22612 27888 22618 27940
rect 22940 27937 22968 27968
rect 22925 27931 22983 27937
rect 22925 27897 22937 27931
rect 22971 27897 22983 27931
rect 22925 27891 22983 27897
rect 23201 27931 23259 27937
rect 23201 27897 23213 27931
rect 23247 27928 23259 27931
rect 24136 27928 24164 28027
rect 23247 27900 24164 27928
rect 23247 27897 23259 27900
rect 23201 27891 23259 27897
rect 21131 27832 22048 27860
rect 22097 27863 22155 27869
rect 21131 27829 21143 27832
rect 21085 27823 21143 27829
rect 22097 27829 22109 27863
rect 22143 27860 22155 27863
rect 22462 27860 22468 27872
rect 22143 27832 22468 27860
rect 22143 27829 22155 27832
rect 22097 27823 22155 27829
rect 22462 27820 22468 27832
rect 22520 27820 22526 27872
rect 22649 27863 22707 27869
rect 22649 27829 22661 27863
rect 22695 27860 22707 27863
rect 23014 27860 23020 27872
rect 22695 27832 23020 27860
rect 22695 27829 22707 27832
rect 22649 27823 22707 27829
rect 23014 27820 23020 27832
rect 23072 27820 23078 27872
rect 23750 27820 23756 27872
rect 23808 27820 23814 27872
rect 24394 27820 24400 27872
rect 24452 27820 24458 27872
rect 1104 27770 24840 27792
rect 1104 27718 3917 27770
rect 3969 27718 3981 27770
rect 4033 27718 4045 27770
rect 4097 27718 4109 27770
rect 4161 27718 4173 27770
rect 4225 27718 9851 27770
rect 9903 27718 9915 27770
rect 9967 27718 9979 27770
rect 10031 27718 10043 27770
rect 10095 27718 10107 27770
rect 10159 27718 15785 27770
rect 15837 27718 15849 27770
rect 15901 27718 15913 27770
rect 15965 27718 15977 27770
rect 16029 27718 16041 27770
rect 16093 27718 21719 27770
rect 21771 27718 21783 27770
rect 21835 27718 21847 27770
rect 21899 27718 21911 27770
rect 21963 27718 21975 27770
rect 22027 27718 24840 27770
rect 1104 27696 24840 27718
rect 474 27616 480 27668
rect 532 27656 538 27668
rect 3326 27656 3332 27668
rect 532 27628 3332 27656
rect 532 27616 538 27628
rect 3326 27616 3332 27628
rect 3384 27616 3390 27668
rect 4522 27616 4528 27668
rect 4580 27656 4586 27668
rect 6362 27656 6368 27668
rect 4580 27628 6368 27656
rect 4580 27616 4586 27628
rect 6362 27616 6368 27628
rect 6420 27616 6426 27668
rect 10318 27616 10324 27668
rect 10376 27656 10382 27668
rect 10376 27628 19380 27656
rect 10376 27616 10382 27628
rect 5813 27591 5871 27597
rect 5813 27557 5825 27591
rect 5859 27557 5871 27591
rect 5813 27551 5871 27557
rect 1394 27480 1400 27532
rect 1452 27480 1458 27532
rect 5828 27520 5856 27551
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 8018 27588 8024 27600
rect 7892 27560 8024 27588
rect 7892 27548 7898 27560
rect 8018 27548 8024 27560
rect 8076 27548 8082 27600
rect 10410 27548 10416 27600
rect 10468 27548 10474 27600
rect 15286 27588 15292 27600
rect 12176 27560 15292 27588
rect 5828 27492 6210 27520
rect 8754 27480 8760 27532
rect 8812 27520 8818 27532
rect 8812 27492 8970 27520
rect 8812 27480 8818 27492
rect 1578 27412 1584 27464
rect 1636 27452 1642 27464
rect 1671 27455 1729 27461
rect 1671 27452 1683 27455
rect 1636 27424 1683 27452
rect 1636 27412 1642 27424
rect 1671 27421 1683 27424
rect 1717 27421 1729 27455
rect 1671 27415 1729 27421
rect 2777 27455 2835 27461
rect 2777 27421 2789 27455
rect 2823 27421 2835 27455
rect 2777 27415 2835 27421
rect 1210 27344 1216 27396
rect 1268 27384 1274 27396
rect 2792 27384 2820 27415
rect 4430 27412 4436 27464
rect 4488 27452 4494 27464
rect 4801 27455 4859 27461
rect 4801 27452 4813 27455
rect 4488 27424 4813 27452
rect 4488 27412 4494 27424
rect 4801 27421 4813 27424
rect 4847 27452 4859 27455
rect 4982 27452 4988 27464
rect 4847 27424 4988 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5075 27455 5133 27461
rect 5075 27421 5087 27455
rect 5121 27452 5133 27455
rect 6546 27452 6552 27464
rect 5121 27424 6552 27452
rect 5121 27421 5133 27424
rect 5075 27415 5133 27421
rect 6546 27412 6552 27424
rect 6604 27412 6610 27464
rect 6822 27412 6828 27464
rect 6880 27412 6886 27464
rect 7098 27412 7104 27464
rect 7156 27452 7162 27464
rect 7834 27452 7840 27464
rect 7156 27424 7840 27452
rect 7156 27412 7162 27424
rect 7834 27412 7840 27424
rect 7892 27412 7898 27464
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27452 9551 27455
rect 9674 27452 9680 27464
rect 9539 27424 9680 27452
rect 9539 27421 9551 27424
rect 9493 27415 9551 27421
rect 9674 27412 9680 27424
rect 9732 27412 9738 27464
rect 11422 27452 11428 27464
rect 9784 27424 11428 27452
rect 1268 27356 2820 27384
rect 6641 27387 6699 27393
rect 1268 27344 1274 27356
rect 6641 27353 6653 27387
rect 6687 27353 6699 27387
rect 6641 27347 6699 27353
rect 6733 27387 6791 27393
rect 6733 27353 6745 27387
rect 6779 27384 6791 27387
rect 6838 27384 6866 27412
rect 6779 27356 6866 27384
rect 7392 27356 9352 27384
rect 6779 27353 6791 27356
rect 6733 27347 6791 27353
rect 2038 27276 2044 27328
rect 2096 27316 2102 27328
rect 2409 27319 2467 27325
rect 2409 27316 2421 27319
rect 2096 27288 2421 27316
rect 2096 27276 2102 27288
rect 2409 27285 2421 27288
rect 2455 27285 2467 27319
rect 2409 27279 2467 27285
rect 2958 27276 2964 27328
rect 3016 27276 3022 27328
rect 4982 27276 4988 27328
rect 5040 27316 5046 27328
rect 6270 27316 6276 27328
rect 5040 27288 6276 27316
rect 5040 27276 5046 27288
rect 6270 27276 6276 27288
rect 6328 27276 6334 27328
rect 6362 27276 6368 27328
rect 6420 27276 6426 27328
rect 6454 27276 6460 27328
rect 6512 27316 6518 27328
rect 6654 27316 6682 27347
rect 6512 27288 6682 27316
rect 6512 27276 6518 27288
rect 6822 27276 6828 27328
rect 6880 27316 6886 27328
rect 7392 27316 7420 27356
rect 6880 27288 7420 27316
rect 6880 27276 6886 27288
rect 7466 27276 7472 27328
rect 7524 27276 7530 27328
rect 7650 27276 7656 27328
rect 7708 27276 7714 27328
rect 9125 27319 9183 27325
rect 9125 27285 9137 27319
rect 9171 27316 9183 27319
rect 9214 27316 9220 27328
rect 9171 27288 9220 27316
rect 9171 27285 9183 27288
rect 9125 27279 9183 27285
rect 9214 27276 9220 27288
rect 9272 27276 9278 27328
rect 9324 27316 9352 27356
rect 9398 27344 9404 27396
rect 9456 27344 9462 27396
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 9784 27384 9812 27424
rect 9640 27356 9812 27384
rect 9640 27344 9646 27356
rect 9858 27344 9864 27396
rect 9916 27344 9922 27396
rect 10244 27393 10272 27424
rect 11422 27412 11428 27424
rect 11480 27412 11486 27464
rect 11514 27412 11520 27464
rect 11572 27412 11578 27464
rect 11775 27425 11833 27431
rect 10229 27387 10287 27393
rect 10229 27353 10241 27387
rect 10275 27353 10287 27387
rect 11775 27391 11787 27425
rect 11821 27422 11833 27425
rect 11821 27396 11834 27422
rect 11775 27385 11796 27391
rect 10229 27347 10287 27353
rect 11790 27344 11796 27385
rect 11848 27384 11854 27396
rect 12066 27384 12072 27396
rect 11848 27356 12072 27384
rect 11848 27344 11854 27356
rect 12066 27344 12072 27356
rect 12124 27344 12130 27396
rect 12176 27316 12204 27560
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 12342 27480 12348 27532
rect 12400 27480 12406 27532
rect 12526 27480 12532 27532
rect 12584 27520 12590 27532
rect 15838 27520 15844 27532
rect 12584 27492 15844 27520
rect 12584 27480 12590 27492
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 19352 27520 19380 27628
rect 22462 27616 22468 27668
rect 22520 27616 22526 27668
rect 22557 27659 22615 27665
rect 22557 27625 22569 27659
rect 22603 27656 22615 27659
rect 22830 27656 22836 27668
rect 22603 27628 22836 27656
rect 22603 27625 22615 27628
rect 22557 27619 22615 27625
rect 22830 27616 22836 27628
rect 22888 27616 22894 27668
rect 23014 27616 23020 27668
rect 23072 27656 23078 27668
rect 23569 27659 23627 27665
rect 23072 27628 23428 27656
rect 23072 27616 23078 27628
rect 19981 27591 20039 27597
rect 19981 27557 19993 27591
rect 20027 27588 20039 27591
rect 20714 27588 20720 27600
rect 20027 27560 20720 27588
rect 20027 27557 20039 27560
rect 19981 27551 20039 27557
rect 20714 27548 20720 27560
rect 20772 27548 20778 27600
rect 20806 27548 20812 27600
rect 20864 27548 20870 27600
rect 20901 27591 20959 27597
rect 20901 27557 20913 27591
rect 20947 27588 20959 27591
rect 21082 27588 21088 27600
rect 20947 27560 21088 27588
rect 20947 27557 20959 27560
rect 20901 27551 20959 27557
rect 21082 27548 21088 27560
rect 21140 27548 21146 27600
rect 19352 27492 20760 27520
rect 12360 27452 12388 27480
rect 13998 27452 14004 27464
rect 12360 27424 14004 27452
rect 13998 27412 14004 27424
rect 14056 27412 14062 27464
rect 14642 27412 14648 27464
rect 14700 27452 14706 27464
rect 15197 27455 15255 27461
rect 15197 27452 15209 27455
rect 14700 27424 15209 27452
rect 14700 27412 14706 27424
rect 15197 27421 15209 27424
rect 15243 27421 15255 27455
rect 15197 27415 15255 27421
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 15562 27452 15568 27464
rect 15344 27424 15568 27452
rect 15344 27412 15350 27424
rect 15562 27412 15568 27424
rect 15620 27412 15626 27464
rect 16482 27461 16488 27464
rect 16209 27455 16267 27461
rect 16209 27421 16221 27455
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 16467 27455 16488 27461
rect 16467 27421 16479 27455
rect 16467 27415 16488 27421
rect 13814 27384 13820 27396
rect 12452 27356 13820 27384
rect 9324 27288 12204 27316
rect 12250 27276 12256 27328
rect 12308 27316 12314 27328
rect 12452 27316 12480 27356
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 16224 27384 16252 27415
rect 16482 27412 16488 27415
rect 16540 27412 16546 27464
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 16592 27424 17601 27452
rect 15212 27356 16252 27384
rect 15212 27328 15240 27356
rect 12308 27288 12480 27316
rect 12529 27319 12587 27325
rect 12308 27276 12314 27288
rect 12529 27285 12541 27319
rect 12575 27316 12587 27319
rect 12710 27316 12716 27328
rect 12575 27288 12716 27316
rect 12575 27285 12587 27288
rect 12529 27279 12587 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 13630 27276 13636 27328
rect 13688 27316 13694 27328
rect 14918 27316 14924 27328
rect 13688 27288 14924 27316
rect 13688 27276 13694 27288
rect 14918 27276 14924 27288
rect 14976 27276 14982 27328
rect 15010 27276 15016 27328
rect 15068 27276 15074 27328
rect 15194 27276 15200 27328
rect 15252 27276 15258 27328
rect 16224 27316 16252 27356
rect 16592 27328 16620 27424
rect 17589 27421 17601 27424
rect 17635 27421 17647 27455
rect 17831 27455 17889 27461
rect 17831 27452 17843 27455
rect 17589 27415 17647 27421
rect 17696 27424 17843 27452
rect 17696 27384 17724 27424
rect 17831 27421 17843 27424
rect 17877 27421 17889 27455
rect 17831 27415 17889 27421
rect 19610 27412 19616 27464
rect 19668 27452 19674 27464
rect 20165 27455 20223 27461
rect 20165 27452 20177 27455
rect 19668 27424 20177 27452
rect 19668 27412 19674 27424
rect 20165 27421 20177 27424
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 17420 27356 17724 27384
rect 20732 27384 20760 27492
rect 20824 27452 20852 27548
rect 22480 27520 22508 27616
rect 22741 27591 22799 27597
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 23109 27591 23167 27597
rect 23109 27588 23121 27591
rect 22787 27560 23121 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 23109 27557 23121 27560
rect 23155 27557 23167 27591
rect 23400 27588 23428 27628
rect 23569 27625 23581 27659
rect 23615 27656 23627 27659
rect 23934 27656 23940 27668
rect 23615 27628 23940 27656
rect 23615 27625 23627 27628
rect 23569 27619 23627 27625
rect 23934 27616 23940 27628
rect 23992 27616 23998 27668
rect 23400 27560 23520 27588
rect 23109 27551 23167 27557
rect 22925 27523 22983 27529
rect 22480 27492 22784 27520
rect 21085 27455 21143 27461
rect 21085 27452 21097 27455
rect 20824 27424 21097 27452
rect 21085 27421 21097 27424
rect 21131 27421 21143 27455
rect 21085 27415 21143 27421
rect 21174 27412 21180 27464
rect 21232 27412 21238 27464
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27421 22707 27455
rect 22756 27452 22784 27492
rect 22925 27489 22937 27523
rect 22971 27520 22983 27523
rect 23385 27523 23443 27529
rect 23385 27520 23397 27523
rect 22971 27492 23397 27520
rect 22971 27489 22983 27492
rect 22925 27483 22983 27489
rect 23385 27489 23397 27492
rect 23431 27489 23443 27523
rect 23385 27483 23443 27489
rect 23492 27461 23520 27560
rect 23566 27480 23572 27532
rect 23624 27520 23630 27532
rect 23624 27492 23980 27520
rect 23624 27480 23630 27492
rect 23952 27461 23980 27492
rect 23017 27455 23075 27461
rect 23017 27452 23029 27455
rect 22756 27424 23029 27452
rect 22649 27415 22707 27421
rect 23017 27421 23029 27424
rect 23063 27421 23075 27455
rect 23017 27415 23075 27421
rect 23293 27455 23351 27461
rect 23293 27421 23305 27455
rect 23339 27421 23351 27455
rect 23293 27415 23351 27421
rect 23477 27455 23535 27461
rect 23477 27421 23489 27455
rect 23523 27421 23535 27455
rect 23477 27415 23535 27421
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27421 23811 27455
rect 23753 27415 23811 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 21422 27387 21480 27393
rect 21422 27384 21434 27387
rect 20732 27356 21434 27384
rect 17420 27328 17448 27356
rect 21422 27353 21434 27356
rect 21468 27384 21480 27387
rect 22002 27384 22008 27396
rect 21468 27356 22008 27384
rect 21468 27353 21480 27356
rect 21422 27347 21480 27353
rect 22002 27344 22008 27356
rect 22060 27344 22066 27396
rect 22664 27384 22692 27415
rect 22830 27384 22836 27396
rect 22664 27356 22836 27384
rect 22830 27344 22836 27356
rect 22888 27384 22894 27396
rect 23308 27384 23336 27415
rect 22888 27356 23336 27384
rect 22888 27344 22894 27356
rect 16574 27316 16580 27328
rect 16224 27288 16580 27316
rect 16574 27276 16580 27288
rect 16632 27276 16638 27328
rect 17218 27276 17224 27328
rect 17276 27276 17282 27328
rect 17402 27276 17408 27328
rect 17460 27276 17466 27328
rect 17862 27276 17868 27328
rect 17920 27316 17926 27328
rect 18601 27319 18659 27325
rect 18601 27316 18613 27319
rect 17920 27288 18613 27316
rect 17920 27276 17926 27288
rect 18601 27285 18613 27288
rect 18647 27285 18659 27319
rect 18601 27279 18659 27285
rect 19334 27276 19340 27328
rect 19392 27316 19398 27328
rect 21174 27316 21180 27328
rect 19392 27288 21180 27316
rect 19392 27276 19398 27288
rect 21174 27276 21180 27288
rect 21232 27276 21238 27328
rect 22922 27276 22928 27328
rect 22980 27276 22986 27328
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23768 27316 23796 27415
rect 23072 27288 23796 27316
rect 24121 27319 24179 27325
rect 23072 27276 23078 27288
rect 24121 27285 24133 27319
rect 24167 27316 24179 27319
rect 25130 27316 25136 27328
rect 24167 27288 25136 27316
rect 24167 27285 24179 27288
rect 24121 27279 24179 27285
rect 25130 27276 25136 27288
rect 25188 27276 25194 27328
rect 1104 27226 25000 27248
rect 1104 27174 6884 27226
rect 6936 27174 6948 27226
rect 7000 27174 7012 27226
rect 7064 27174 7076 27226
rect 7128 27174 7140 27226
rect 7192 27174 12818 27226
rect 12870 27174 12882 27226
rect 12934 27174 12946 27226
rect 12998 27174 13010 27226
rect 13062 27174 13074 27226
rect 13126 27174 18752 27226
rect 18804 27174 18816 27226
rect 18868 27174 18880 27226
rect 18932 27174 18944 27226
rect 18996 27174 19008 27226
rect 19060 27174 24686 27226
rect 24738 27174 24750 27226
rect 24802 27174 24814 27226
rect 24866 27174 24878 27226
rect 24930 27174 24942 27226
rect 24994 27174 25000 27226
rect 1104 27152 25000 27174
rect 1670 27072 1676 27124
rect 1728 27112 1734 27124
rect 2041 27115 2099 27121
rect 2041 27112 2053 27115
rect 1728 27084 2053 27112
rect 1728 27072 1734 27084
rect 2041 27081 2053 27084
rect 2087 27081 2099 27115
rect 2774 27112 2780 27124
rect 2041 27075 2099 27081
rect 2240 27084 2780 27112
rect 2240 26976 2268 27084
rect 2774 27072 2780 27084
rect 2832 27072 2838 27124
rect 2958 27072 2964 27124
rect 3016 27112 3022 27124
rect 3145 27115 3203 27121
rect 3145 27112 3157 27115
rect 3016 27084 3157 27112
rect 3016 27072 3022 27084
rect 3145 27081 3157 27084
rect 3191 27081 3203 27115
rect 3145 27075 3203 27081
rect 3326 27072 3332 27124
rect 3384 27072 3390 27124
rect 3697 27115 3755 27121
rect 3697 27081 3709 27115
rect 3743 27112 3755 27115
rect 3743 27084 5396 27112
rect 3743 27081 3755 27084
rect 3697 27075 3755 27081
rect 2590 27004 2596 27056
rect 2648 27044 2654 27056
rect 2648 27016 3556 27044
rect 2648 27004 2654 27016
rect 2317 26979 2375 26985
rect 2317 26976 2329 26979
rect 2240 26948 2329 26976
rect 2317 26945 2329 26948
rect 2363 26945 2375 26979
rect 2317 26939 2375 26945
rect 2406 26936 2412 26988
rect 2464 26936 2470 26988
rect 3528 26985 3556 27016
rect 4522 27004 4528 27056
rect 4580 27044 4586 27056
rect 4982 27044 4988 27056
rect 4580 27016 4752 27044
rect 4580 27004 4586 27016
rect 4724 27006 4752 27016
rect 4908 27016 4988 27044
rect 4783 27009 4841 27015
rect 4783 27006 4795 27009
rect 2777 26979 2835 26985
rect 2777 26945 2789 26979
rect 2823 26976 2835 26979
rect 3513 26979 3571 26985
rect 2823 26948 3464 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 2044 26920 2096 26926
rect 3436 26908 3464 26948
rect 3513 26945 3525 26979
rect 3559 26945 3571 26979
rect 3513 26939 3571 26945
rect 3786 26936 3792 26988
rect 3844 26936 3850 26988
rect 4724 26978 4795 27006
rect 4783 26975 4795 26978
rect 4829 27006 4841 27009
rect 4908 27006 4936 27016
rect 4829 26978 4936 27006
rect 4982 27004 4988 27016
rect 5040 27004 5046 27056
rect 5368 27044 5396 27084
rect 5442 27072 5448 27124
rect 5500 27112 5506 27124
rect 5537 27115 5595 27121
rect 5537 27112 5549 27115
rect 5500 27084 5549 27112
rect 5500 27072 5506 27084
rect 5537 27081 5549 27084
rect 5583 27081 5595 27115
rect 5537 27075 5595 27081
rect 8110 27072 8116 27124
rect 8168 27112 8174 27124
rect 8478 27112 8484 27124
rect 8168 27084 8484 27112
rect 8168 27072 8174 27084
rect 8478 27072 8484 27084
rect 8536 27072 8542 27124
rect 8754 27072 8760 27124
rect 8812 27072 8818 27124
rect 9398 27072 9404 27124
rect 9456 27112 9462 27124
rect 10502 27112 10508 27124
rect 9456 27084 10508 27112
rect 9456 27072 9462 27084
rect 10502 27072 10508 27084
rect 10560 27072 10566 27124
rect 11606 27072 11612 27124
rect 11664 27112 11670 27124
rect 12526 27112 12532 27124
rect 11664 27084 12532 27112
rect 11664 27072 11670 27084
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 13630 27112 13636 27124
rect 12820 27084 13636 27112
rect 12618 27044 12624 27056
rect 5368 27016 12624 27044
rect 12618 27004 12624 27016
rect 12676 27044 12682 27056
rect 12820 27044 12848 27084
rect 13630 27072 13636 27084
rect 13688 27072 13694 27124
rect 13998 27072 14004 27124
rect 14056 27112 14062 27124
rect 14645 27115 14703 27121
rect 14056 27084 14596 27112
rect 14056 27072 14062 27084
rect 12676 27016 12848 27044
rect 12676 27004 12682 27016
rect 8019 26979 8077 26985
rect 4829 26975 4841 26978
rect 4783 26969 4841 26975
rect 8019 26945 8031 26979
rect 8065 26976 8077 26979
rect 8110 26976 8116 26988
rect 8065 26948 8116 26976
rect 8065 26945 8077 26948
rect 8019 26939 8077 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 12820 26985 12848 27016
rect 14568 27044 14596 27084
rect 14645 27081 14657 27115
rect 14691 27112 14703 27115
rect 19334 27112 19340 27124
rect 14691 27084 19340 27112
rect 14691 27081 14703 27084
rect 14645 27075 14703 27081
rect 19334 27072 19340 27084
rect 19392 27072 19398 27124
rect 19812 27084 22094 27112
rect 19812 27056 19840 27084
rect 15194 27044 15200 27056
rect 14568 27016 15200 27044
rect 12805 26979 12863 26985
rect 12805 26945 12817 26979
rect 12851 26945 12863 26979
rect 12805 26939 12863 26945
rect 13814 26936 13820 26988
rect 13872 26985 13878 26988
rect 13872 26979 13900 26985
rect 13888 26945 13900 26979
rect 14568 26976 14596 27016
rect 15194 27004 15200 27016
rect 15252 27004 15258 27056
rect 15838 27004 15844 27056
rect 15896 27004 15902 27056
rect 19794 27004 19800 27056
rect 19852 27004 19858 27056
rect 21082 27004 21088 27056
rect 21140 27044 21146 27056
rect 21634 27044 21640 27056
rect 21140 27016 21640 27044
rect 21140 27004 21146 27016
rect 21634 27004 21640 27016
rect 21692 27004 21698 27056
rect 22066 27044 22094 27084
rect 22830 27072 22836 27124
rect 22888 27072 22894 27124
rect 23014 27072 23020 27124
rect 23072 27072 23078 27124
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27112 23351 27115
rect 23566 27112 23572 27124
rect 23339 27084 23572 27112
rect 23339 27081 23351 27084
rect 23293 27075 23351 27081
rect 23566 27072 23572 27084
rect 23624 27072 23630 27124
rect 23750 27072 23756 27124
rect 23808 27072 23814 27124
rect 23937 27115 23995 27121
rect 23937 27081 23949 27115
rect 23983 27081 23995 27115
rect 23937 27075 23995 27081
rect 23032 27044 23060 27072
rect 23768 27044 23796 27072
rect 22066 27016 23060 27044
rect 23492 27016 23796 27044
rect 23952 27044 23980 27075
rect 23952 27016 24256 27044
rect 14737 26979 14795 26985
rect 14737 26976 14749 26979
rect 14568 26948 14749 26976
rect 13872 26939 13900 26945
rect 14737 26945 14749 26948
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 13872 26936 13878 26939
rect 14918 26936 14924 26988
rect 14976 26976 14982 26988
rect 15011 26979 15069 26985
rect 15011 26976 15023 26979
rect 14976 26948 15023 26976
rect 14976 26936 14982 26948
rect 15011 26945 15023 26948
rect 15057 26945 15069 26979
rect 15011 26939 15069 26945
rect 3602 26908 3608 26920
rect 3436 26880 3608 26908
rect 3602 26868 3608 26880
rect 3660 26868 3666 26920
rect 3804 26908 3832 26936
rect 4522 26908 4528 26920
rect 3804 26880 4528 26908
rect 4522 26868 4528 26880
rect 4580 26868 4586 26920
rect 7742 26868 7748 26920
rect 7800 26868 7806 26920
rect 9214 26868 9220 26920
rect 9272 26908 9278 26920
rect 9766 26908 9772 26920
rect 9272 26880 9772 26908
rect 9272 26868 9278 26880
rect 9766 26868 9772 26880
rect 9824 26868 9830 26920
rect 9858 26868 9864 26920
rect 9916 26908 9922 26920
rect 12250 26908 12256 26920
rect 9916 26880 12256 26908
rect 9916 26868 9922 26880
rect 12250 26868 12256 26880
rect 12308 26868 12314 26920
rect 12989 26911 13047 26917
rect 12989 26877 13001 26911
rect 13035 26908 13047 26911
rect 13354 26908 13360 26920
rect 13035 26880 13360 26908
rect 13035 26877 13047 26880
rect 12989 26871 13047 26877
rect 13354 26868 13360 26880
rect 13412 26868 13418 26920
rect 13446 26868 13452 26920
rect 13504 26868 13510 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13556 26880 13737 26908
rect 2044 26862 2096 26868
rect 12894 26840 12900 26852
rect 9324 26812 12900 26840
rect 9324 26784 9352 26812
rect 12894 26800 12900 26812
rect 12952 26840 12958 26852
rect 13556 26840 13584 26880
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 14001 26911 14059 26917
rect 14001 26877 14013 26911
rect 14047 26908 14059 26911
rect 15856 26908 15884 27004
rect 16758 26936 16764 26988
rect 16816 26976 16822 26988
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16816 26948 16865 26976
rect 16816 26936 16822 26948
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 17862 26936 17868 26988
rect 17920 26936 17926 26988
rect 20070 26936 20076 26988
rect 20128 26976 20134 26988
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 20128 26948 21833 26976
rect 20128 26936 20134 26948
rect 21821 26945 21833 26948
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 22095 26979 22153 26985
rect 22095 26945 22107 26979
rect 22141 26976 22153 26979
rect 23014 26976 23020 26988
rect 22141 26948 23020 26976
rect 22141 26945 22153 26948
rect 22095 26939 22153 26945
rect 23014 26936 23020 26948
rect 23072 26936 23078 26988
rect 23492 26985 23520 27016
rect 23477 26979 23535 26985
rect 23477 26945 23489 26979
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 23750 26936 23756 26988
rect 23808 26936 23814 26988
rect 24228 26985 24256 27016
rect 24121 26979 24179 26985
rect 24121 26945 24133 26979
rect 24167 26945 24179 26979
rect 24121 26939 24179 26945
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26945 24271 26979
rect 24213 26939 24271 26945
rect 16574 26908 16580 26920
rect 14047 26880 14504 26908
rect 15856 26880 16580 26908
rect 14047 26877 14059 26880
rect 14001 26871 14059 26877
rect 12952 26812 13584 26840
rect 14476 26840 14504 26880
rect 16574 26868 16580 26880
rect 16632 26908 16638 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 16632 26880 16681 26908
rect 16632 26868 16638 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 16942 26868 16948 26920
rect 17000 26868 17006 26920
rect 17218 26868 17224 26920
rect 17276 26908 17282 26920
rect 17770 26917 17776 26920
rect 17313 26911 17371 26917
rect 17313 26908 17325 26911
rect 17276 26880 17325 26908
rect 17276 26868 17282 26880
rect 17313 26877 17325 26880
rect 17359 26877 17371 26911
rect 17589 26911 17647 26917
rect 17589 26908 17601 26911
rect 17313 26871 17371 26877
rect 17420 26880 17601 26908
rect 16960 26840 16988 26868
rect 17126 26840 17132 26852
rect 14476 26812 14654 26840
rect 16960 26812 17132 26840
rect 12952 26800 12958 26812
rect 3234 26732 3240 26784
rect 3292 26772 3298 26784
rect 8018 26772 8024 26784
rect 3292 26744 8024 26772
rect 3292 26732 3298 26744
rect 8018 26732 8024 26744
rect 8076 26732 8082 26784
rect 9306 26732 9312 26784
rect 9364 26732 9370 26784
rect 14626 26772 14654 26812
rect 17126 26800 17132 26812
rect 17184 26840 17190 26852
rect 17420 26840 17448 26880
rect 17589 26877 17601 26880
rect 17635 26877 17647 26911
rect 17589 26871 17647 26877
rect 17727 26911 17776 26917
rect 17727 26877 17739 26911
rect 17773 26877 17776 26911
rect 17727 26871 17776 26877
rect 17770 26868 17776 26871
rect 17828 26868 17834 26920
rect 21082 26868 21088 26920
rect 21140 26908 21146 26920
rect 21542 26908 21548 26920
rect 21140 26880 21548 26908
rect 21140 26868 21146 26880
rect 21542 26868 21548 26880
rect 21600 26868 21606 26920
rect 24136 26908 24164 26939
rect 24854 26936 24860 26988
rect 24912 26976 24918 26988
rect 25590 26976 25596 26988
rect 24912 26948 25596 26976
rect 24912 26936 24918 26948
rect 25590 26936 25596 26948
rect 25648 26936 25654 26988
rect 23584 26880 24164 26908
rect 23584 26849 23612 26880
rect 17184 26812 17448 26840
rect 23569 26843 23627 26849
rect 17184 26800 17190 26812
rect 23569 26809 23581 26843
rect 23615 26809 23627 26843
rect 23569 26803 23627 26809
rect 15749 26775 15807 26781
rect 15749 26772 15761 26775
rect 14626 26744 15761 26772
rect 15749 26741 15761 26744
rect 15795 26741 15807 26775
rect 15749 26735 15807 26741
rect 18509 26775 18567 26781
rect 18509 26741 18521 26775
rect 18555 26772 18567 26775
rect 19426 26772 19432 26784
rect 18555 26744 19432 26772
rect 18555 26741 18567 26744
rect 18509 26735 18567 26741
rect 19426 26732 19432 26744
rect 19484 26732 19490 26784
rect 22922 26732 22928 26784
rect 22980 26772 22986 26784
rect 24118 26772 24124 26784
rect 22980 26744 24124 26772
rect 22980 26732 22986 26744
rect 24118 26732 24124 26744
rect 24176 26732 24182 26784
rect 24394 26732 24400 26784
rect 24452 26732 24458 26784
rect 1104 26682 24840 26704
rect 1104 26630 3917 26682
rect 3969 26630 3981 26682
rect 4033 26630 4045 26682
rect 4097 26630 4109 26682
rect 4161 26630 4173 26682
rect 4225 26630 9851 26682
rect 9903 26630 9915 26682
rect 9967 26630 9979 26682
rect 10031 26630 10043 26682
rect 10095 26630 10107 26682
rect 10159 26630 15785 26682
rect 15837 26630 15849 26682
rect 15901 26630 15913 26682
rect 15965 26630 15977 26682
rect 16029 26630 16041 26682
rect 16093 26630 21719 26682
rect 21771 26630 21783 26682
rect 21835 26630 21847 26682
rect 21899 26630 21911 26682
rect 21963 26630 21975 26682
rect 22027 26630 24840 26682
rect 1104 26608 24840 26630
rect 2406 26528 2412 26580
rect 2464 26568 2470 26580
rect 2593 26571 2651 26577
rect 2593 26568 2605 26571
rect 2464 26540 2605 26568
rect 2464 26528 2470 26540
rect 2593 26537 2605 26540
rect 2639 26537 2651 26571
rect 2593 26531 2651 26537
rect 3237 26571 3295 26577
rect 3237 26537 3249 26571
rect 3283 26568 3295 26571
rect 3510 26568 3516 26580
rect 3283 26540 3516 26568
rect 3283 26537 3295 26540
rect 3237 26531 3295 26537
rect 3510 26528 3516 26540
rect 3568 26528 3574 26580
rect 3973 26571 4031 26577
rect 3973 26537 3985 26571
rect 4019 26568 4031 26571
rect 8662 26568 8668 26580
rect 4019 26540 8668 26568
rect 4019 26537 4031 26540
rect 3973 26531 4031 26537
rect 8662 26528 8668 26540
rect 8720 26528 8726 26580
rect 9232 26540 10824 26568
rect 3145 26503 3203 26509
rect 3145 26469 3157 26503
rect 3191 26469 3203 26503
rect 3145 26463 3203 26469
rect 1394 26392 1400 26444
rect 1452 26432 1458 26444
rect 1581 26435 1639 26441
rect 1581 26432 1593 26435
rect 1452 26404 1593 26432
rect 1452 26392 1458 26404
rect 1581 26401 1593 26404
rect 1627 26401 1639 26435
rect 1581 26395 1639 26401
rect 1839 26337 1897 26343
rect 1839 26303 1851 26337
rect 1885 26334 1897 26337
rect 1885 26303 1900 26334
rect 2866 26324 2872 26376
rect 2924 26364 2930 26376
rect 2961 26367 3019 26373
rect 2961 26364 2973 26367
rect 2924 26336 2973 26364
rect 2924 26324 2930 26336
rect 2961 26333 2973 26336
rect 3007 26333 3019 26367
rect 3160 26364 3188 26463
rect 3510 26392 3516 26444
rect 3568 26432 3574 26444
rect 4246 26432 4252 26444
rect 3568 26404 4252 26432
rect 3568 26392 3574 26404
rect 4246 26392 4252 26404
rect 4304 26392 4310 26444
rect 4522 26392 4528 26444
rect 4580 26432 4586 26444
rect 6546 26432 6552 26444
rect 4580 26404 6552 26432
rect 4580 26392 4586 26404
rect 6546 26392 6552 26404
rect 6604 26392 6610 26444
rect 9232 26441 9260 26540
rect 9674 26460 9680 26512
rect 9732 26500 9738 26512
rect 9861 26503 9919 26509
rect 9861 26500 9873 26503
rect 9732 26472 9873 26500
rect 9732 26460 9738 26472
rect 9861 26469 9873 26472
rect 9907 26469 9919 26503
rect 9861 26463 9919 26469
rect 9217 26435 9275 26441
rect 9217 26401 9229 26435
rect 9263 26401 9275 26435
rect 9217 26395 9275 26401
rect 9950 26392 9956 26444
rect 10008 26432 10014 26444
rect 10254 26435 10312 26441
rect 10254 26432 10266 26435
rect 10008 26404 10266 26432
rect 10008 26392 10014 26404
rect 10254 26401 10266 26404
rect 10300 26401 10312 26435
rect 10796 26432 10824 26540
rect 10962 26528 10968 26580
rect 11020 26568 11026 26580
rect 11057 26571 11115 26577
rect 11057 26568 11069 26571
rect 11020 26540 11069 26568
rect 11020 26528 11026 26540
rect 11057 26537 11069 26540
rect 11103 26537 11115 26571
rect 16298 26568 16304 26580
rect 11057 26531 11115 26537
rect 15580 26540 16304 26568
rect 10796 26404 11008 26432
rect 10254 26395 10312 26401
rect 3160 26336 3372 26364
rect 2961 26327 3019 26333
rect 1839 26297 1900 26303
rect 1872 26296 1900 26297
rect 3234 26296 3240 26308
rect 1872 26268 3240 26296
rect 3234 26256 3240 26268
rect 3292 26256 3298 26308
rect 3344 26296 3372 26336
rect 3418 26324 3424 26376
rect 3476 26324 3482 26376
rect 3786 26324 3792 26376
rect 3844 26324 3850 26376
rect 6730 26324 6736 26376
rect 6788 26364 6794 26376
rect 6823 26367 6881 26373
rect 6823 26364 6835 26367
rect 6788 26336 6835 26364
rect 6788 26324 6794 26336
rect 6823 26333 6835 26336
rect 6869 26333 6881 26367
rect 6823 26327 6881 26333
rect 7466 26324 7472 26376
rect 7524 26364 7530 26376
rect 8202 26364 8208 26376
rect 7524 26336 8208 26364
rect 7524 26324 7530 26336
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 9306 26324 9312 26376
rect 9364 26364 9370 26376
rect 9401 26367 9459 26373
rect 9401 26364 9413 26367
rect 9364 26336 9413 26364
rect 9364 26324 9370 26336
rect 9401 26333 9413 26336
rect 9447 26333 9459 26367
rect 9401 26327 9459 26333
rect 10134 26324 10140 26376
rect 10192 26324 10198 26376
rect 10410 26324 10416 26376
rect 10468 26324 10474 26376
rect 10980 26364 11008 26404
rect 11054 26392 11060 26444
rect 11112 26432 11118 26444
rect 11112 26404 11362 26432
rect 11112 26392 11118 26404
rect 11790 26364 11796 26376
rect 10980 26336 11796 26364
rect 11790 26324 11796 26336
rect 11848 26324 11854 26376
rect 11882 26324 11888 26376
rect 11940 26324 11946 26376
rect 13906 26324 13912 26376
rect 13964 26364 13970 26376
rect 14090 26364 14096 26376
rect 13964 26336 14096 26364
rect 13964 26324 13970 26336
rect 14090 26324 14096 26336
rect 14148 26364 14154 26376
rect 14921 26367 14979 26373
rect 14921 26364 14933 26367
rect 14148 26336 14933 26364
rect 14148 26324 14154 26336
rect 14921 26333 14933 26336
rect 14967 26333 14979 26367
rect 14921 26327 14979 26333
rect 15194 26324 15200 26376
rect 15252 26364 15258 26376
rect 15580 26364 15608 26540
rect 16298 26528 16304 26540
rect 16356 26528 16362 26580
rect 16761 26571 16819 26577
rect 16761 26537 16773 26571
rect 16807 26568 16819 26571
rect 19702 26568 19708 26580
rect 16807 26540 19708 26568
rect 16807 26537 16819 26540
rect 16761 26531 16819 26537
rect 19702 26528 19708 26540
rect 19760 26528 19766 26580
rect 22741 26571 22799 26577
rect 22741 26537 22753 26571
rect 22787 26568 22799 26571
rect 23750 26568 23756 26580
rect 22787 26540 23756 26568
rect 22787 26537 22799 26540
rect 22741 26531 22799 26537
rect 23750 26528 23756 26540
rect 23808 26528 23814 26580
rect 15930 26460 15936 26512
rect 15988 26500 15994 26512
rect 19061 26503 19119 26509
rect 15988 26472 16344 26500
rect 15988 26460 15994 26472
rect 16316 26441 16344 26472
rect 19061 26469 19073 26503
rect 19107 26500 19119 26503
rect 19518 26500 19524 26512
rect 19107 26472 19524 26500
rect 19107 26469 19119 26472
rect 19061 26463 19119 26469
rect 19518 26460 19524 26472
rect 19576 26460 19582 26512
rect 20438 26460 20444 26512
rect 20496 26500 20502 26512
rect 20496 26472 22094 26500
rect 20496 26460 20502 26472
rect 16301 26435 16359 26441
rect 16301 26401 16313 26435
rect 16347 26401 16359 26435
rect 16301 26395 16359 26401
rect 17678 26392 17684 26444
rect 17736 26392 17742 26444
rect 22066 26432 22094 26472
rect 23566 26460 23572 26512
rect 23624 26500 23630 26512
rect 24486 26500 24492 26512
rect 23624 26472 24492 26500
rect 23624 26460 23630 26472
rect 24486 26460 24492 26472
rect 24544 26460 24550 26512
rect 24854 26460 24860 26512
rect 24912 26460 24918 26512
rect 24872 26432 24900 26460
rect 22066 26404 24900 26432
rect 15252 26336 15608 26364
rect 15252 26324 15258 26336
rect 15654 26324 15660 26376
rect 15712 26364 15718 26376
rect 16485 26367 16543 26373
rect 16485 26364 16497 26367
rect 15712 26336 16497 26364
rect 15712 26324 15718 26336
rect 16485 26333 16497 26336
rect 16531 26333 16543 26367
rect 17948 26367 18006 26373
rect 16485 26327 16543 26333
rect 16776 26336 17908 26364
rect 12158 26296 12164 26308
rect 3344 26268 9444 26296
rect 5350 26188 5356 26240
rect 5408 26228 5414 26240
rect 5810 26228 5816 26240
rect 5408 26200 5816 26228
rect 5408 26188 5414 26200
rect 5810 26188 5816 26200
rect 5868 26188 5874 26240
rect 7561 26231 7619 26237
rect 7561 26197 7573 26231
rect 7607 26228 7619 26231
rect 7650 26228 7656 26240
rect 7607 26200 7656 26228
rect 7607 26197 7619 26200
rect 7561 26191 7619 26197
rect 7650 26188 7656 26200
rect 7708 26188 7714 26240
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 8294 26228 8300 26240
rect 7800 26200 8300 26228
rect 7800 26188 7806 26200
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 9416 26228 9444 26268
rect 10888 26268 12164 26296
rect 10888 26228 10916 26268
rect 12158 26256 12164 26268
rect 12216 26296 12222 26308
rect 12253 26299 12311 26305
rect 12253 26296 12265 26299
rect 12216 26268 12265 26296
rect 12216 26256 12222 26268
rect 12253 26265 12265 26268
rect 12299 26265 12311 26299
rect 16776 26296 16804 26336
rect 12253 26259 12311 26265
rect 12820 26268 16804 26296
rect 9416 26200 10916 26228
rect 10962 26188 10968 26240
rect 11020 26228 11026 26240
rect 11422 26228 11428 26240
rect 11020 26200 11428 26228
rect 11020 26188 11026 26200
rect 11422 26188 11428 26200
rect 11480 26228 11486 26240
rect 11517 26231 11575 26237
rect 11517 26228 11529 26231
rect 11480 26200 11529 26228
rect 11480 26188 11486 26200
rect 11517 26197 11529 26200
rect 11563 26197 11575 26231
rect 11517 26191 11575 26197
rect 12618 26188 12624 26240
rect 12676 26188 12682 26240
rect 12820 26237 12848 26268
rect 16850 26256 16856 26308
rect 16908 26256 16914 26308
rect 17880 26296 17908 26336
rect 17948 26333 17960 26367
rect 17994 26364 18006 26367
rect 19426 26364 19432 26376
rect 17994 26336 19432 26364
rect 17994 26333 18006 26336
rect 17948 26327 18006 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 20530 26324 20536 26376
rect 20588 26324 20594 26376
rect 20714 26324 20720 26376
rect 20772 26364 20778 26376
rect 22925 26367 22983 26373
rect 22925 26364 22937 26367
rect 20772 26336 22937 26364
rect 20772 26324 20778 26336
rect 22925 26333 22937 26336
rect 22971 26333 22983 26367
rect 22925 26327 22983 26333
rect 23474 26324 23480 26376
rect 23532 26324 23538 26376
rect 23566 26324 23572 26376
rect 23624 26364 23630 26376
rect 23661 26367 23719 26373
rect 23661 26364 23673 26367
rect 23624 26336 23673 26364
rect 23624 26324 23630 26336
rect 23661 26333 23673 26336
rect 23707 26333 23719 26367
rect 23661 26327 23719 26333
rect 19610 26296 19616 26308
rect 17880 26268 19616 26296
rect 19610 26256 19616 26268
rect 19668 26256 19674 26308
rect 20548 26296 20576 26324
rect 23845 26299 23903 26305
rect 23845 26296 23857 26299
rect 20548 26268 23857 26296
rect 23845 26265 23857 26268
rect 23891 26265 23903 26299
rect 23845 26259 23903 26265
rect 24213 26299 24271 26305
rect 24213 26265 24225 26299
rect 24259 26296 24271 26299
rect 25130 26296 25136 26308
rect 24259 26268 25136 26296
rect 24259 26265 24271 26268
rect 24213 26259 24271 26265
rect 25130 26256 25136 26268
rect 25188 26256 25194 26308
rect 12805 26231 12863 26237
rect 12805 26197 12817 26231
rect 12851 26197 12863 26231
rect 12805 26191 12863 26197
rect 12894 26188 12900 26240
rect 12952 26228 12958 26240
rect 13262 26228 13268 26240
rect 12952 26200 13268 26228
rect 12952 26188 12958 26200
rect 13262 26188 13268 26200
rect 13320 26188 13326 26240
rect 14826 26188 14832 26240
rect 14884 26228 14890 26240
rect 16114 26228 16120 26240
rect 14884 26200 16120 26228
rect 14884 26188 14890 26200
rect 16114 26188 16120 26200
rect 16172 26188 16178 26240
rect 19242 26188 19248 26240
rect 19300 26188 19306 26240
rect 23658 26188 23664 26240
rect 23716 26188 23722 26240
rect 1104 26138 25000 26160
rect 1104 26086 6884 26138
rect 6936 26086 6948 26138
rect 7000 26086 7012 26138
rect 7064 26086 7076 26138
rect 7128 26086 7140 26138
rect 7192 26086 12818 26138
rect 12870 26086 12882 26138
rect 12934 26086 12946 26138
rect 12998 26086 13010 26138
rect 13062 26086 13074 26138
rect 13126 26086 18752 26138
rect 18804 26086 18816 26138
rect 18868 26086 18880 26138
rect 18932 26086 18944 26138
rect 18996 26086 19008 26138
rect 19060 26086 24686 26138
rect 24738 26086 24750 26138
rect 24802 26086 24814 26138
rect 24866 26086 24878 26138
rect 24930 26086 24942 26138
rect 24994 26086 25000 26138
rect 1104 26064 25000 26086
rect 2406 25984 2412 26036
rect 2464 26024 2470 26036
rect 2501 26027 2559 26033
rect 2501 26024 2513 26027
rect 2464 25996 2513 26024
rect 2464 25984 2470 25996
rect 2501 25993 2513 25996
rect 2547 25993 2559 26027
rect 2501 25987 2559 25993
rect 3053 26027 3111 26033
rect 3053 25993 3065 26027
rect 3099 26024 3111 26027
rect 3329 26027 3387 26033
rect 3099 25996 3280 26024
rect 3099 25993 3111 25996
rect 3053 25987 3111 25993
rect 1302 25916 1308 25968
rect 1360 25956 1366 25968
rect 3252 25956 3280 25996
rect 3329 25993 3341 26027
rect 3375 26024 3387 26027
rect 11606 26024 11612 26036
rect 3375 25996 8616 26024
rect 3375 25993 3387 25996
rect 3329 25987 3387 25993
rect 5994 25956 6000 25968
rect 1360 25928 3188 25956
rect 3252 25928 6000 25956
rect 1360 25916 1366 25928
rect 1394 25848 1400 25900
rect 1452 25888 1458 25900
rect 1489 25891 1547 25897
rect 1489 25888 1501 25891
rect 1452 25860 1501 25888
rect 1452 25848 1458 25860
rect 1489 25857 1501 25860
rect 1535 25857 1547 25891
rect 1489 25851 1547 25857
rect 1763 25891 1821 25897
rect 1763 25857 1775 25891
rect 1809 25888 1821 25891
rect 2774 25888 2780 25900
rect 1809 25860 2780 25888
rect 1809 25857 1821 25860
rect 1763 25851 1821 25857
rect 2774 25848 2780 25860
rect 2832 25848 2838 25900
rect 3160 25897 3188 25928
rect 5994 25916 6000 25928
rect 6052 25916 6058 25968
rect 7101 25959 7159 25965
rect 6840 25928 7052 25956
rect 2869 25891 2927 25897
rect 2869 25857 2881 25891
rect 2915 25857 2927 25891
rect 2869 25851 2927 25857
rect 3145 25891 3203 25897
rect 3145 25857 3157 25891
rect 3191 25857 3203 25891
rect 3145 25851 3203 25857
rect 3695 25891 3753 25897
rect 3695 25857 3707 25891
rect 3741 25888 3753 25891
rect 4246 25888 4252 25900
rect 3741 25860 4252 25888
rect 3741 25857 3753 25860
rect 3695 25851 3753 25857
rect 2884 25752 2912 25851
rect 4246 25848 4252 25860
rect 4304 25848 4310 25900
rect 5075 25891 5133 25897
rect 5075 25857 5087 25891
rect 5121 25888 5133 25891
rect 6270 25888 6276 25900
rect 5121 25860 6276 25888
rect 5121 25857 5133 25860
rect 5075 25851 5133 25857
rect 6270 25848 6276 25860
rect 6328 25848 6334 25900
rect 6840 25897 6868 25928
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25857 6883 25891
rect 7024 25888 7052 25928
rect 7101 25925 7113 25959
rect 7147 25956 7159 25959
rect 7282 25956 7288 25968
rect 7147 25928 7288 25956
rect 7147 25925 7159 25928
rect 7101 25919 7159 25925
rect 7282 25916 7288 25928
rect 7340 25956 7346 25968
rect 7650 25956 7656 25968
rect 7340 25928 7656 25956
rect 7340 25916 7346 25928
rect 7650 25916 7656 25928
rect 7708 25916 7714 25968
rect 7834 25916 7840 25968
rect 7892 25916 7898 25968
rect 8202 25916 8208 25968
rect 8260 25916 8266 25968
rect 7377 25891 7435 25897
rect 7377 25888 7389 25891
rect 7024 25860 7389 25888
rect 6825 25851 6883 25857
rect 7377 25857 7389 25860
rect 7423 25857 7435 25891
rect 7377 25851 7435 25857
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25888 7527 25891
rect 7742 25888 7748 25900
rect 7515 25860 7748 25888
rect 7515 25857 7527 25860
rect 7469 25851 7527 25857
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 3421 25823 3479 25829
rect 3421 25789 3433 25823
rect 3467 25789 3479 25823
rect 3421 25783 3479 25789
rect 4801 25823 4859 25829
rect 4801 25789 4813 25823
rect 4847 25789 4859 25823
rect 4801 25783 4859 25789
rect 2148 25724 2912 25752
rect 1210 25644 1216 25696
rect 1268 25684 1274 25696
rect 2148 25684 2176 25724
rect 1268 25656 2176 25684
rect 1268 25644 1274 25656
rect 2222 25644 2228 25696
rect 2280 25684 2286 25696
rect 2590 25684 2596 25696
rect 2280 25656 2596 25684
rect 2280 25644 2286 25656
rect 2590 25644 2596 25656
rect 2648 25644 2654 25696
rect 2774 25644 2780 25696
rect 2832 25684 2838 25696
rect 3142 25684 3148 25696
rect 2832 25656 3148 25684
rect 2832 25644 2838 25656
rect 3142 25644 3148 25656
rect 3200 25644 3206 25696
rect 3436 25684 3464 25783
rect 3694 25684 3700 25696
rect 3436 25656 3700 25684
rect 3694 25644 3700 25656
rect 3752 25644 3758 25696
rect 4430 25644 4436 25696
rect 4488 25644 4494 25696
rect 4816 25684 4844 25783
rect 7558 25780 7564 25832
rect 7616 25780 7622 25832
rect 5258 25684 5264 25696
rect 4816 25656 5264 25684
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 5810 25644 5816 25696
rect 5868 25644 5874 25696
rect 8386 25644 8392 25696
rect 8444 25644 8450 25696
rect 8588 25684 8616 25996
rect 9048 25996 11612 26024
rect 8754 25780 8760 25832
rect 8812 25820 8818 25832
rect 9048 25829 9076 25996
rect 11606 25984 11612 25996
rect 11664 25984 11670 26036
rect 11790 25984 11796 26036
rect 11848 25984 11854 26036
rect 11882 25984 11888 26036
rect 11940 26024 11946 26036
rect 14826 26024 14832 26036
rect 11940 25996 14832 26024
rect 11940 25984 11946 25996
rect 14826 25984 14832 25996
rect 14884 25984 14890 26036
rect 15010 25984 15016 26036
rect 15068 25984 15074 26036
rect 15654 25984 15660 26036
rect 15712 25984 15718 26036
rect 15930 25984 15936 26036
rect 15988 25984 15994 26036
rect 16025 26027 16083 26033
rect 16025 25993 16037 26027
rect 16071 26024 16083 26027
rect 16850 26024 16856 26036
rect 16071 25996 16856 26024
rect 16071 25993 16083 25996
rect 16025 25987 16083 25993
rect 16850 25984 16856 25996
rect 16908 25984 16914 26036
rect 22373 26027 22431 26033
rect 22373 25993 22385 26027
rect 22419 25993 22431 26027
rect 22373 25987 22431 25993
rect 23477 26027 23535 26033
rect 23477 25993 23489 26027
rect 23523 26024 23535 26027
rect 23566 26024 23572 26036
rect 23523 25996 23572 26024
rect 23523 25993 23535 25996
rect 23477 25987 23535 25993
rect 11808 25956 11836 25984
rect 15028 25956 15056 25984
rect 11808 25928 13124 25956
rect 15028 25928 15608 25956
rect 11514 25848 11520 25900
rect 11572 25848 11578 25900
rect 11791 25891 11849 25897
rect 11791 25857 11803 25891
rect 11837 25888 11849 25891
rect 12250 25888 12256 25900
rect 11837 25860 12256 25888
rect 11837 25857 11849 25860
rect 11791 25851 11849 25857
rect 12250 25848 12256 25860
rect 12308 25848 12314 25900
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 8812 25792 9045 25820
rect 8812 25780 8818 25792
rect 9033 25789 9045 25792
rect 9079 25789 9091 25823
rect 9033 25783 9091 25789
rect 9217 25823 9275 25829
rect 9217 25789 9229 25823
rect 9263 25820 9275 25823
rect 9582 25820 9588 25832
rect 9263 25792 9588 25820
rect 9263 25789 9275 25792
rect 9217 25783 9275 25789
rect 9582 25780 9588 25792
rect 9640 25780 9646 25832
rect 9766 25780 9772 25832
rect 9824 25820 9830 25832
rect 9953 25823 10011 25829
rect 9953 25820 9965 25823
rect 9824 25792 9965 25820
rect 9824 25780 9830 25792
rect 9953 25789 9965 25792
rect 9999 25789 10011 25823
rect 9953 25783 10011 25789
rect 10042 25780 10048 25832
rect 10100 25829 10106 25832
rect 10100 25823 10128 25829
rect 10116 25789 10128 25823
rect 10100 25783 10128 25789
rect 10229 25823 10287 25829
rect 10229 25789 10241 25823
rect 10275 25820 10287 25823
rect 10410 25820 10416 25832
rect 10275 25792 10416 25820
rect 10275 25789 10287 25792
rect 10229 25783 10287 25789
rect 10100 25780 10106 25783
rect 10410 25780 10416 25792
rect 10468 25780 10474 25832
rect 13096 25829 13124 25928
rect 13262 25848 13268 25900
rect 13320 25848 13326 25900
rect 13998 25848 14004 25900
rect 14056 25848 14062 25900
rect 14274 25848 14280 25900
rect 14332 25848 14338 25900
rect 15580 25897 15608 25928
rect 14921 25891 14979 25897
rect 14921 25857 14933 25891
rect 14967 25888 14979 25891
rect 15473 25891 15531 25897
rect 15473 25888 15485 25891
rect 14967 25860 15485 25888
rect 14967 25857 14979 25860
rect 14921 25851 14979 25857
rect 15473 25857 15485 25860
rect 15519 25857 15531 25891
rect 15473 25851 15531 25857
rect 15565 25891 15623 25897
rect 15565 25857 15577 25891
rect 15611 25857 15623 25891
rect 15565 25851 15623 25857
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25888 15899 25891
rect 15948 25888 15976 25984
rect 17126 25916 17132 25968
rect 17184 25956 17190 25968
rect 20714 25956 20720 25968
rect 17184 25928 20720 25956
rect 17184 25916 17190 25928
rect 20714 25916 20720 25928
rect 20772 25916 20778 25968
rect 22388 25956 22416 25987
rect 23566 25984 23572 25996
rect 23624 25984 23630 26036
rect 23937 26027 23995 26033
rect 23937 25993 23949 26027
rect 23983 26024 23995 26027
rect 24302 26024 24308 26036
rect 23983 25996 24308 26024
rect 23983 25993 23995 25996
rect 23937 25987 23995 25993
rect 24302 25984 24308 25996
rect 24360 25984 24366 26036
rect 22388 25928 23060 25956
rect 15887 25860 15976 25888
rect 16025 25891 16083 25897
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16025 25857 16037 25891
rect 16071 25857 16083 25891
rect 16025 25851 16083 25857
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25820 13139 25823
rect 13127 25792 13308 25820
rect 13127 25789 13139 25792
rect 13081 25783 13139 25789
rect 9674 25712 9680 25764
rect 9732 25712 9738 25764
rect 10686 25712 10692 25764
rect 10744 25752 10750 25764
rect 10873 25755 10931 25761
rect 10873 25752 10885 25755
rect 10744 25724 10885 25752
rect 10744 25712 10750 25724
rect 10873 25721 10885 25724
rect 10919 25721 10931 25755
rect 12986 25752 12992 25764
rect 10873 25715 10931 25721
rect 12406 25724 12992 25752
rect 12406 25684 12434 25724
rect 12986 25712 12992 25724
rect 13044 25712 13050 25764
rect 13280 25696 13308 25792
rect 13722 25780 13728 25832
rect 13780 25780 13786 25832
rect 14139 25823 14197 25829
rect 14139 25789 14151 25823
rect 14185 25820 14197 25823
rect 16040 25820 16068 25851
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18843 25891 18901 25897
rect 18843 25888 18855 25891
rect 18012 25860 18855 25888
rect 18012 25848 18018 25860
rect 18843 25857 18855 25860
rect 18889 25857 18901 25891
rect 19981 25891 20039 25897
rect 19981 25888 19993 25891
rect 18843 25851 18901 25857
rect 19628 25860 19993 25888
rect 14185 25792 14688 25820
rect 14185 25789 14197 25792
rect 14139 25783 14197 25789
rect 8588 25656 12434 25684
rect 12526 25644 12532 25696
rect 12584 25644 12590 25696
rect 13262 25644 13268 25696
rect 13320 25644 13326 25696
rect 13446 25644 13452 25696
rect 13504 25684 13510 25696
rect 14660 25684 14688 25792
rect 15304 25792 16068 25820
rect 15304 25761 15332 25792
rect 16114 25780 16120 25832
rect 16172 25820 16178 25832
rect 16482 25820 16488 25832
rect 16172 25792 16488 25820
rect 16172 25780 16178 25792
rect 16482 25780 16488 25792
rect 16540 25780 16546 25832
rect 18601 25823 18659 25829
rect 18601 25789 18613 25823
rect 18647 25789 18659 25823
rect 18601 25783 18659 25789
rect 15289 25755 15347 25761
rect 15289 25721 15301 25755
rect 15335 25721 15347 25755
rect 15289 25715 15347 25721
rect 15654 25712 15660 25764
rect 15712 25752 15718 25764
rect 16666 25752 16672 25764
rect 15712 25724 16672 25752
rect 15712 25712 15718 25724
rect 16666 25712 16672 25724
rect 16724 25712 16730 25764
rect 18616 25752 18644 25783
rect 19628 25761 19656 25860
rect 19981 25857 19993 25860
rect 20027 25888 20039 25891
rect 20349 25891 20407 25897
rect 20349 25888 20361 25891
rect 20027 25860 20361 25888
rect 20027 25857 20039 25860
rect 19981 25851 20039 25857
rect 20349 25857 20361 25860
rect 20395 25857 20407 25891
rect 20349 25851 20407 25857
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25857 20591 25891
rect 20533 25851 20591 25857
rect 20257 25823 20315 25829
rect 20257 25789 20269 25823
rect 20303 25820 20315 25823
rect 20441 25823 20499 25829
rect 20441 25820 20453 25823
rect 20303 25792 20453 25820
rect 20303 25789 20315 25792
rect 20257 25783 20315 25789
rect 20441 25789 20453 25792
rect 20487 25789 20499 25823
rect 20441 25783 20499 25789
rect 19613 25755 19671 25761
rect 18616 25724 18736 25752
rect 13504 25656 14688 25684
rect 13504 25644 13510 25656
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 17402 25684 17408 25696
rect 14884 25656 17408 25684
rect 14884 25644 14890 25656
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 18708 25684 18736 25724
rect 19613 25721 19625 25755
rect 19659 25721 19671 25755
rect 19613 25715 19671 25721
rect 20346 25712 20352 25764
rect 20404 25752 20410 25764
rect 20548 25752 20576 25851
rect 21358 25848 21364 25900
rect 21416 25848 21422 25900
rect 21542 25848 21548 25900
rect 21600 25848 21606 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 23032 25897 23060 25928
rect 23842 25916 23848 25968
rect 23900 25956 23906 25968
rect 24121 25959 24179 25965
rect 24121 25956 24133 25959
rect 23900 25928 24133 25956
rect 23900 25916 23906 25928
rect 24121 25925 24133 25928
rect 24167 25925 24179 25959
rect 24121 25919 24179 25925
rect 22557 25891 22615 25897
rect 22557 25888 22569 25891
rect 22152 25860 22569 25888
rect 22152 25848 22158 25860
rect 22557 25857 22569 25860
rect 22603 25857 22615 25891
rect 22557 25851 22615 25857
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25857 23075 25891
rect 23017 25851 23075 25857
rect 23566 25848 23572 25900
rect 23624 25888 23630 25900
rect 23661 25891 23719 25897
rect 23661 25888 23673 25891
rect 23624 25860 23673 25888
rect 23624 25848 23630 25860
rect 23661 25857 23673 25860
rect 23707 25857 23719 25891
rect 23661 25851 23719 25857
rect 23753 25891 23811 25897
rect 23753 25857 23765 25891
rect 23799 25857 23811 25891
rect 23753 25851 23811 25857
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 23768 25820 23796 25851
rect 23440 25792 23796 25820
rect 23440 25780 23446 25792
rect 20404 25724 20576 25752
rect 20404 25712 20410 25724
rect 19426 25684 19432 25696
rect 18708 25656 19432 25684
rect 19426 25644 19432 25656
rect 19484 25684 19490 25696
rect 19978 25684 19984 25696
rect 19484 25656 19984 25684
rect 19484 25644 19490 25656
rect 19978 25644 19984 25656
rect 20036 25644 20042 25696
rect 20070 25644 20076 25696
rect 20128 25644 20134 25696
rect 20165 25687 20223 25693
rect 20165 25653 20177 25687
rect 20211 25684 20223 25687
rect 21082 25684 21088 25696
rect 20211 25656 21088 25684
rect 20211 25653 20223 25656
rect 20165 25647 20223 25653
rect 21082 25644 21088 25656
rect 21140 25644 21146 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 23106 25644 23112 25696
rect 23164 25644 23170 25696
rect 24394 25644 24400 25696
rect 24452 25644 24458 25696
rect 1104 25594 24840 25616
rect 1104 25542 3917 25594
rect 3969 25542 3981 25594
rect 4033 25542 4045 25594
rect 4097 25542 4109 25594
rect 4161 25542 4173 25594
rect 4225 25542 9851 25594
rect 9903 25542 9915 25594
rect 9967 25542 9979 25594
rect 10031 25542 10043 25594
rect 10095 25542 10107 25594
rect 10159 25542 15785 25594
rect 15837 25542 15849 25594
rect 15901 25542 15913 25594
rect 15965 25542 15977 25594
rect 16029 25542 16041 25594
rect 16093 25542 21719 25594
rect 21771 25542 21783 25594
rect 21835 25542 21847 25594
rect 21899 25542 21911 25594
rect 21963 25542 21975 25594
rect 22027 25542 24840 25594
rect 1104 25520 24840 25542
rect 1581 25483 1639 25489
rect 1581 25449 1593 25483
rect 1627 25480 1639 25483
rect 2222 25480 2228 25492
rect 1627 25452 2228 25480
rect 1627 25449 1639 25452
rect 1581 25443 1639 25449
rect 2222 25440 2228 25452
rect 2280 25440 2286 25492
rect 2332 25452 3740 25480
rect 2332 25353 2360 25452
rect 3712 25424 3740 25452
rect 7742 25440 7748 25492
rect 7800 25480 7806 25492
rect 8297 25483 8355 25489
rect 8297 25480 8309 25483
rect 7800 25452 8309 25480
rect 7800 25440 7806 25452
rect 8297 25449 8309 25452
rect 8343 25449 8355 25483
rect 8297 25443 8355 25449
rect 8404 25452 10364 25480
rect 3329 25415 3387 25421
rect 3329 25381 3341 25415
rect 3375 25381 3387 25415
rect 3329 25375 3387 25381
rect 2317 25347 2375 25353
rect 2056 25316 2268 25344
rect 2056 25288 2084 25316
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 1670 25236 1676 25288
rect 1728 25236 1734 25288
rect 2038 25236 2044 25288
rect 2096 25236 2102 25288
rect 2130 25236 2136 25288
rect 2188 25236 2194 25288
rect 2240 25276 2268 25316
rect 2317 25313 2329 25347
rect 2363 25313 2375 25347
rect 3344 25344 3372 25375
rect 3694 25372 3700 25424
rect 3752 25372 3758 25424
rect 8404 25412 8432 25452
rect 8128 25384 8432 25412
rect 10336 25412 10364 25452
rect 10410 25440 10416 25492
rect 10468 25480 10474 25492
rect 10505 25483 10563 25489
rect 10505 25480 10517 25483
rect 10468 25452 10517 25480
rect 10468 25440 10474 25452
rect 10505 25449 10517 25452
rect 10551 25449 10563 25483
rect 10505 25443 10563 25449
rect 11146 25440 11152 25492
rect 11204 25440 11210 25492
rect 12986 25440 12992 25492
rect 13044 25440 13050 25492
rect 16574 25440 16580 25492
rect 16632 25480 16638 25492
rect 16850 25480 16856 25492
rect 16632 25452 16856 25480
rect 16632 25440 16638 25452
rect 16850 25440 16856 25452
rect 16908 25480 16914 25492
rect 19337 25483 19395 25489
rect 16908 25452 17448 25480
rect 16908 25440 16914 25452
rect 11164 25412 11192 25440
rect 10336 25384 11192 25412
rect 3344 25316 3818 25344
rect 2317 25307 2375 25313
rect 5258 25304 5264 25356
rect 5316 25344 5322 25356
rect 5445 25347 5503 25353
rect 5445 25344 5457 25347
rect 5316 25316 5457 25344
rect 5316 25304 5322 25316
rect 5445 25313 5457 25316
rect 5491 25313 5503 25347
rect 5445 25307 5503 25313
rect 2559 25279 2617 25285
rect 2559 25276 2571 25279
rect 2240 25248 2571 25276
rect 2559 25245 2571 25248
rect 2605 25245 2617 25279
rect 3510 25276 3516 25288
rect 2559 25239 2617 25245
rect 2792 25248 3516 25276
rect 2314 25168 2320 25220
rect 2372 25208 2378 25220
rect 2792 25208 2820 25248
rect 3510 25236 3516 25248
rect 3568 25236 3574 25288
rect 4709 25279 4767 25285
rect 4709 25276 4721 25279
rect 3712 25248 4721 25276
rect 2372 25180 2820 25208
rect 2372 25168 2378 25180
rect 3712 25152 3740 25248
rect 4709 25245 4721 25248
rect 4755 25245 4767 25279
rect 4709 25239 4767 25245
rect 5074 25236 5080 25288
rect 5132 25236 5138 25288
rect 4249 25211 4307 25217
rect 4249 25177 4261 25211
rect 4295 25177 4307 25211
rect 4249 25171 4307 25177
rect 4341 25211 4399 25217
rect 4341 25177 4353 25211
rect 4387 25208 4399 25211
rect 4430 25208 4436 25220
rect 4387 25180 4436 25208
rect 4387 25177 4399 25180
rect 4341 25171 4399 25177
rect 1854 25100 1860 25152
rect 1912 25100 1918 25152
rect 1949 25143 2007 25149
rect 1949 25109 1961 25143
rect 1995 25140 2007 25143
rect 3694 25140 3700 25152
rect 1995 25112 3700 25140
rect 1995 25109 2007 25112
rect 1949 25103 2007 25109
rect 3694 25100 3700 25112
rect 3752 25100 3758 25152
rect 3878 25100 3884 25152
rect 3936 25140 3942 25152
rect 3973 25143 4031 25149
rect 3973 25140 3985 25143
rect 3936 25112 3985 25140
rect 3936 25100 3942 25112
rect 3973 25109 3985 25112
rect 4019 25109 4031 25143
rect 3973 25103 4031 25109
rect 4062 25100 4068 25152
rect 4120 25140 4126 25152
rect 4264 25140 4292 25171
rect 4430 25168 4436 25180
rect 4488 25168 4494 25220
rect 5092 25149 5120 25236
rect 5460 25208 5488 25307
rect 6178 25304 6184 25356
rect 6236 25344 6242 25356
rect 6546 25344 6552 25356
rect 6236 25316 6552 25344
rect 6236 25304 6242 25316
rect 6546 25304 6552 25316
rect 6604 25344 6610 25356
rect 7285 25347 7343 25353
rect 7285 25344 7297 25347
rect 6604 25316 7297 25344
rect 6604 25304 6610 25316
rect 7285 25313 7297 25316
rect 7331 25313 7343 25347
rect 7285 25307 7343 25313
rect 5719 25279 5777 25285
rect 5719 25245 5731 25279
rect 5765 25276 5777 25279
rect 7006 25276 7012 25288
rect 5765 25248 7012 25276
rect 5765 25245 5777 25248
rect 5719 25239 5777 25245
rect 7006 25236 7012 25248
rect 7064 25236 7070 25288
rect 7300 25208 7328 25307
rect 7559 25279 7617 25285
rect 7559 25245 7571 25279
rect 7605 25276 7617 25279
rect 8018 25276 8024 25288
rect 7605 25248 8024 25276
rect 7605 25245 7617 25248
rect 7559 25239 7617 25245
rect 8018 25236 8024 25248
rect 8076 25236 8082 25288
rect 8128 25208 8156 25384
rect 12526 25344 12532 25356
rect 12466 25316 12532 25344
rect 12526 25304 12532 25316
rect 12584 25304 12590 25356
rect 13004 25344 13032 25440
rect 15378 25372 15384 25424
rect 15436 25412 15442 25424
rect 16482 25412 16488 25424
rect 15436 25384 16488 25412
rect 15436 25372 15442 25384
rect 16482 25372 16488 25384
rect 16540 25412 16546 25424
rect 16540 25384 16896 25412
rect 16540 25372 16546 25384
rect 16669 25347 16727 25353
rect 16669 25344 16681 25347
rect 13004 25316 16681 25344
rect 16669 25313 16681 25316
rect 16715 25344 16727 25347
rect 16758 25344 16764 25356
rect 16715 25316 16764 25344
rect 16715 25313 16727 25316
rect 16669 25307 16727 25313
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 16868 25353 16896 25384
rect 16853 25347 16911 25353
rect 16853 25313 16865 25347
rect 16899 25313 16911 25347
rect 16853 25307 16911 25313
rect 17310 25304 17316 25356
rect 17368 25304 17374 25356
rect 17420 25344 17448 25452
rect 19337 25449 19349 25483
rect 19383 25480 19395 25483
rect 20070 25480 20076 25492
rect 19383 25452 20076 25480
rect 19383 25449 19395 25452
rect 19337 25443 19395 25449
rect 20070 25440 20076 25452
rect 20128 25440 20134 25492
rect 20346 25440 20352 25492
rect 20404 25440 20410 25492
rect 21358 25440 21364 25492
rect 21416 25440 21422 25492
rect 23106 25440 23112 25492
rect 23164 25480 23170 25492
rect 23477 25483 23535 25489
rect 23477 25480 23489 25483
rect 23164 25452 23489 25480
rect 23164 25440 23170 25452
rect 23477 25449 23489 25452
rect 23523 25449 23535 25483
rect 23477 25443 23535 25449
rect 23566 25440 23572 25492
rect 23624 25440 23630 25492
rect 23658 25440 23664 25492
rect 23716 25440 23722 25492
rect 19518 25372 19524 25424
rect 19576 25372 19582 25424
rect 19613 25415 19671 25421
rect 19613 25381 19625 25415
rect 19659 25412 19671 25415
rect 20364 25412 20392 25440
rect 19659 25384 20392 25412
rect 23201 25415 23259 25421
rect 19659 25381 19671 25384
rect 19613 25375 19671 25381
rect 23201 25381 23213 25415
rect 23247 25412 23259 25415
rect 23584 25412 23612 25440
rect 23247 25384 23612 25412
rect 23247 25381 23259 25384
rect 23201 25375 23259 25381
rect 17706 25347 17764 25353
rect 17706 25344 17718 25347
rect 17420 25316 17718 25344
rect 17706 25313 17718 25316
rect 17752 25313 17764 25347
rect 17706 25307 17764 25313
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 8536 25248 9505 25276
rect 8536 25236 8542 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 9767 25279 9825 25285
rect 9767 25245 9779 25279
rect 9813 25276 9825 25279
rect 10318 25276 10324 25288
rect 9813 25248 10324 25276
rect 9813 25245 9825 25248
rect 9767 25239 9825 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11698 25276 11704 25288
rect 11112 25248 11704 25276
rect 11112 25236 11118 25248
rect 11698 25236 11704 25248
rect 11756 25236 11762 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25276 11851 25279
rect 12710 25276 12716 25288
rect 11839 25248 12716 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 17586 25236 17592 25288
rect 17644 25236 17650 25288
rect 17862 25236 17868 25288
rect 17920 25236 17926 25288
rect 19242 25236 19248 25288
rect 19300 25236 19306 25288
rect 19536 25276 19564 25372
rect 19978 25304 19984 25356
rect 20036 25344 20042 25356
rect 20349 25347 20407 25353
rect 20349 25344 20361 25347
rect 20036 25316 20361 25344
rect 20036 25304 20042 25316
rect 20349 25313 20361 25316
rect 20395 25313 20407 25347
rect 20349 25307 20407 25313
rect 23474 25304 23480 25356
rect 23532 25304 23538 25356
rect 23676 25353 23704 25440
rect 23661 25347 23719 25353
rect 23661 25313 23673 25347
rect 23707 25313 23719 25347
rect 23661 25307 23719 25313
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19536 25248 19809 25276
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 20070 25236 20076 25288
rect 20128 25276 20134 25288
rect 20128 25255 20650 25276
rect 20128 25249 20665 25255
rect 20128 25248 20619 25249
rect 20128 25236 20134 25248
rect 5460 25180 7236 25208
rect 7300 25180 8156 25208
rect 4120 25112 4292 25140
rect 5077 25143 5135 25149
rect 4120 25100 4126 25112
rect 5077 25109 5089 25143
rect 5123 25109 5135 25143
rect 5077 25103 5135 25109
rect 5258 25100 5264 25152
rect 5316 25100 5322 25152
rect 6362 25100 6368 25152
rect 6420 25140 6426 25152
rect 6457 25143 6515 25149
rect 6457 25140 6469 25143
rect 6420 25112 6469 25140
rect 6420 25100 6426 25112
rect 6457 25109 6469 25112
rect 6503 25109 6515 25143
rect 7208 25140 7236 25180
rect 8754 25168 8760 25220
rect 8812 25208 8818 25220
rect 8812 25180 11560 25208
rect 8812 25168 8818 25180
rect 7282 25140 7288 25152
rect 7208 25112 7288 25140
rect 6457 25103 6515 25109
rect 7282 25100 7288 25112
rect 7340 25100 7346 25152
rect 9766 25100 9772 25152
rect 9824 25140 9830 25152
rect 11054 25140 11060 25152
rect 9824 25112 11060 25140
rect 9824 25100 9830 25112
rect 11054 25100 11060 25112
rect 11112 25100 11118 25152
rect 11330 25100 11336 25152
rect 11388 25140 11394 25152
rect 11425 25143 11483 25149
rect 11425 25140 11437 25143
rect 11388 25112 11437 25140
rect 11388 25100 11394 25112
rect 11425 25109 11437 25112
rect 11471 25109 11483 25143
rect 11532 25140 11560 25180
rect 11606 25168 11612 25220
rect 11664 25208 11670 25220
rect 11664 25180 12020 25208
rect 11664 25168 11670 25180
rect 11882 25140 11888 25152
rect 11532 25112 11888 25140
rect 11425 25103 11483 25109
rect 11882 25100 11888 25112
rect 11940 25100 11946 25152
rect 11992 25140 12020 25180
rect 12158 25168 12164 25220
rect 12216 25168 12222 25220
rect 19150 25208 19156 25220
rect 18432 25180 19156 25208
rect 12529 25143 12587 25149
rect 12529 25140 12541 25143
rect 11992 25112 12541 25140
rect 12529 25109 12541 25112
rect 12575 25140 12587 25143
rect 12618 25140 12624 25152
rect 12575 25112 12624 25140
rect 12575 25109 12587 25112
rect 12529 25103 12587 25109
rect 12618 25100 12624 25112
rect 12676 25100 12682 25152
rect 12713 25143 12771 25149
rect 12713 25109 12725 25143
rect 12759 25140 12771 25143
rect 18432 25140 18460 25180
rect 19150 25168 19156 25180
rect 19208 25168 19214 25220
rect 20607 25215 20619 25248
rect 20653 25215 20665 25249
rect 21174 25236 21180 25288
rect 21232 25276 21238 25288
rect 21821 25279 21879 25285
rect 21821 25276 21833 25279
rect 21232 25248 21833 25276
rect 21232 25236 21238 25248
rect 21821 25245 21833 25248
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 22554 25236 22560 25288
rect 22612 25236 22618 25288
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25276 23443 25279
rect 23492 25276 23520 25304
rect 23431 25248 23520 25276
rect 23431 25245 23443 25248
rect 23385 25239 23443 25245
rect 20607 25209 20665 25215
rect 21726 25168 21732 25220
rect 21784 25208 21790 25220
rect 22094 25217 22100 25220
rect 22088 25208 22100 25217
rect 21784 25180 22100 25208
rect 21784 25168 21790 25180
rect 22088 25171 22100 25180
rect 22094 25168 22100 25171
rect 22152 25168 22158 25220
rect 22572 25208 22600 25236
rect 23845 25211 23903 25217
rect 23845 25208 23857 25211
rect 22572 25180 23857 25208
rect 23845 25177 23857 25180
rect 23891 25177 23903 25211
rect 23845 25171 23903 25177
rect 24213 25211 24271 25217
rect 24213 25177 24225 25211
rect 24259 25208 24271 25211
rect 25130 25208 25136 25220
rect 24259 25180 25136 25208
rect 24259 25177 24271 25180
rect 24213 25171 24271 25177
rect 25130 25168 25136 25180
rect 25188 25168 25194 25220
rect 12759 25112 18460 25140
rect 18509 25143 18567 25149
rect 12759 25109 12771 25112
rect 12713 25103 12771 25109
rect 18509 25109 18521 25143
rect 18555 25140 18567 25143
rect 19426 25140 19432 25152
rect 18555 25112 19432 25140
rect 18555 25109 18567 25112
rect 18509 25103 18567 25109
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 19702 25100 19708 25152
rect 19760 25140 19766 25152
rect 22554 25140 22560 25152
rect 19760 25112 22560 25140
rect 19760 25100 19766 25112
rect 22554 25100 22560 25112
rect 22612 25100 22618 25152
rect 23661 25143 23719 25149
rect 23661 25109 23673 25143
rect 23707 25140 23719 25143
rect 23750 25140 23756 25152
rect 23707 25112 23756 25140
rect 23707 25109 23719 25112
rect 23661 25103 23719 25109
rect 23750 25100 23756 25112
rect 23808 25100 23814 25152
rect 1104 25050 25000 25072
rect 1104 24998 6884 25050
rect 6936 24998 6948 25050
rect 7000 24998 7012 25050
rect 7064 24998 7076 25050
rect 7128 24998 7140 25050
rect 7192 24998 12818 25050
rect 12870 24998 12882 25050
rect 12934 24998 12946 25050
rect 12998 24998 13010 25050
rect 13062 24998 13074 25050
rect 13126 24998 18752 25050
rect 18804 24998 18816 25050
rect 18868 24998 18880 25050
rect 18932 24998 18944 25050
rect 18996 24998 19008 25050
rect 19060 24998 24686 25050
rect 24738 24998 24750 25050
rect 24802 24998 24814 25050
rect 24866 24998 24878 25050
rect 24930 24998 24942 25050
rect 24994 24998 25000 25050
rect 1104 24976 25000 24998
rect 1118 24896 1124 24948
rect 1176 24936 1182 24948
rect 1302 24936 1308 24948
rect 1176 24908 1308 24936
rect 1176 24896 1182 24908
rect 1302 24896 1308 24908
rect 1360 24896 1366 24948
rect 1578 24896 1584 24948
rect 1636 24896 1642 24948
rect 1946 24896 1952 24948
rect 2004 24936 2010 24948
rect 2004 24908 3648 24936
rect 2004 24896 2010 24908
rect 1026 24828 1032 24880
rect 1084 24868 1090 24880
rect 3620 24877 3648 24908
rect 3694 24896 3700 24948
rect 3752 24936 3758 24948
rect 3973 24939 4031 24945
rect 3973 24936 3985 24939
rect 3752 24908 3985 24936
rect 3752 24896 3758 24908
rect 3973 24905 3985 24908
rect 4019 24905 4031 24939
rect 3973 24899 4031 24905
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 4982 24936 4988 24948
rect 4764 24908 4988 24936
rect 4764 24896 4770 24908
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 5258 24896 5264 24948
rect 5316 24936 5322 24948
rect 5316 24908 17264 24936
rect 5316 24896 5322 24908
rect 2869 24871 2927 24877
rect 1084 24840 1808 24868
rect 1084 24828 1090 24840
rect 750 24760 756 24812
rect 808 24800 814 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 808 24772 1409 24800
rect 808 24760 814 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 1578 24760 1584 24812
rect 1636 24800 1642 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 1636 24772 1685 24800
rect 1636 24760 1642 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 1780 24800 1808 24840
rect 2869 24837 2881 24871
rect 2915 24837 2927 24871
rect 3605 24871 3663 24877
rect 2869 24831 2927 24837
rect 3160 24840 3372 24868
rect 1949 24803 2007 24809
rect 1949 24800 1961 24803
rect 1780 24772 1961 24800
rect 1673 24763 1731 24769
rect 1949 24769 1961 24772
rect 1995 24769 2007 24803
rect 1949 24763 2007 24769
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24769 2283 24803
rect 2884 24800 2912 24831
rect 3050 24800 3056 24812
rect 2884 24772 3056 24800
rect 2225 24763 2283 24769
rect 1118 24692 1124 24744
rect 1176 24732 1182 24744
rect 2240 24732 2268 24763
rect 3050 24760 3056 24772
rect 3108 24760 3114 24812
rect 3160 24809 3188 24840
rect 3145 24803 3203 24809
rect 3145 24769 3157 24803
rect 3191 24769 3203 24803
rect 3145 24763 3203 24769
rect 3234 24760 3240 24812
rect 3292 24760 3298 24812
rect 3344 24800 3372 24840
rect 3605 24837 3617 24871
rect 3651 24868 3663 24871
rect 3878 24868 3884 24880
rect 3651 24840 3884 24868
rect 3651 24837 3663 24840
rect 3605 24831 3663 24837
rect 3878 24828 3884 24840
rect 3936 24828 3942 24880
rect 6270 24828 6276 24880
rect 6328 24868 6334 24880
rect 6328 24840 8248 24868
rect 6328 24828 6334 24840
rect 3418 24800 3424 24812
rect 3344 24772 3424 24800
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 3896 24800 3924 24828
rect 4341 24803 4399 24809
rect 4341 24800 4353 24803
rect 3896 24772 4353 24800
rect 4341 24769 4353 24772
rect 4387 24769 4399 24803
rect 4341 24763 4399 24769
rect 6181 24803 6239 24809
rect 6181 24769 6193 24803
rect 6227 24800 6239 24803
rect 6914 24800 6920 24812
rect 6227 24772 6920 24800
rect 6227 24769 6239 24772
rect 6181 24763 6239 24769
rect 6914 24760 6920 24772
rect 6972 24760 6978 24812
rect 8220 24744 8248 24840
rect 8386 24828 8392 24880
rect 8444 24868 8450 24880
rect 17126 24868 17132 24880
rect 8444 24840 17132 24868
rect 8444 24828 8450 24840
rect 17126 24828 17132 24840
rect 17184 24828 17190 24880
rect 17236 24868 17264 24908
rect 17310 24896 17316 24948
rect 17368 24936 17374 24948
rect 17681 24939 17739 24945
rect 17681 24936 17693 24939
rect 17368 24908 17693 24936
rect 17368 24896 17374 24908
rect 17681 24905 17693 24908
rect 17727 24905 17739 24939
rect 19702 24936 19708 24948
rect 17681 24899 17739 24905
rect 17788 24908 19708 24936
rect 17788 24868 17816 24908
rect 19702 24896 19708 24908
rect 19760 24896 19766 24948
rect 19978 24896 19984 24948
rect 20036 24936 20042 24948
rect 20036 24908 21496 24936
rect 20036 24896 20042 24908
rect 17236 24840 17816 24868
rect 17954 24828 17960 24880
rect 18012 24868 18018 24880
rect 18012 24840 18164 24868
rect 18012 24828 18018 24840
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8755 24803 8813 24809
rect 8755 24800 8767 24803
rect 8720 24772 8767 24800
rect 8720 24760 8726 24772
rect 8755 24769 8767 24772
rect 8801 24769 8813 24803
rect 8755 24763 8813 24769
rect 8846 24760 8852 24812
rect 8904 24800 8910 24812
rect 11514 24800 11520 24812
rect 8904 24772 11520 24800
rect 8904 24760 8910 24772
rect 11514 24760 11520 24772
rect 11572 24760 11578 24812
rect 11606 24760 11612 24812
rect 11664 24800 11670 24812
rect 12435 24803 12493 24809
rect 12435 24800 12447 24803
rect 11664 24772 12447 24800
rect 11664 24760 11670 24772
rect 12435 24769 12447 24772
rect 12481 24800 12493 24803
rect 13630 24800 13636 24812
rect 12481 24772 13636 24800
rect 12481 24769 12493 24772
rect 12435 24763 12493 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 13906 24760 13912 24812
rect 13964 24800 13970 24812
rect 15470 24800 15476 24812
rect 13964 24772 15476 24800
rect 13964 24760 13970 24772
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 16943 24803 17001 24809
rect 16943 24769 16955 24803
rect 16989 24800 17001 24803
rect 17402 24800 17408 24812
rect 16989 24772 17408 24800
rect 16989 24769 17001 24772
rect 16943 24763 17001 24769
rect 17402 24760 17408 24772
rect 17460 24760 17466 24812
rect 17494 24760 17500 24812
rect 17552 24800 17558 24812
rect 18049 24803 18107 24809
rect 18049 24800 18061 24803
rect 17552 24772 18061 24800
rect 17552 24760 17558 24772
rect 18049 24769 18061 24772
rect 18095 24769 18107 24803
rect 18136 24800 18164 24840
rect 19426 24828 19432 24880
rect 19484 24868 19490 24880
rect 21468 24868 21496 24908
rect 21542 24896 21548 24948
rect 21600 24936 21606 24948
rect 21821 24939 21879 24945
rect 21821 24936 21833 24939
rect 21600 24908 21833 24936
rect 21600 24896 21606 24908
rect 21821 24905 21833 24908
rect 21867 24905 21879 24939
rect 21821 24899 21879 24905
rect 23474 24896 23480 24948
rect 23532 24896 23538 24948
rect 19484 24840 20116 24868
rect 21468 24840 22122 24868
rect 19484 24828 19490 24840
rect 18291 24803 18349 24809
rect 18291 24800 18303 24803
rect 18136 24772 18303 24800
rect 18049 24763 18107 24769
rect 18291 24769 18303 24772
rect 18337 24769 18349 24803
rect 20088 24800 20116 24840
rect 20162 24809 20168 24812
rect 20145 24803 20168 24809
rect 20145 24800 20157 24803
rect 20088 24772 20157 24800
rect 18291 24763 18349 24769
rect 20145 24769 20157 24772
rect 20145 24763 20168 24769
rect 20162 24760 20168 24763
rect 20220 24760 20226 24812
rect 21358 24760 21364 24812
rect 21416 24760 21422 24812
rect 22005 24803 22063 24809
rect 22005 24800 22017 24803
rect 21468 24772 22017 24800
rect 1176 24704 2268 24732
rect 1176 24692 1182 24704
rect 3510 24692 3516 24744
rect 3568 24692 3574 24744
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 4706 24732 4712 24744
rect 4571 24704 4712 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 4706 24692 4712 24704
rect 4764 24732 4770 24744
rect 5074 24732 5080 24744
rect 4764 24704 5080 24732
rect 4764 24692 4770 24704
rect 5074 24692 5080 24704
rect 5132 24692 5138 24744
rect 5258 24692 5264 24744
rect 5316 24692 5322 24744
rect 5442 24741 5448 24744
rect 5399 24735 5448 24741
rect 5399 24701 5411 24735
rect 5445 24701 5448 24735
rect 5399 24695 5448 24701
rect 5442 24692 5448 24695
rect 5500 24692 5506 24744
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24732 5595 24735
rect 6362 24732 6368 24744
rect 5583 24704 6368 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 6362 24692 6368 24704
rect 6420 24692 6426 24744
rect 8202 24692 8208 24744
rect 8260 24692 8266 24744
rect 8478 24692 8484 24744
rect 8536 24692 8542 24744
rect 11146 24692 11152 24744
rect 11204 24732 11210 24744
rect 12158 24732 12164 24744
rect 11204 24704 12164 24732
rect 11204 24692 11210 24704
rect 12158 24692 12164 24704
rect 12216 24692 12222 24744
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 16666 24732 16672 24744
rect 14332 24704 16672 24732
rect 14332 24692 14338 24704
rect 16666 24692 16672 24704
rect 16724 24692 16730 24744
rect 19889 24735 19947 24741
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 2133 24667 2191 24673
rect 2133 24633 2145 24667
rect 2179 24664 2191 24667
rect 2314 24664 2320 24676
rect 2179 24636 2320 24664
rect 2179 24633 2191 24636
rect 2133 24627 2191 24633
rect 2314 24624 2320 24636
rect 2372 24624 2378 24676
rect 4062 24624 4068 24676
rect 4120 24664 4126 24676
rect 4614 24664 4620 24676
rect 4120 24636 4620 24664
rect 4120 24624 4126 24636
rect 4614 24624 4620 24636
rect 4672 24624 4678 24676
rect 4985 24667 5043 24673
rect 4985 24633 4997 24667
rect 5031 24633 5043 24667
rect 4985 24627 5043 24633
rect 1762 24556 1768 24608
rect 1820 24596 1826 24608
rect 1857 24599 1915 24605
rect 1857 24596 1869 24599
rect 1820 24568 1869 24596
rect 1820 24556 1826 24568
rect 1857 24565 1869 24568
rect 1903 24565 1915 24599
rect 1857 24559 1915 24565
rect 2409 24599 2467 24605
rect 2409 24565 2421 24599
rect 2455 24596 2467 24599
rect 2774 24596 2780 24608
rect 2455 24568 2780 24596
rect 2455 24565 2467 24568
rect 2409 24559 2467 24565
rect 2774 24556 2780 24568
rect 2832 24556 2838 24608
rect 4157 24599 4215 24605
rect 4157 24565 4169 24599
rect 4203 24596 4215 24599
rect 4890 24596 4896 24608
rect 4203 24568 4896 24596
rect 4203 24565 4215 24568
rect 4157 24559 4215 24565
rect 4890 24556 4896 24568
rect 4948 24556 4954 24608
rect 5000 24596 5028 24627
rect 6546 24624 6552 24676
rect 6604 24664 6610 24676
rect 7926 24664 7932 24676
rect 6604 24636 7932 24664
rect 6604 24624 6610 24636
rect 7926 24624 7932 24636
rect 7984 24624 7990 24676
rect 9493 24667 9551 24673
rect 9493 24633 9505 24667
rect 9539 24664 9551 24667
rect 9674 24664 9680 24676
rect 9539 24636 9680 24664
rect 9539 24633 9551 24636
rect 9493 24627 9551 24633
rect 9674 24624 9680 24636
rect 9732 24624 9738 24676
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 11882 24664 11888 24676
rect 10376 24636 11888 24664
rect 10376 24624 10382 24636
rect 11882 24624 11888 24636
rect 11940 24624 11946 24676
rect 13096 24636 14504 24664
rect 5718 24596 5724 24608
rect 5000 24568 5724 24596
rect 5718 24556 5724 24568
rect 5776 24556 5782 24608
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 13096 24596 13124 24636
rect 14476 24608 14504 24636
rect 17862 24624 17868 24676
rect 17920 24624 17926 24676
rect 6328 24568 13124 24596
rect 6328 24556 6334 24568
rect 13170 24556 13176 24608
rect 13228 24556 13234 24608
rect 14458 24556 14464 24608
rect 14516 24556 14522 24608
rect 15378 24556 15384 24608
rect 15436 24596 15442 24608
rect 16114 24596 16120 24608
rect 15436 24568 16120 24596
rect 15436 24556 15442 24568
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 16574 24556 16580 24608
rect 16632 24596 16638 24608
rect 17770 24596 17776 24608
rect 16632 24568 17776 24596
rect 16632 24556 16638 24568
rect 17770 24556 17776 24568
rect 17828 24556 17834 24608
rect 17880 24596 17908 24624
rect 19061 24599 19119 24605
rect 19061 24596 19073 24599
rect 17880 24568 19073 24596
rect 19061 24565 19073 24568
rect 19107 24565 19119 24599
rect 19904 24596 19932 24695
rect 21269 24667 21327 24673
rect 21269 24633 21281 24667
rect 21315 24664 21327 24667
rect 21468 24664 21496 24772
rect 22005 24769 22017 24772
rect 22051 24769 22063 24803
rect 22005 24763 22063 24769
rect 21542 24692 21548 24744
rect 21600 24732 21606 24744
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21600 24704 21649 24732
rect 21600 24692 21606 24704
rect 21637 24701 21649 24704
rect 21683 24701 21695 24735
rect 22094 24732 22122 24840
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 22707 24803 22765 24809
rect 22707 24800 22719 24803
rect 22428 24772 22719 24800
rect 22428 24760 22434 24772
rect 22707 24769 22719 24772
rect 22753 24769 22765 24803
rect 22707 24763 22765 24769
rect 24121 24803 24179 24809
rect 24121 24769 24133 24803
rect 24167 24800 24179 24803
rect 24210 24800 24216 24812
rect 24167 24772 24216 24800
rect 24167 24769 24179 24772
rect 24121 24763 24179 24769
rect 24210 24760 24216 24772
rect 24268 24760 24274 24812
rect 22186 24732 22192 24744
rect 22094 24704 22192 24732
rect 21637 24695 21695 24701
rect 22186 24692 22192 24704
rect 22244 24732 22250 24744
rect 22465 24735 22523 24741
rect 22465 24732 22477 24735
rect 22244 24704 22477 24732
rect 22244 24692 22250 24704
rect 22465 24701 22477 24704
rect 22511 24701 22523 24735
rect 22465 24695 22523 24701
rect 21315 24636 21496 24664
rect 21560 24636 22094 24664
rect 21315 24633 21327 24636
rect 21269 24627 21327 24633
rect 20622 24596 20628 24608
rect 19904 24568 20628 24596
rect 19061 24559 19119 24565
rect 20622 24556 20628 24568
rect 20680 24596 20686 24608
rect 21174 24596 21180 24608
rect 20680 24568 21180 24596
rect 20680 24556 20686 24568
rect 21174 24556 21180 24568
rect 21232 24556 21238 24608
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 21560 24605 21588 24636
rect 21545 24599 21603 24605
rect 21545 24565 21557 24599
rect 21591 24565 21603 24599
rect 22066 24596 22094 24636
rect 24302 24624 24308 24676
rect 24360 24624 24366 24676
rect 24320 24596 24348 24624
rect 22066 24568 24348 24596
rect 21545 24559 21603 24565
rect 24394 24556 24400 24608
rect 24452 24556 24458 24608
rect 1104 24506 24840 24528
rect 1104 24454 3917 24506
rect 3969 24454 3981 24506
rect 4033 24454 4045 24506
rect 4097 24454 4109 24506
rect 4161 24454 4173 24506
rect 4225 24454 9851 24506
rect 9903 24454 9915 24506
rect 9967 24454 9979 24506
rect 10031 24454 10043 24506
rect 10095 24454 10107 24506
rect 10159 24454 15785 24506
rect 15837 24454 15849 24506
rect 15901 24454 15913 24506
rect 15965 24454 15977 24506
rect 16029 24454 16041 24506
rect 16093 24454 21719 24506
rect 21771 24454 21783 24506
rect 21835 24454 21847 24506
rect 21899 24454 21911 24506
rect 21963 24454 21975 24506
rect 22027 24454 24840 24506
rect 1104 24432 24840 24454
rect 2774 24352 2780 24404
rect 2832 24352 2838 24404
rect 2866 24352 2872 24404
rect 2924 24352 2930 24404
rect 3050 24352 3056 24404
rect 3108 24352 3114 24404
rect 6914 24352 6920 24404
rect 6972 24352 6978 24404
rect 7009 24395 7067 24401
rect 7009 24361 7021 24395
rect 7055 24392 7067 24395
rect 9030 24392 9036 24404
rect 7055 24364 7604 24392
rect 7055 24361 7067 24364
rect 7009 24355 7067 24361
rect 2406 24216 2412 24268
rect 2464 24216 2470 24268
rect 2792 24256 2820 24352
rect 3068 24324 3096 24352
rect 5442 24324 5448 24336
rect 3068 24296 5448 24324
rect 5442 24284 5448 24296
rect 5500 24284 5506 24336
rect 5810 24284 5816 24336
rect 5868 24284 5874 24336
rect 4154 24256 4160 24268
rect 2792 24228 4160 24256
rect 4154 24216 4160 24228
rect 4212 24216 4218 24268
rect 4522 24216 4528 24268
rect 4580 24256 4586 24268
rect 4798 24256 4804 24268
rect 4580 24228 4804 24256
rect 4580 24216 4586 24228
rect 4798 24216 4804 24228
rect 4856 24256 4862 24268
rect 5169 24259 5227 24265
rect 5169 24256 5181 24259
rect 4856 24228 5181 24256
rect 4856 24216 4862 24228
rect 5169 24225 5181 24228
rect 5215 24225 5227 24259
rect 5169 24219 5227 24225
rect 5258 24216 5264 24268
rect 5316 24256 5322 24268
rect 6206 24259 6264 24265
rect 6206 24256 6218 24259
rect 5316 24228 6218 24256
rect 5316 24216 5322 24228
rect 6206 24225 6218 24228
rect 6252 24225 6264 24259
rect 6206 24219 6264 24225
rect 6362 24216 6368 24268
rect 6420 24216 6426 24268
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24188 2007 24191
rect 2498 24188 2504 24200
rect 1995 24160 2504 24188
rect 1995 24157 2007 24160
rect 1949 24151 2007 24157
rect 2498 24148 2504 24160
rect 2556 24148 2562 24200
rect 2700 24160 3372 24188
rect 1486 24080 1492 24132
rect 1544 24120 1550 24132
rect 1581 24123 1639 24129
rect 1581 24120 1593 24123
rect 1544 24092 1593 24120
rect 1544 24080 1550 24092
rect 1581 24089 1593 24092
rect 1627 24089 1639 24123
rect 1581 24083 1639 24089
rect 1854 24080 1860 24132
rect 1912 24080 1918 24132
rect 2700 24129 2728 24160
rect 2317 24123 2375 24129
rect 2317 24089 2329 24123
rect 2363 24089 2375 24123
rect 2317 24083 2375 24089
rect 2685 24123 2743 24129
rect 2685 24089 2697 24123
rect 2731 24089 2743 24123
rect 3344 24120 3372 24160
rect 3418 24148 3424 24200
rect 3476 24188 3482 24200
rect 3694 24188 3700 24200
rect 3476 24160 3700 24188
rect 3476 24148 3482 24160
rect 3694 24148 3700 24160
rect 3752 24188 3758 24200
rect 4982 24188 4988 24200
rect 3752 24160 4988 24188
rect 3752 24148 3758 24160
rect 4982 24148 4988 24160
rect 5040 24188 5046 24200
rect 5353 24191 5411 24197
rect 5353 24188 5365 24191
rect 5040 24160 5365 24188
rect 5040 24148 5046 24160
rect 5353 24157 5365 24160
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 6086 24148 6092 24200
rect 6144 24148 6150 24200
rect 6932 24188 6960 24352
rect 7101 24327 7159 24333
rect 7101 24293 7113 24327
rect 7147 24324 7159 24327
rect 7147 24296 7512 24324
rect 7147 24293 7159 24296
rect 7101 24287 7159 24293
rect 7484 24197 7512 24296
rect 7285 24191 7343 24197
rect 7285 24188 7297 24191
rect 6932 24160 7297 24188
rect 7285 24157 7297 24160
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24157 7527 24191
rect 7576 24188 7604 24364
rect 8404 24364 9036 24392
rect 8404 24336 8432 24364
rect 9030 24352 9036 24364
rect 9088 24392 9094 24404
rect 10318 24392 10324 24404
rect 9088 24364 10324 24392
rect 9088 24352 9094 24364
rect 10318 24352 10324 24364
rect 10376 24352 10382 24404
rect 10962 24392 10968 24404
rect 10612 24364 10968 24392
rect 8386 24284 8392 24336
rect 8444 24284 8450 24336
rect 9766 24216 9772 24268
rect 9824 24256 9830 24268
rect 10226 24256 10232 24268
rect 9824 24228 10232 24256
rect 9824 24216 9830 24228
rect 10226 24216 10232 24228
rect 10284 24216 10290 24268
rect 10612 24265 10640 24364
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 11514 24352 11520 24404
rect 11572 24392 11578 24404
rect 16574 24392 16580 24404
rect 11572 24364 16580 24392
rect 11572 24352 11578 24364
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 17957 24395 18015 24401
rect 17957 24392 17969 24395
rect 16868 24364 17969 24392
rect 14090 24284 14096 24336
rect 14148 24324 14154 24336
rect 16868 24324 16896 24364
rect 17957 24361 17969 24364
rect 18003 24361 18015 24395
rect 17957 24355 18015 24361
rect 19521 24395 19579 24401
rect 19521 24361 19533 24395
rect 19567 24392 19579 24395
rect 20993 24395 21051 24401
rect 19567 24364 20024 24392
rect 19567 24361 19579 24364
rect 19521 24355 19579 24361
rect 14148 24296 15792 24324
rect 14148 24284 14154 24296
rect 10597 24259 10655 24265
rect 10597 24225 10609 24259
rect 10643 24225 10655 24259
rect 10597 24219 10655 24225
rect 12158 24216 12164 24268
rect 12216 24256 12222 24268
rect 12621 24259 12679 24265
rect 12621 24256 12633 24259
rect 12216 24228 12633 24256
rect 12216 24216 12222 24228
rect 12621 24225 12633 24228
rect 12667 24225 12679 24259
rect 12621 24219 12679 24225
rect 13538 24216 13544 24268
rect 13596 24256 13602 24268
rect 14918 24256 14924 24268
rect 13596 24228 14924 24256
rect 13596 24216 13602 24228
rect 14918 24216 14924 24228
rect 14976 24216 14982 24268
rect 15013 24259 15071 24265
rect 15013 24225 15025 24259
rect 15059 24256 15071 24259
rect 15102 24256 15108 24268
rect 15059 24228 15108 24256
rect 15059 24225 15071 24228
rect 15013 24219 15071 24225
rect 15102 24216 15108 24228
rect 15160 24216 15166 24268
rect 15197 24259 15255 24265
rect 15197 24225 15209 24259
rect 15243 24256 15255 24259
rect 15286 24256 15292 24268
rect 15243 24228 15292 24256
rect 15243 24225 15255 24228
rect 15197 24219 15255 24225
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 15654 24216 15660 24268
rect 15712 24216 15718 24268
rect 15764 24256 15792 24296
rect 16684 24296 16896 24324
rect 16209 24259 16267 24265
rect 15764 24228 16068 24256
rect 16040 24200 16068 24228
rect 16209 24225 16221 24259
rect 16255 24256 16267 24259
rect 16684 24256 16712 24296
rect 16255 24228 16712 24256
rect 16255 24225 16267 24228
rect 16209 24219 16267 24225
rect 16758 24216 16764 24268
rect 16816 24256 16822 24268
rect 16945 24259 17003 24265
rect 16945 24256 16957 24259
rect 16816 24228 16957 24256
rect 16816 24216 16822 24228
rect 16945 24225 16957 24228
rect 16991 24225 17003 24259
rect 16945 24219 17003 24225
rect 17604 24228 19932 24256
rect 7929 24191 7987 24197
rect 7929 24188 7941 24191
rect 7576 24160 7941 24188
rect 7469 24151 7527 24157
rect 7929 24157 7941 24160
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 8294 24148 8300 24200
rect 8352 24188 8358 24200
rect 8941 24191 8999 24197
rect 8941 24188 8953 24191
rect 8352 24160 8953 24188
rect 8352 24148 8358 24160
rect 8941 24157 8953 24160
rect 8987 24157 8999 24191
rect 8941 24151 8999 24157
rect 9215 24191 9273 24197
rect 9215 24157 9227 24191
rect 9261 24188 9273 24191
rect 9582 24188 9588 24200
rect 9261 24160 9588 24188
rect 9261 24157 9273 24160
rect 9215 24151 9273 24157
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 10870 24188 10876 24200
rect 10831 24160 10876 24188
rect 10870 24148 10876 24160
rect 10928 24148 10934 24200
rect 11882 24148 11888 24200
rect 11940 24188 11946 24200
rect 12895 24191 12953 24197
rect 12895 24188 12907 24191
rect 11940 24160 12907 24188
rect 11940 24148 11946 24160
rect 12895 24157 12907 24160
rect 12941 24188 12953 24191
rect 12941 24160 14596 24188
rect 12941 24157 12953 24160
rect 12895 24151 12953 24157
rect 4430 24120 4436 24132
rect 3344 24092 4436 24120
rect 2685 24083 2743 24089
rect 2332 24052 2360 24083
rect 4430 24080 4436 24092
rect 4488 24080 4494 24132
rect 4614 24080 4620 24132
rect 4672 24120 4678 24132
rect 5258 24120 5264 24132
rect 4672 24092 5264 24120
rect 4672 24080 4678 24092
rect 5258 24080 5264 24092
rect 5316 24080 5322 24132
rect 10318 24120 10324 24132
rect 6838 24092 10324 24120
rect 2590 24052 2596 24064
rect 2332 24024 2596 24052
rect 2590 24012 2596 24024
rect 2648 24012 2654 24064
rect 4154 24012 4160 24064
rect 4212 24052 4218 24064
rect 6838 24052 6866 24092
rect 10318 24080 10324 24092
rect 10376 24080 10382 24132
rect 12250 24080 12256 24132
rect 12308 24120 12314 24132
rect 14458 24120 14464 24132
rect 12308 24092 14464 24120
rect 12308 24080 12314 24092
rect 14458 24080 14464 24092
rect 14516 24080 14522 24132
rect 14568 24064 14596 24160
rect 15930 24148 15936 24200
rect 15988 24148 15994 24200
rect 16022 24148 16028 24200
rect 16080 24197 16086 24200
rect 16080 24191 16108 24197
rect 16096 24157 16108 24191
rect 17187 24191 17245 24197
rect 17187 24188 17199 24191
rect 16080 24151 16108 24157
rect 17052 24160 17199 24188
rect 16080 24148 16086 24151
rect 17052 24120 17080 24160
rect 17187 24157 17199 24160
rect 17233 24157 17245 24191
rect 17187 24151 17245 24157
rect 16684 24092 17080 24120
rect 4212 24024 6866 24052
rect 4212 24012 4218 24024
rect 7558 24012 7564 24064
rect 7616 24012 7622 24064
rect 7742 24012 7748 24064
rect 7800 24012 7806 24064
rect 9674 24012 9680 24064
rect 9732 24052 9738 24064
rect 9953 24055 10011 24061
rect 9953 24052 9965 24055
rect 9732 24024 9965 24052
rect 9732 24012 9738 24024
rect 9953 24021 9965 24024
rect 9999 24021 10011 24055
rect 9953 24015 10011 24021
rect 11238 24012 11244 24064
rect 11296 24052 11302 24064
rect 11609 24055 11667 24061
rect 11609 24052 11621 24055
rect 11296 24024 11621 24052
rect 11296 24012 11302 24024
rect 11609 24021 11621 24024
rect 11655 24021 11667 24055
rect 11609 24015 11667 24021
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 13814 24052 13820 24064
rect 13679 24024 13820 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14550 24012 14556 24064
rect 14608 24012 14614 24064
rect 14918 24012 14924 24064
rect 14976 24052 14982 24064
rect 16684 24052 16712 24092
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 17604 24120 17632 24228
rect 19242 24148 19248 24200
rect 19300 24188 19306 24200
rect 19705 24191 19763 24197
rect 19705 24188 19717 24191
rect 19300 24160 19717 24188
rect 19300 24148 19306 24160
rect 19705 24157 19717 24160
rect 19751 24157 19763 24191
rect 19705 24151 19763 24157
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 17552 24092 17632 24120
rect 17552 24080 17558 24092
rect 14976 24024 16712 24052
rect 16853 24055 16911 24061
rect 14976 24012 14982 24024
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 17402 24052 17408 24064
rect 16899 24024 17408 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 17402 24012 17408 24024
rect 17460 24012 17466 24064
rect 19610 24012 19616 24064
rect 19668 24052 19674 24064
rect 19812 24052 19840 24151
rect 19904 24120 19932 24228
rect 19996 24197 20024 24364
rect 20993 24361 21005 24395
rect 21039 24392 21051 24395
rect 21450 24392 21456 24404
rect 21039 24364 21456 24392
rect 21039 24361 21051 24364
rect 20993 24355 21051 24361
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 22370 24392 22376 24404
rect 22066 24364 22376 24392
rect 22066 24324 22094 24364
rect 22370 24352 22376 24364
rect 22428 24352 22434 24404
rect 22646 24352 22652 24404
rect 22704 24352 22710 24404
rect 23382 24352 23388 24404
rect 23440 24352 23446 24404
rect 20088 24296 22094 24324
rect 22664 24324 22692 24352
rect 23845 24327 23903 24333
rect 23845 24324 23857 24327
rect 22664 24296 23857 24324
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24157 20039 24191
rect 19981 24151 20039 24157
rect 20088 24120 20116 24296
rect 23845 24293 23857 24296
rect 23891 24293 23903 24327
rect 23845 24287 23903 24293
rect 21082 24216 21088 24268
rect 21140 24256 21146 24268
rect 21140 24228 23980 24256
rect 21140 24216 21146 24228
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20533 24191 20591 24197
rect 20533 24188 20545 24191
rect 20220 24160 20545 24188
rect 20220 24148 20226 24160
rect 20533 24157 20545 24160
rect 20579 24157 20591 24191
rect 20533 24151 20591 24157
rect 20901 24191 20959 24197
rect 20901 24157 20913 24191
rect 20947 24157 20959 24191
rect 20901 24151 20959 24157
rect 20916 24120 20944 24151
rect 22462 24148 22468 24200
rect 22520 24188 22526 24200
rect 23290 24188 23296 24200
rect 22520 24160 23296 24188
rect 22520 24148 22526 24160
rect 23290 24148 23296 24160
rect 23348 24148 23354 24200
rect 23566 24148 23572 24200
rect 23624 24148 23630 24200
rect 23658 24148 23664 24200
rect 23716 24148 23722 24200
rect 23952 24197 23980 24228
rect 23937 24191 23995 24197
rect 23937 24157 23949 24191
rect 23983 24157 23995 24191
rect 23937 24151 23995 24157
rect 19904 24092 20116 24120
rect 20364 24092 20944 24120
rect 19668 24024 19840 24052
rect 19668 24012 19674 24024
rect 19886 24012 19892 24064
rect 19944 24012 19950 24064
rect 20364 24061 20392 24092
rect 20349 24055 20407 24061
rect 20349 24021 20361 24055
rect 20395 24021 20407 24055
rect 20349 24015 20407 24021
rect 20898 24012 20904 24064
rect 20956 24052 20962 24064
rect 21174 24052 21180 24064
rect 20956 24024 21180 24052
rect 20956 24012 20962 24024
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 24121 24055 24179 24061
rect 24121 24021 24133 24055
rect 24167 24052 24179 24055
rect 25130 24052 25136 24064
rect 24167 24024 25136 24052
rect 24167 24021 24179 24024
rect 24121 24015 24179 24021
rect 25130 24012 25136 24024
rect 25188 24012 25194 24064
rect 1104 23962 25000 23984
rect 1104 23910 6884 23962
rect 6936 23910 6948 23962
rect 7000 23910 7012 23962
rect 7064 23910 7076 23962
rect 7128 23910 7140 23962
rect 7192 23910 12818 23962
rect 12870 23910 12882 23962
rect 12934 23910 12946 23962
rect 12998 23910 13010 23962
rect 13062 23910 13074 23962
rect 13126 23910 18752 23962
rect 18804 23910 18816 23962
rect 18868 23910 18880 23962
rect 18932 23910 18944 23962
rect 18996 23910 19008 23962
rect 19060 23910 24686 23962
rect 24738 23910 24750 23962
rect 24802 23910 24814 23962
rect 24866 23910 24878 23962
rect 24930 23910 24942 23962
rect 24994 23910 25000 23962
rect 1104 23888 25000 23910
rect 1854 23808 1860 23860
rect 1912 23848 1918 23860
rect 1912 23820 3464 23848
rect 1912 23808 1918 23820
rect 3436 23780 3464 23820
rect 3510 23808 3516 23860
rect 3568 23808 3574 23860
rect 4062 23808 4068 23860
rect 4120 23808 4126 23860
rect 4890 23808 4896 23860
rect 4948 23848 4954 23860
rect 9766 23848 9772 23860
rect 4948 23820 9772 23848
rect 4948 23808 4954 23820
rect 9766 23808 9772 23820
rect 9824 23808 9830 23860
rect 9858 23808 9864 23860
rect 9916 23848 9922 23860
rect 9953 23851 10011 23857
rect 9953 23848 9965 23851
rect 9916 23820 9965 23848
rect 9916 23808 9922 23820
rect 9953 23817 9965 23820
rect 9999 23817 10011 23851
rect 9953 23811 10011 23817
rect 10318 23808 10324 23860
rect 10376 23848 10382 23860
rect 13354 23848 13360 23860
rect 10376 23820 13360 23848
rect 10376 23808 10382 23820
rect 3602 23780 3608 23792
rect 3436 23752 3608 23780
rect 3602 23740 3608 23752
rect 3660 23780 3666 23792
rect 6086 23780 6092 23792
rect 3660 23752 6092 23780
rect 3660 23740 3666 23752
rect 6086 23740 6092 23752
rect 6144 23780 6150 23792
rect 6362 23780 6368 23792
rect 6144 23752 6368 23780
rect 6144 23740 6150 23752
rect 6362 23740 6368 23752
rect 6420 23740 6426 23792
rect 7282 23780 7288 23792
rect 6932 23752 7288 23780
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 3881 23715 3939 23721
rect 3881 23712 3893 23715
rect 2832 23684 2875 23712
rect 3528 23684 3893 23712
rect 2832 23672 2838 23684
rect 1394 23604 1400 23656
rect 1452 23604 1458 23656
rect 1673 23647 1731 23653
rect 1673 23613 1685 23647
rect 1719 23613 1731 23647
rect 1673 23607 1731 23613
rect 1688 23508 1716 23607
rect 2222 23604 2228 23656
rect 2280 23644 2286 23656
rect 2501 23647 2559 23653
rect 2501 23644 2513 23647
rect 2280 23616 2513 23644
rect 2280 23604 2286 23616
rect 2501 23613 2513 23616
rect 2547 23613 2559 23647
rect 2501 23607 2559 23613
rect 3528 23588 3556 23684
rect 3881 23681 3893 23684
rect 3927 23712 3939 23715
rect 5442 23712 5448 23724
rect 3927 23684 5448 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 5442 23672 5448 23684
rect 5500 23672 5506 23724
rect 6932 23721 6960 23752
rect 7282 23740 7288 23752
rect 7340 23740 7346 23792
rect 7742 23740 7748 23792
rect 7800 23780 7806 23792
rect 7800 23752 8524 23780
rect 7800 23740 7806 23752
rect 6917 23715 6975 23721
rect 6917 23681 6929 23715
rect 6963 23681 6975 23715
rect 6917 23675 6975 23681
rect 7191 23715 7249 23721
rect 7191 23681 7203 23715
rect 7237 23712 7249 23715
rect 7237 23684 7880 23712
rect 7237 23681 7249 23684
rect 7191 23675 7249 23681
rect 7852 23644 7880 23684
rect 8110 23672 8116 23724
rect 8168 23712 8174 23724
rect 8496 23721 8524 23752
rect 8846 23740 8852 23792
rect 8904 23740 8910 23792
rect 9125 23783 9183 23789
rect 9125 23749 9137 23783
rect 9171 23749 9183 23783
rect 9125 23743 9183 23749
rect 8297 23715 8355 23721
rect 8297 23712 8309 23715
rect 8168 23684 8309 23712
rect 8168 23672 8174 23684
rect 8297 23681 8309 23684
rect 8343 23681 8355 23715
rect 8297 23675 8355 23681
rect 8481 23715 8539 23721
rect 8481 23681 8493 23715
rect 8527 23681 8539 23715
rect 9140 23712 9168 23743
rect 9214 23740 9220 23792
rect 9272 23740 9278 23792
rect 10134 23780 10140 23792
rect 9416 23752 10140 23780
rect 9416 23712 9444 23752
rect 10134 23740 10140 23752
rect 10192 23780 10198 23792
rect 11790 23780 11796 23792
rect 10192 23752 11796 23780
rect 10192 23740 10198 23752
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 12250 23740 12256 23792
rect 12308 23740 12314 23792
rect 9582 23712 9588 23724
rect 9640 23722 9646 23724
rect 9766 23722 9772 23724
rect 9140 23684 9444 23712
rect 9543 23684 9588 23712
rect 8481 23675 8539 23681
rect 9582 23672 9588 23684
rect 9640 23694 9772 23722
rect 9640 23684 9674 23694
rect 9640 23672 9646 23684
rect 9766 23672 9772 23694
rect 9824 23672 9830 23724
rect 11606 23672 11612 23724
rect 11664 23712 11670 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11664 23684 11897 23712
rect 11664 23672 11670 23684
rect 11885 23681 11897 23684
rect 11931 23712 11943 23715
rect 12268 23712 12296 23740
rect 11931 23684 12296 23712
rect 12621 23715 12679 23721
rect 11931 23681 11943 23684
rect 11885 23675 11943 23681
rect 12621 23681 12633 23715
rect 12667 23712 12679 23715
rect 12818 23712 12846 23820
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 15654 23808 15660 23860
rect 15712 23808 15718 23860
rect 15930 23808 15936 23860
rect 15988 23808 15994 23860
rect 19242 23808 19248 23860
rect 19300 23808 19306 23860
rect 19702 23848 19708 23860
rect 19536 23820 19708 23848
rect 13722 23721 13728 23724
rect 12667 23684 12846 23712
rect 13679 23715 13728 23721
rect 12667 23681 12679 23684
rect 12621 23675 12679 23681
rect 13679 23681 13691 23715
rect 13725 23681 13728 23715
rect 13679 23675 13728 23681
rect 13722 23672 13728 23675
rect 13780 23672 13786 23724
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 14458 23672 14464 23724
rect 14516 23712 14522 23724
rect 14887 23715 14945 23721
rect 14887 23712 14899 23715
rect 14516 23684 14899 23712
rect 14516 23672 14522 23684
rect 14887 23681 14899 23684
rect 14933 23681 14945 23715
rect 15948 23712 15976 23808
rect 16574 23740 16580 23792
rect 16632 23780 16638 23792
rect 19536 23780 19564 23820
rect 19702 23808 19708 23820
rect 19760 23808 19766 23860
rect 22554 23808 22560 23860
rect 22612 23808 22618 23860
rect 22833 23851 22891 23857
rect 22833 23817 22845 23851
rect 22879 23817 22891 23851
rect 22833 23811 22891 23817
rect 19978 23780 19984 23792
rect 16632 23752 19564 23780
rect 19700 23752 19984 23780
rect 16632 23740 16638 23752
rect 19700 23742 19728 23752
rect 19628 23731 19728 23742
rect 19978 23740 19984 23752
rect 20036 23740 20042 23792
rect 19611 23725 19728 23731
rect 16209 23715 16267 23721
rect 16209 23712 16221 23715
rect 15948 23684 16221 23712
rect 14887 23675 14945 23681
rect 16209 23681 16221 23684
rect 16255 23681 16267 23715
rect 16209 23675 16267 23681
rect 17678 23672 17684 23724
rect 17736 23712 17742 23724
rect 17865 23715 17923 23721
rect 17865 23712 17877 23715
rect 17736 23684 17877 23712
rect 17736 23672 17742 23684
rect 17865 23681 17877 23684
rect 17911 23681 17923 23715
rect 18121 23715 18179 23721
rect 18121 23712 18133 23715
rect 17865 23675 17923 23681
rect 17972 23684 18133 23712
rect 8386 23644 8392 23656
rect 7852 23616 8392 23644
rect 8386 23604 8392 23616
rect 8444 23604 8450 23656
rect 9674 23604 9680 23656
rect 9732 23604 9738 23656
rect 11974 23604 11980 23656
rect 12032 23644 12038 23656
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12032 23616 12817 23644
rect 12032 23604 12038 23616
rect 12636 23588 12664 23616
rect 12805 23613 12817 23616
rect 12851 23613 12863 23647
rect 12805 23607 12863 23613
rect 13170 23604 13176 23656
rect 13228 23644 13234 23656
rect 13265 23647 13323 23653
rect 13265 23644 13277 23647
rect 13228 23616 13277 23644
rect 13228 23604 13234 23616
rect 13265 23613 13277 23616
rect 13311 23613 13323 23647
rect 13265 23607 13323 23613
rect 13354 23604 13360 23656
rect 13412 23644 13418 23656
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 13412 23616 13553 23644
rect 13412 23604 13418 23616
rect 13541 23613 13553 23616
rect 13587 23613 13599 23647
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 13541 23607 13599 23613
rect 14384 23616 14657 23644
rect 3510 23536 3516 23588
rect 3568 23536 3574 23588
rect 10134 23536 10140 23588
rect 10192 23536 10198 23588
rect 12618 23536 12624 23588
rect 12676 23536 12682 23588
rect 6546 23508 6552 23520
rect 1688 23480 6552 23508
rect 6546 23468 6552 23480
rect 6604 23468 6610 23520
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 8110 23508 8116 23520
rect 7984 23480 8116 23508
rect 7984 23468 7990 23480
rect 8110 23468 8116 23480
rect 8168 23468 8174 23520
rect 8386 23468 8392 23520
rect 8444 23468 8450 23520
rect 11514 23468 11520 23520
rect 11572 23508 11578 23520
rect 12069 23511 12127 23517
rect 12069 23508 12081 23511
rect 11572 23480 12081 23508
rect 11572 23468 11578 23480
rect 12069 23477 12081 23480
rect 12115 23477 12127 23511
rect 12069 23471 12127 23477
rect 13814 23468 13820 23520
rect 13872 23508 13878 23520
rect 14274 23508 14280 23520
rect 13872 23480 14280 23508
rect 13872 23468 13878 23480
rect 14274 23468 14280 23480
rect 14332 23508 14338 23520
rect 14384 23508 14412 23616
rect 14645 23613 14657 23616
rect 14691 23613 14703 23647
rect 17972 23644 18000 23684
rect 18121 23681 18133 23684
rect 18167 23712 18179 23715
rect 18414 23712 18420 23724
rect 18167 23684 18420 23712
rect 18167 23681 18179 23684
rect 18121 23675 18179 23681
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 19611 23691 19623 23725
rect 19657 23714 19728 23725
rect 19657 23691 19669 23714
rect 19611 23685 19669 23691
rect 22572 23712 22600 23808
rect 22848 23780 22876 23811
rect 23290 23808 23296 23860
rect 23348 23848 23354 23860
rect 23348 23820 24164 23848
rect 23348 23808 23354 23820
rect 24136 23789 24164 23820
rect 24121 23783 24179 23789
rect 22848 23752 23520 23780
rect 22646 23712 22652 23724
rect 22572 23684 22652 23712
rect 22646 23672 22652 23684
rect 22704 23712 22710 23724
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22704 23684 23029 23712
rect 22704 23672 22710 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23492 23721 23520 23752
rect 24121 23749 24133 23783
rect 24167 23749 24179 23783
rect 24121 23743 24179 23749
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23681 23443 23715
rect 23385 23675 23443 23681
rect 23477 23715 23535 23721
rect 23477 23681 23489 23715
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 14645 23607 14703 23613
rect 17880 23616 18000 23644
rect 19337 23647 19395 23653
rect 16022 23536 16028 23588
rect 16080 23576 16086 23588
rect 16206 23576 16212 23588
rect 16080 23548 16212 23576
rect 16080 23536 16086 23548
rect 16206 23536 16212 23548
rect 16264 23536 16270 23588
rect 14332 23480 14412 23508
rect 14461 23511 14519 23517
rect 14332 23468 14338 23480
rect 14461 23477 14473 23511
rect 14507 23508 14519 23511
rect 17880 23508 17908 23616
rect 19337 23613 19349 23647
rect 19383 23613 19395 23647
rect 23400 23644 23428 23675
rect 23934 23672 23940 23724
rect 23992 23672 23998 23724
rect 23400 23616 23796 23644
rect 19337 23607 19395 23613
rect 19352 23576 19380 23607
rect 23768 23585 23796 23616
rect 23753 23579 23811 23585
rect 19352 23548 19472 23576
rect 19444 23520 19472 23548
rect 23753 23545 23765 23579
rect 23799 23545 23811 23579
rect 23753 23539 23811 23545
rect 14507 23480 17908 23508
rect 14507 23477 14519 23480
rect 14461 23471 14519 23477
rect 19426 23468 19432 23520
rect 19484 23468 19490 23520
rect 19610 23468 19616 23520
rect 19668 23508 19674 23520
rect 20349 23511 20407 23517
rect 20349 23508 20361 23511
rect 19668 23480 20361 23508
rect 19668 23468 19674 23480
rect 20349 23477 20361 23480
rect 20395 23477 20407 23511
rect 20349 23471 20407 23477
rect 23290 23468 23296 23520
rect 23348 23468 23354 23520
rect 23566 23468 23572 23520
rect 23624 23468 23630 23520
rect 24394 23468 24400 23520
rect 24452 23468 24458 23520
rect 566 23400 572 23452
rect 624 23400 630 23452
rect 1104 23418 24840 23440
rect 584 23248 612 23400
rect 1104 23366 3917 23418
rect 3969 23366 3981 23418
rect 4033 23366 4045 23418
rect 4097 23366 4109 23418
rect 4161 23366 4173 23418
rect 4225 23366 9851 23418
rect 9903 23366 9915 23418
rect 9967 23366 9979 23418
rect 10031 23366 10043 23418
rect 10095 23366 10107 23418
rect 10159 23366 15785 23418
rect 15837 23366 15849 23418
rect 15901 23366 15913 23418
rect 15965 23366 15977 23418
rect 16029 23366 16041 23418
rect 16093 23366 21719 23418
rect 21771 23366 21783 23418
rect 21835 23366 21847 23418
rect 21899 23366 21911 23418
rect 21963 23366 21975 23418
rect 22027 23366 24840 23418
rect 1104 23344 24840 23366
rect 676 23276 2360 23304
rect 676 23248 704 23276
rect 566 23196 572 23248
rect 624 23196 630 23248
rect 658 23196 664 23248
rect 716 23196 722 23248
rect 2332 23236 2360 23276
rect 2406 23264 2412 23316
rect 2464 23264 2470 23316
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2924 23276 2973 23304
rect 2924 23264 2930 23276
rect 2961 23273 2973 23276
rect 3007 23273 3019 23307
rect 2961 23267 3019 23273
rect 3418 23264 3424 23316
rect 3476 23304 3482 23316
rect 5718 23304 5724 23316
rect 3476 23276 5724 23304
rect 3476 23264 3482 23276
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 19886 23264 19892 23316
rect 19944 23264 19950 23316
rect 23753 23307 23811 23313
rect 23753 23273 23765 23307
rect 23799 23304 23811 23307
rect 23934 23304 23940 23316
rect 23799 23276 23940 23304
rect 23799 23273 23811 23276
rect 23753 23267 23811 23273
rect 23934 23264 23940 23276
rect 23992 23264 23998 23316
rect 24394 23264 24400 23316
rect 24452 23304 24458 23316
rect 25406 23304 25412 23316
rect 24452 23276 25412 23304
rect 24452 23264 24458 23276
rect 25406 23264 25412 23276
rect 25464 23264 25470 23316
rect 3510 23236 3516 23248
rect 2332 23208 3516 23236
rect 3510 23196 3516 23208
rect 3568 23196 3574 23248
rect 3970 23196 3976 23248
rect 4028 23236 4034 23248
rect 5626 23236 5632 23248
rect 4028 23208 5632 23236
rect 4028 23196 4034 23208
rect 5626 23196 5632 23208
rect 5684 23196 5690 23248
rect 18417 23239 18475 23245
rect 18417 23205 18429 23239
rect 18463 23205 18475 23239
rect 18417 23199 18475 23205
rect 2866 23168 2872 23180
rect 2700 23140 2872 23168
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 1671 23103 1729 23109
rect 1671 23069 1683 23103
rect 1717 23100 1729 23103
rect 2700 23100 2728 23140
rect 2866 23128 2872 23140
rect 2924 23168 2930 23180
rect 4614 23168 4620 23180
rect 2924 23140 4620 23168
rect 2924 23128 2930 23140
rect 4614 23128 4620 23140
rect 4672 23128 4678 23180
rect 7576 23140 7880 23168
rect 7576 23112 7604 23140
rect 1717 23072 2728 23100
rect 2777 23103 2835 23109
rect 1717 23069 1729 23072
rect 1671 23063 1729 23069
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 1302 22992 1308 23044
rect 1360 23032 1366 23044
rect 2792 23032 2820 23063
rect 1360 23004 2820 23032
rect 1360 22992 1366 23004
rect 2866 22992 2872 23044
rect 2924 23032 2930 23044
rect 3068 23032 3096 23063
rect 5258 23060 5264 23112
rect 5316 23100 5322 23112
rect 5442 23100 5448 23112
rect 5316 23072 5448 23100
rect 5316 23060 5322 23072
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 7466 23060 7472 23112
rect 7524 23060 7530 23112
rect 7558 23060 7564 23112
rect 7616 23060 7622 23112
rect 7852 23109 7880 23140
rect 7926 23128 7932 23180
rect 7984 23128 7990 23180
rect 11054 23128 11060 23180
rect 11112 23128 11118 23180
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 13262 23168 13268 23180
rect 12216 23140 13268 23168
rect 12216 23128 12222 23140
rect 13262 23128 13268 23140
rect 13320 23168 13326 23180
rect 13814 23168 13820 23180
rect 13320 23140 13820 23168
rect 13320 23128 13326 23140
rect 13814 23128 13820 23140
rect 13872 23168 13878 23180
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13872 23140 14105 23168
rect 13872 23128 13878 23140
rect 14093 23137 14105 23140
rect 14139 23137 14151 23171
rect 18432 23168 18460 23199
rect 19904 23177 19932 23264
rect 19337 23171 19395 23177
rect 18432 23140 19288 23168
rect 14093 23131 14151 23137
rect 7837 23103 7895 23109
rect 7837 23069 7849 23103
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 8205 23103 8263 23109
rect 8205 23069 8217 23103
rect 8251 23100 8263 23103
rect 8386 23100 8392 23112
rect 8251 23072 8392 23100
rect 8251 23069 8263 23072
rect 8205 23063 8263 23069
rect 8386 23060 8392 23072
rect 8444 23060 8450 23112
rect 10686 23060 10692 23112
rect 10744 23100 10750 23112
rect 10873 23103 10931 23109
rect 10873 23100 10885 23103
rect 10744 23072 10885 23100
rect 10744 23060 10750 23072
rect 10873 23069 10885 23072
rect 10919 23069 10931 23103
rect 10873 23063 10931 23069
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23100 11023 23103
rect 11238 23100 11244 23112
rect 11011 23072 11244 23100
rect 11011 23069 11023 23072
rect 10965 23063 11023 23069
rect 11238 23060 11244 23072
rect 11296 23060 11302 23112
rect 11333 23103 11391 23109
rect 11333 23069 11345 23103
rect 11379 23100 11391 23103
rect 11790 23100 11796 23112
rect 11379 23072 11796 23100
rect 11379 23069 11391 23072
rect 11333 23063 11391 23069
rect 11790 23060 11796 23072
rect 11848 23060 11854 23112
rect 14366 23100 14372 23112
rect 14327 23072 14372 23100
rect 14366 23060 14372 23072
rect 14424 23100 14430 23112
rect 14826 23100 14832 23112
rect 14424 23072 14832 23100
rect 14424 23060 14430 23072
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 18414 23060 18420 23112
rect 18472 23100 18478 23112
rect 19260 23109 19288 23140
rect 19337 23137 19349 23171
rect 19383 23168 19395 23171
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 19383 23140 19717 23168
rect 19383 23137 19395 23140
rect 19337 23131 19395 23137
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23137 19947 23171
rect 19889 23131 19947 23137
rect 18601 23103 18659 23109
rect 18601 23100 18613 23103
rect 18472 23072 18613 23100
rect 18472 23060 18478 23072
rect 18601 23069 18613 23072
rect 18647 23069 18659 23103
rect 18601 23063 18659 23069
rect 19245 23103 19303 23109
rect 19245 23069 19257 23103
rect 19291 23069 19303 23103
rect 19245 23063 19303 23069
rect 19610 23060 19616 23112
rect 19668 23060 19674 23112
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 20680 23072 21016 23100
rect 20680 23060 20686 23072
rect 7484 23032 7512 23060
rect 2924 23004 3096 23032
rect 3160 23004 7512 23032
rect 2924 22992 2930 23004
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 3160 22964 3188 23004
rect 8110 22992 8116 23044
rect 8168 22992 8174 23044
rect 10134 22992 10140 23044
rect 10192 23032 10198 23044
rect 11701 23035 11759 23041
rect 11701 23032 11713 23035
rect 10192 23004 11713 23032
rect 10192 22992 10198 23004
rect 11701 23001 11713 23004
rect 11747 23001 11759 23035
rect 11701 22995 11759 23001
rect 14274 22992 14280 23044
rect 14332 23032 14338 23044
rect 18046 23032 18052 23044
rect 14332 23004 18052 23032
rect 14332 22992 14338 23004
rect 18046 22992 18052 23004
rect 18104 22992 18110 23044
rect 19334 22992 19340 23044
rect 19392 23032 19398 23044
rect 20530 23032 20536 23044
rect 19392 23004 20536 23032
rect 19392 22992 19398 23004
rect 20530 22992 20536 23004
rect 20588 23032 20594 23044
rect 20870 23035 20928 23041
rect 20870 23032 20882 23035
rect 20588 23004 20882 23032
rect 20588 22992 20594 23004
rect 20870 23001 20882 23004
rect 20916 23001 20928 23035
rect 20988 23032 21016 23072
rect 21726 23060 21732 23112
rect 21784 23100 21790 23112
rect 22097 23103 22155 23109
rect 22097 23100 22109 23103
rect 21784 23072 22109 23100
rect 21784 23060 21790 23072
rect 22097 23069 22109 23072
rect 22143 23069 22155 23103
rect 22097 23063 22155 23069
rect 22370 23060 22376 23112
rect 22428 23060 22434 23112
rect 22646 23109 22652 23112
rect 22640 23100 22652 23109
rect 22607 23072 22652 23100
rect 22640 23063 22652 23072
rect 22646 23060 22652 23063
rect 22704 23060 22710 23112
rect 23750 23060 23756 23112
rect 23808 23100 23814 23112
rect 23937 23103 23995 23109
rect 23937 23100 23949 23103
rect 23808 23072 23949 23100
rect 23808 23060 23814 23072
rect 23937 23069 23949 23072
rect 23983 23069 23995 23103
rect 23937 23063 23995 23069
rect 22388 23032 22416 23060
rect 20988 23004 22416 23032
rect 20870 22995 20928 23001
rect 1728 22936 3188 22964
rect 3237 22967 3295 22973
rect 1728 22924 1734 22936
rect 3237 22933 3249 22967
rect 3283 22964 3295 22967
rect 6638 22964 6644 22976
rect 3283 22936 6644 22964
rect 3283 22933 3295 22936
rect 3237 22927 3295 22933
rect 6638 22924 6644 22936
rect 6696 22964 6702 22976
rect 7466 22964 7472 22976
rect 6696 22936 7472 22964
rect 6696 22924 6702 22936
rect 7466 22924 7472 22936
rect 7524 22924 7530 22976
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 10410 22964 10416 22976
rect 9456 22936 10416 22964
rect 9456 22924 9462 22936
rect 10410 22924 10416 22936
rect 10468 22924 10474 22976
rect 10597 22967 10655 22973
rect 10597 22933 10609 22967
rect 10643 22964 10655 22967
rect 11606 22964 11612 22976
rect 10643 22936 11612 22964
rect 10643 22933 10655 22936
rect 10597 22927 10655 22933
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 11885 22967 11943 22973
rect 11885 22933 11897 22967
rect 11931 22964 11943 22967
rect 14458 22964 14464 22976
rect 11931 22936 14464 22964
rect 11931 22933 11943 22936
rect 11885 22927 11943 22933
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 15105 22967 15163 22973
rect 15105 22933 15117 22967
rect 15151 22964 15163 22967
rect 15286 22964 15292 22976
rect 15151 22936 15292 22964
rect 15151 22933 15163 22936
rect 15105 22927 15163 22933
rect 15286 22924 15292 22936
rect 15344 22924 15350 22976
rect 19889 22967 19947 22973
rect 19889 22933 19901 22967
rect 19935 22964 19947 22967
rect 21266 22964 21272 22976
rect 19935 22936 21272 22964
rect 19935 22933 19947 22936
rect 19889 22927 19947 22933
rect 21266 22924 21272 22936
rect 21324 22924 21330 22976
rect 22005 22967 22063 22973
rect 22005 22933 22017 22967
rect 22051 22964 22063 22967
rect 22094 22964 22100 22976
rect 22051 22936 22100 22964
rect 22051 22933 22063 22936
rect 22005 22927 22063 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 22186 22924 22192 22976
rect 22244 22924 22250 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24026 22964 24032 22976
rect 23532 22936 24032 22964
rect 23532 22924 23538 22936
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 24121 22967 24179 22973
rect 24121 22933 24133 22967
rect 24167 22964 24179 22967
rect 25130 22964 25136 22976
rect 24167 22936 25136 22964
rect 24167 22933 24179 22936
rect 24121 22927 24179 22933
rect 25130 22924 25136 22936
rect 25188 22924 25194 22976
rect 1104 22874 25000 22896
rect 1104 22822 6884 22874
rect 6936 22822 6948 22874
rect 7000 22822 7012 22874
rect 7064 22822 7076 22874
rect 7128 22822 7140 22874
rect 7192 22822 12818 22874
rect 12870 22822 12882 22874
rect 12934 22822 12946 22874
rect 12998 22822 13010 22874
rect 13062 22822 13074 22874
rect 13126 22822 18752 22874
rect 18804 22822 18816 22874
rect 18868 22822 18880 22874
rect 18932 22822 18944 22874
rect 18996 22822 19008 22874
rect 19060 22822 24686 22874
rect 24738 22822 24750 22874
rect 24802 22822 24814 22874
rect 24866 22822 24878 22874
rect 24930 22822 24942 22874
rect 24994 22822 25000 22874
rect 1104 22800 25000 22822
rect 198 22720 204 22772
rect 256 22760 262 22772
rect 3050 22760 3056 22772
rect 256 22732 3056 22760
rect 256 22720 262 22732
rect 3050 22720 3056 22732
rect 3108 22720 3114 22772
rect 3142 22720 3148 22772
rect 3200 22720 3206 22772
rect 3234 22720 3240 22772
rect 3292 22760 3298 22772
rect 3789 22763 3847 22769
rect 3789 22760 3801 22763
rect 3292 22732 3801 22760
rect 3292 22720 3298 22732
rect 3789 22729 3801 22732
rect 3835 22729 3847 22763
rect 3789 22723 3847 22729
rect 4338 22720 4344 22772
rect 4396 22720 4402 22772
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 5626 22760 5632 22772
rect 4488 22732 5632 22760
rect 4488 22720 4494 22732
rect 5626 22720 5632 22732
rect 5684 22720 5690 22772
rect 6546 22720 6552 22772
rect 6604 22760 6610 22772
rect 7558 22760 7564 22772
rect 6604 22732 7564 22760
rect 6604 22720 6610 22732
rect 7558 22720 7564 22732
rect 7616 22720 7622 22772
rect 9214 22720 9220 22772
rect 9272 22760 9278 22772
rect 9677 22763 9735 22769
rect 9677 22760 9689 22763
rect 9272 22732 9689 22760
rect 9272 22720 9278 22732
rect 9677 22729 9689 22732
rect 9723 22729 9735 22763
rect 9677 22723 9735 22729
rect 11054 22720 11060 22772
rect 11112 22720 11118 22772
rect 13998 22720 14004 22772
rect 14056 22760 14062 22772
rect 16022 22760 16028 22772
rect 14056 22732 16028 22760
rect 14056 22720 14062 22732
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 19518 22720 19524 22772
rect 19576 22760 19582 22772
rect 20070 22760 20076 22772
rect 19576 22732 20076 22760
rect 19576 22720 19582 22732
rect 20070 22720 20076 22732
rect 20128 22720 20134 22772
rect 20530 22720 20536 22772
rect 20588 22720 20594 22772
rect 21085 22763 21143 22769
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 21726 22760 21732 22772
rect 21131 22732 21732 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 21726 22720 21732 22732
rect 21784 22720 21790 22772
rect 22020 22732 22416 22760
rect 1946 22692 1952 22704
rect 1686 22664 1952 22692
rect 1686 22663 1714 22664
rect 1655 22657 1714 22663
rect 1655 22623 1667 22657
rect 1701 22626 1714 22657
rect 1946 22652 1952 22664
rect 2004 22652 2010 22704
rect 1701 22623 1713 22626
rect 1655 22617 1713 22623
rect 2222 22584 2228 22636
rect 2280 22624 2286 22636
rect 2777 22627 2835 22633
rect 2777 22624 2789 22627
rect 2280 22596 2789 22624
rect 2280 22584 2286 22596
rect 2777 22593 2789 22596
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 3051 22627 3109 22633
rect 3051 22593 3063 22627
rect 3097 22624 3109 22627
rect 3160 22624 3188 22720
rect 4246 22692 4252 22704
rect 4080 22664 4252 22692
rect 4080 22624 4108 22664
rect 4246 22652 4252 22664
rect 4304 22652 4310 22704
rect 3097 22596 4108 22624
rect 4157 22627 4215 22633
rect 3097 22593 3109 22596
rect 3051 22587 3109 22593
rect 4157 22593 4169 22627
rect 4203 22624 4215 22627
rect 4356 22624 4384 22720
rect 4614 22652 4620 22704
rect 4672 22692 4678 22704
rect 12066 22692 12072 22704
rect 4672 22664 6316 22692
rect 4672 22652 4678 22664
rect 4203 22596 4384 22624
rect 4431 22627 4489 22633
rect 4203 22593 4215 22596
rect 4157 22587 4215 22593
rect 4431 22593 4443 22627
rect 4477 22624 4489 22627
rect 4890 22624 4896 22636
rect 4477 22596 4896 22624
rect 4477 22593 4489 22596
rect 4431 22587 4489 22593
rect 1394 22516 1400 22568
rect 1452 22516 1458 22568
rect 2792 22432 2820 22587
rect 2406 22380 2412 22432
rect 2464 22380 2470 22432
rect 2774 22380 2780 22432
rect 2832 22380 2838 22432
rect 4172 22420 4200 22587
rect 4890 22584 4896 22596
rect 4948 22584 4954 22636
rect 6178 22584 6184 22636
rect 6236 22584 6242 22636
rect 6288 22624 6316 22664
rect 8956 22664 12072 22692
rect 8956 22663 8984 22664
rect 8923 22657 8984 22663
rect 6607 22627 6665 22633
rect 6607 22624 6619 22627
rect 6288 22596 6619 22624
rect 6607 22593 6619 22596
rect 6653 22593 6665 22627
rect 8923 22623 8935 22657
rect 8969 22626 8984 22657
rect 12066 22652 12072 22664
rect 12124 22652 12130 22704
rect 16868 22692 16896 22720
rect 16500 22664 16896 22692
rect 8969 22623 8981 22626
rect 8923 22617 8981 22623
rect 6607 22587 6665 22593
rect 10318 22584 10324 22636
rect 10376 22624 10382 22636
rect 10376 22596 15608 22624
rect 10376 22584 10382 22596
rect 6196 22556 6224 22584
rect 6365 22559 6423 22565
rect 6365 22556 6377 22559
rect 6196 22528 6377 22556
rect 6365 22525 6377 22528
rect 6411 22525 6423 22559
rect 6365 22519 6423 22525
rect 8294 22516 8300 22568
rect 8352 22556 8358 22568
rect 8665 22559 8723 22565
rect 8665 22556 8677 22559
rect 8352 22528 8677 22556
rect 8352 22516 8358 22528
rect 8665 22525 8677 22528
rect 8711 22525 8723 22559
rect 8665 22519 8723 22525
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22525 10103 22559
rect 10045 22519 10103 22525
rect 7282 22448 7288 22500
rect 7340 22488 7346 22500
rect 8110 22488 8116 22500
rect 7340 22460 8116 22488
rect 7340 22448 7346 22460
rect 8110 22448 8116 22460
rect 8168 22448 8174 22500
rect 4614 22420 4620 22432
rect 4172 22392 4620 22420
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 5166 22380 5172 22432
rect 5224 22380 5230 22432
rect 6730 22380 6736 22432
rect 6788 22420 6794 22432
rect 7377 22423 7435 22429
rect 7377 22420 7389 22423
rect 6788 22392 7389 22420
rect 6788 22380 6794 22392
rect 7377 22389 7389 22392
rect 7423 22389 7435 22423
rect 10060 22420 10088 22519
rect 10962 22516 10968 22568
rect 11020 22516 11026 22568
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 11330 22556 11336 22568
rect 11112 22528 11336 22556
rect 11112 22516 11118 22528
rect 11330 22516 11336 22528
rect 11388 22516 11394 22568
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 12158 22556 12164 22568
rect 11756 22528 12164 22556
rect 11756 22516 11762 22528
rect 12158 22516 12164 22528
rect 12216 22516 12222 22568
rect 12342 22516 12348 22568
rect 12400 22556 12406 22568
rect 15470 22556 15476 22568
rect 12400 22528 15476 22556
rect 12400 22516 12406 22528
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 10980 22420 11008 22516
rect 14182 22448 14188 22500
rect 14240 22488 14246 22500
rect 14366 22488 14372 22500
rect 14240 22460 14372 22488
rect 14240 22448 14246 22460
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 11606 22420 11612 22432
rect 10060 22392 11612 22420
rect 7377 22383 7435 22389
rect 11606 22380 11612 22392
rect 11664 22380 11670 22432
rect 14826 22380 14832 22432
rect 14884 22380 14890 22432
rect 15580 22420 15608 22596
rect 15654 22516 15660 22568
rect 15712 22516 15718 22568
rect 16500 22556 16528 22664
rect 16574 22584 16580 22636
rect 16632 22624 16638 22636
rect 16850 22624 16856 22636
rect 16632 22596 16856 22624
rect 16632 22584 16638 22596
rect 16850 22584 16856 22596
rect 16908 22584 16914 22636
rect 17770 22633 17776 22636
rect 17727 22627 17776 22633
rect 17727 22593 17739 22627
rect 17773 22593 17776 22627
rect 17727 22587 17776 22593
rect 17770 22584 17776 22587
rect 17828 22584 17834 22636
rect 20548 22624 20576 22720
rect 22020 22636 22048 22732
rect 22278 22692 22284 22704
rect 22204 22664 22284 22692
rect 22095 22637 22153 22643
rect 21269 22627 21327 22633
rect 21269 22624 21281 22627
rect 20548 22596 21281 22624
rect 21269 22593 21281 22596
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21450 22584 21456 22636
rect 21508 22584 21514 22636
rect 21637 22627 21695 22633
rect 21637 22593 21649 22627
rect 21683 22624 21695 22627
rect 21726 22624 21732 22636
rect 21683 22596 21732 22624
rect 21683 22593 21695 22596
rect 21637 22587 21695 22593
rect 21726 22584 21732 22596
rect 21784 22584 21790 22636
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22624 21879 22627
rect 22002 22624 22008 22636
rect 21867 22596 22008 22624
rect 21867 22593 21879 22596
rect 21821 22587 21879 22593
rect 22002 22584 22008 22596
rect 22060 22584 22066 22636
rect 22095 22603 22107 22637
rect 22141 22634 22153 22637
rect 22204 22634 22232 22664
rect 22278 22652 22284 22664
rect 22336 22652 22342 22704
rect 22141 22606 22232 22634
rect 22388 22624 22416 22732
rect 23198 22720 23204 22772
rect 23256 22760 23262 22772
rect 24213 22763 24271 22769
rect 24213 22760 24225 22763
rect 23256 22732 24225 22760
rect 23256 22720 23262 22732
rect 24213 22729 24225 22732
rect 24259 22729 24271 22763
rect 24213 22723 24271 22729
rect 23842 22652 23848 22704
rect 23900 22692 23906 22704
rect 24486 22692 24492 22704
rect 23900 22664 24492 22692
rect 23900 22652 23906 22664
rect 24486 22652 24492 22664
rect 24544 22652 24550 22704
rect 22554 22624 22560 22636
rect 22141 22603 22153 22606
rect 22095 22597 22153 22603
rect 22388 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22624 22618 22636
rect 23201 22627 23259 22633
rect 23201 22624 23213 22627
rect 22612 22596 23213 22624
rect 22612 22584 22618 22596
rect 23201 22593 23213 22596
rect 23247 22593 23259 22627
rect 23201 22587 23259 22593
rect 23474 22584 23480 22636
rect 23532 22584 23538 22636
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16500 22528 16681 22556
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 17589 22559 17647 22565
rect 17589 22556 17601 22559
rect 16669 22519 16727 22525
rect 16776 22528 17601 22556
rect 15672 22488 15700 22516
rect 16776 22488 16804 22528
rect 17589 22525 17601 22528
rect 17635 22525 17647 22559
rect 17589 22519 17647 22525
rect 17862 22516 17868 22568
rect 17920 22516 17926 22568
rect 15672 22460 16804 22488
rect 17310 22448 17316 22500
rect 17368 22448 17374 22500
rect 16666 22420 16672 22432
rect 15580 22392 16672 22420
rect 16666 22380 16672 22392
rect 16724 22420 16730 22432
rect 17218 22420 17224 22432
rect 16724 22392 17224 22420
rect 16724 22380 16730 22392
rect 17218 22380 17224 22392
rect 17276 22380 17282 22432
rect 18506 22380 18512 22432
rect 18564 22380 18570 22432
rect 21545 22423 21603 22429
rect 21545 22389 21557 22423
rect 21591 22420 21603 22423
rect 22278 22420 22284 22432
rect 21591 22392 22284 22420
rect 21591 22389 21603 22392
rect 21545 22383 21603 22389
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 22830 22380 22836 22432
rect 22888 22380 22894 22432
rect 1104 22330 24840 22352
rect 1104 22278 3917 22330
rect 3969 22278 3981 22330
rect 4033 22278 4045 22330
rect 4097 22278 4109 22330
rect 4161 22278 4173 22330
rect 4225 22278 9851 22330
rect 9903 22278 9915 22330
rect 9967 22278 9979 22330
rect 10031 22278 10043 22330
rect 10095 22278 10107 22330
rect 10159 22278 15785 22330
rect 15837 22278 15849 22330
rect 15901 22278 15913 22330
rect 15965 22278 15977 22330
rect 16029 22278 16041 22330
rect 16093 22278 21719 22330
rect 21771 22278 21783 22330
rect 21835 22278 21847 22330
rect 21899 22278 21911 22330
rect 21963 22278 21975 22330
rect 22027 22278 24840 22330
rect 1104 22256 24840 22278
rect 3050 22176 3056 22228
rect 3108 22176 3114 22228
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 3510 22216 3516 22228
rect 3292 22188 3516 22216
rect 3292 22176 3298 22188
rect 3510 22176 3516 22188
rect 3568 22176 3574 22228
rect 3602 22176 3608 22228
rect 3660 22176 3666 22228
rect 3786 22176 3792 22228
rect 3844 22216 3850 22228
rect 3973 22219 4031 22225
rect 3973 22216 3985 22219
rect 3844 22188 3985 22216
rect 3844 22176 3850 22188
rect 3973 22185 3985 22188
rect 4019 22185 4031 22219
rect 9030 22216 9036 22228
rect 3973 22179 4031 22185
rect 6012 22188 9036 22216
rect 3620 22148 3648 22176
rect 6012 22157 6040 22188
rect 9030 22176 9036 22188
rect 9088 22176 9094 22228
rect 9122 22176 9128 22228
rect 9180 22216 9186 22228
rect 9490 22216 9496 22228
rect 9180 22188 9496 22216
rect 9180 22176 9186 22188
rect 9490 22176 9496 22188
rect 9548 22176 9554 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10870 22216 10876 22228
rect 10008 22188 10876 22216
rect 10008 22176 10014 22188
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 11057 22219 11115 22225
rect 11057 22185 11069 22219
rect 11103 22216 11115 22219
rect 19150 22216 19156 22228
rect 11103 22188 11468 22216
rect 11103 22185 11115 22188
rect 11057 22179 11115 22185
rect 5997 22151 6055 22157
rect 3620 22120 4476 22148
rect 2314 22040 2320 22092
rect 2372 22040 2378 22092
rect 3160 22052 4016 22080
rect 2133 22015 2191 22021
rect 2133 21981 2145 22015
rect 2179 22012 2191 22015
rect 2406 22012 2412 22024
rect 2179 21984 2412 22012
rect 2179 21981 2191 21984
rect 2133 21975 2191 21981
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 22012 2559 22015
rect 3160 22012 3188 22052
rect 2547 21984 3188 22012
rect 3237 22015 3295 22021
rect 2547 21981 2559 21984
rect 2501 21975 2559 21981
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 3602 22012 3608 22024
rect 3283 21984 3608 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3602 21972 3608 21984
rect 3660 21972 3666 22024
rect 3789 22015 3847 22021
rect 3789 21981 3801 22015
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 1762 21904 1768 21956
rect 1820 21904 1826 21956
rect 2038 21904 2044 21956
rect 2096 21904 2102 21956
rect 3804 21944 3832 21975
rect 3988 21956 4016 22052
rect 4448 22012 4476 22120
rect 5997 22117 6009 22151
rect 6043 22117 6055 22151
rect 5997 22111 6055 22117
rect 6178 22108 6184 22160
rect 6236 22108 6242 22160
rect 6546 22108 6552 22160
rect 6604 22108 6610 22160
rect 7650 22108 7656 22160
rect 7708 22148 7714 22160
rect 7708 22120 8064 22148
rect 7708 22108 7714 22120
rect 5166 22040 5172 22092
rect 5224 22040 5230 22092
rect 6196 22080 6224 22108
rect 6641 22083 6699 22089
rect 6641 22080 6653 22083
rect 6196 22052 6653 22080
rect 6564 22024 6592 22052
rect 6641 22049 6653 22052
rect 6687 22049 6699 22083
rect 6641 22043 6699 22049
rect 8036 22024 8064 22120
rect 11440 22066 11468 22188
rect 12912 22188 19156 22216
rect 12912 22157 12940 22188
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 20622 22216 20628 22228
rect 19260 22188 20628 22216
rect 12897 22151 12955 22157
rect 12897 22117 12909 22151
rect 12943 22117 12955 22151
rect 12897 22111 12955 22117
rect 17310 22108 17316 22160
rect 17368 22108 17374 22160
rect 18506 22108 18512 22160
rect 18564 22108 18570 22160
rect 14734 22040 14740 22092
rect 14792 22040 14798 22092
rect 14826 22040 14832 22092
rect 14884 22080 14890 22092
rect 15013 22083 15071 22089
rect 15013 22080 15025 22083
rect 14884 22052 15025 22080
rect 14884 22040 14890 22052
rect 15013 22049 15025 22052
rect 15059 22049 15071 22083
rect 15013 22043 15071 22049
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 4985 22015 5043 22021
rect 4985 22012 4997 22015
rect 4448 21984 4997 22012
rect 4985 21981 4997 21984
rect 5031 21981 5043 22015
rect 4985 21975 5043 21981
rect 5074 21972 5080 22024
rect 5132 21972 5138 22024
rect 5258 21972 5264 22024
rect 5316 22012 5322 22024
rect 5316 21984 6040 22012
rect 5316 21972 5322 21984
rect 2746 21916 3832 21944
rect 1210 21836 1216 21888
rect 1268 21876 1274 21888
rect 2746 21876 2774 21916
rect 3970 21904 3976 21956
rect 4028 21904 4034 21956
rect 5166 21904 5172 21956
rect 5224 21944 5230 21956
rect 5445 21947 5503 21953
rect 5445 21944 5457 21947
rect 5224 21916 5457 21944
rect 5224 21904 5230 21916
rect 5445 21913 5457 21916
rect 5491 21944 5503 21947
rect 5626 21944 5632 21956
rect 5491 21916 5632 21944
rect 5491 21913 5503 21916
rect 5445 21907 5503 21913
rect 5626 21904 5632 21916
rect 5684 21904 5690 21956
rect 6012 21944 6040 21984
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6915 22015 6973 22021
rect 6915 21981 6927 22015
rect 6961 22012 6973 22015
rect 7650 22012 7656 22024
rect 6961 21984 7656 22012
rect 6961 21981 6973 21984
rect 6915 21975 6973 21981
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 8018 21972 8024 22024
rect 8076 21972 8082 22024
rect 9582 21972 9588 22024
rect 9640 22008 9646 22024
rect 10042 22012 10048 22024
rect 9692 22008 10048 22012
rect 9640 21984 10048 22008
rect 9640 21980 9720 21984
rect 9640 21972 9646 21980
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10319 22015 10377 22021
rect 10319 21981 10331 22015
rect 10365 22012 10377 22015
rect 10410 22012 10416 22024
rect 10365 21984 10416 22012
rect 10365 21981 10377 21984
rect 10319 21975 10377 21981
rect 10410 21972 10416 21984
rect 10468 21972 10474 22024
rect 13354 22012 13360 22024
rect 11072 21984 13360 22012
rect 11072 21944 11100 21984
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14093 21975 14151 21981
rect 14200 21984 14289 22012
rect 6012 21916 9674 21944
rect 1268 21848 2774 21876
rect 2869 21879 2927 21885
rect 1268 21836 1274 21848
rect 2869 21845 2881 21879
rect 2915 21876 2927 21879
rect 3050 21876 3056 21888
rect 2915 21848 3056 21876
rect 2915 21845 2927 21848
rect 2869 21839 2927 21845
rect 3050 21836 3056 21848
rect 3108 21836 3114 21888
rect 3421 21879 3479 21885
rect 3421 21845 3433 21879
rect 3467 21876 3479 21879
rect 3988 21876 4016 21904
rect 3467 21848 4016 21876
rect 3467 21845 3479 21848
rect 3421 21839 3479 21845
rect 4062 21836 4068 21888
rect 4120 21876 4126 21888
rect 4706 21876 4712 21888
rect 4120 21848 4712 21876
rect 4120 21836 4126 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5813 21879 5871 21885
rect 5813 21845 5825 21879
rect 5859 21876 5871 21879
rect 5994 21876 6000 21888
rect 5859 21848 6000 21876
rect 5859 21845 5871 21848
rect 5813 21839 5871 21845
rect 5994 21836 6000 21848
rect 6052 21836 6058 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7432 21848 7665 21876
rect 7432 21836 7438 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 9646 21876 9674 21916
rect 9876 21916 11100 21944
rect 11164 21916 11744 21944
rect 9876 21876 9904 21916
rect 9646 21848 9904 21876
rect 7653 21839 7711 21845
rect 10594 21836 10600 21888
rect 10652 21876 10658 21888
rect 11164 21876 11192 21916
rect 10652 21848 11192 21876
rect 10652 21836 10658 21848
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 11609 21879 11667 21885
rect 11609 21876 11621 21879
rect 11296 21848 11621 21876
rect 11296 21836 11302 21848
rect 11609 21845 11621 21848
rect 11655 21845 11667 21879
rect 11716 21876 11744 21916
rect 11882 21904 11888 21956
rect 11940 21904 11946 21956
rect 11974 21904 11980 21956
rect 12032 21904 12038 21956
rect 12158 21904 12164 21956
rect 12216 21944 12222 21956
rect 12345 21947 12403 21953
rect 12345 21944 12357 21947
rect 12216 21916 12357 21944
rect 12216 21904 12222 21916
rect 12345 21913 12357 21916
rect 12391 21944 12403 21947
rect 14108 21944 14136 21975
rect 12391 21916 14136 21944
rect 12391 21913 12403 21916
rect 12345 21907 12403 21913
rect 12713 21879 12771 21885
rect 12713 21876 12725 21879
rect 11716 21848 12725 21876
rect 11609 21839 11667 21845
rect 12713 21845 12725 21848
rect 12759 21876 12771 21879
rect 14200 21876 14228 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 15102 21972 15108 22024
rect 15160 22021 15166 22024
rect 15160 22015 15188 22021
rect 15176 21981 15188 22015
rect 15160 21975 15188 21981
rect 15160 21972 15166 21975
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16301 22015 16359 22021
rect 16301 22012 16313 22015
rect 16172 21984 16313 22012
rect 16172 21972 16178 21984
rect 16301 21981 16313 21984
rect 16347 21981 16359 22015
rect 16574 22012 16580 22024
rect 16535 21984 16580 22012
rect 16301 21975 16359 21981
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 18417 22015 18475 22021
rect 16684 21984 17632 22012
rect 16684 21944 16712 21984
rect 15764 21916 16712 21944
rect 12759 21848 14228 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 14826 21836 14832 21888
rect 14884 21876 14890 21888
rect 15764 21876 15792 21916
rect 17218 21904 17224 21956
rect 17276 21944 17282 21956
rect 17494 21944 17500 21956
rect 17276 21916 17500 21944
rect 17276 21904 17282 21916
rect 17494 21904 17500 21916
rect 17552 21904 17558 21956
rect 17604 21944 17632 21984
rect 18417 21981 18429 22015
rect 18463 22012 18475 22015
rect 18524 22012 18552 22108
rect 19260 22024 19288 22188
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 22002 22216 22008 22228
rect 20772 22188 22008 22216
rect 20772 22176 20778 22188
rect 22002 22176 22008 22188
rect 22060 22176 22066 22228
rect 22097 22219 22155 22225
rect 22097 22185 22109 22219
rect 22143 22216 22155 22219
rect 22186 22216 22192 22228
rect 22143 22188 22192 22216
rect 22143 22185 22155 22188
rect 22097 22179 22155 22185
rect 22186 22176 22192 22188
rect 22244 22176 22250 22228
rect 22830 22216 22836 22228
rect 22296 22188 22836 22216
rect 21450 22108 21456 22160
rect 21508 22148 21514 22160
rect 22296 22148 22324 22188
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 23201 22219 23259 22225
rect 23201 22185 23213 22219
rect 23247 22216 23259 22219
rect 23566 22216 23572 22228
rect 23247 22188 23572 22216
rect 23247 22185 23259 22188
rect 23201 22179 23259 22185
rect 23566 22176 23572 22188
rect 23624 22176 23630 22228
rect 21508 22120 22324 22148
rect 22373 22151 22431 22157
rect 21508 22108 21514 22120
rect 20254 22040 20260 22092
rect 20312 22080 20318 22092
rect 20312 22052 21128 22080
rect 20312 22040 20318 22052
rect 19242 22012 19248 22024
rect 18463 21984 18552 22012
rect 19203 21984 19248 22012
rect 18463 21981 18475 21984
rect 18417 21975 18475 21981
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19512 22015 19570 22021
rect 19512 21981 19524 22015
rect 19558 22012 19570 22015
rect 19794 22012 19800 22024
rect 19558 21984 19800 22012
rect 19558 21981 19570 21984
rect 19512 21975 19570 21981
rect 19794 21972 19800 21984
rect 19852 22012 19858 22024
rect 20070 22012 20076 22024
rect 19852 21984 20076 22012
rect 19852 21972 19858 21984
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 20806 21972 20812 22024
rect 20864 21972 20870 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 19886 21944 19892 21956
rect 17604 21916 19892 21944
rect 19886 21904 19892 21916
rect 19944 21944 19950 21956
rect 20346 21944 20352 21956
rect 19944 21916 20352 21944
rect 19944 21904 19950 21916
rect 20346 21904 20352 21916
rect 20404 21904 20410 21956
rect 20714 21904 20720 21956
rect 20772 21944 20778 21956
rect 21008 21944 21036 21975
rect 20772 21916 21036 21944
rect 21100 21944 21128 22052
rect 22020 22021 22048 22120
rect 22373 22117 22385 22151
rect 22419 22148 22431 22151
rect 22462 22148 22468 22160
rect 22419 22120 22468 22148
rect 22419 22117 22431 22120
rect 22373 22111 22431 22117
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 22278 22040 22284 22092
rect 22336 22040 22342 22092
rect 23382 22040 23388 22092
rect 23440 22040 23446 22092
rect 24026 22080 24032 22092
rect 23584 22052 24032 22080
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 21981 22063 22015
rect 22005 21975 22063 21981
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22152 21984 22569 22012
rect 22152 21972 22158 21984
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 22557 21975 22615 21981
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 23584 22021 23612 22052
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23750 21972 23756 22024
rect 23808 21972 23814 22024
rect 24210 21972 24216 22024
rect 24268 21972 24274 22024
rect 23474 21944 23480 21956
rect 21100 21916 23480 21944
rect 20772 21904 20778 21916
rect 23474 21904 23480 21916
rect 23532 21904 23538 21956
rect 14884 21848 15792 21876
rect 15933 21879 15991 21885
rect 14884 21836 14890 21848
rect 15933 21845 15945 21879
rect 15979 21876 15991 21879
rect 17770 21876 17776 21888
rect 15979 21848 17776 21876
rect 15979 21845 15991 21848
rect 15933 21839 15991 21845
rect 17770 21836 17776 21848
rect 17828 21836 17834 21888
rect 18233 21879 18291 21885
rect 18233 21845 18245 21879
rect 18279 21876 18291 21879
rect 18598 21876 18604 21888
rect 18279 21848 18604 21876
rect 18279 21845 18291 21848
rect 18233 21839 18291 21845
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 20625 21879 20683 21885
rect 20625 21845 20637 21879
rect 20671 21876 20683 21879
rect 20898 21876 20904 21888
rect 20671 21848 20904 21876
rect 20671 21845 20683 21848
rect 20625 21839 20683 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 20990 21836 20996 21888
rect 21048 21836 21054 21888
rect 22278 21836 22284 21888
rect 22336 21836 22342 21888
rect 23382 21836 23388 21888
rect 23440 21836 23446 21888
rect 23768 21876 23796 21972
rect 23937 21947 23995 21953
rect 23937 21913 23949 21947
rect 23983 21944 23995 21947
rect 25130 21944 25136 21956
rect 23983 21916 25136 21944
rect 23983 21913 23995 21916
rect 23937 21907 23995 21913
rect 25130 21904 25136 21916
rect 25188 21904 25194 21956
rect 24029 21879 24087 21885
rect 24029 21876 24041 21879
rect 23768 21848 24041 21876
rect 24029 21845 24041 21848
rect 24075 21845 24087 21879
rect 24029 21839 24087 21845
rect 1104 21786 25000 21808
rect 1104 21734 6884 21786
rect 6936 21734 6948 21786
rect 7000 21734 7012 21786
rect 7064 21734 7076 21786
rect 7128 21734 7140 21786
rect 7192 21734 12818 21786
rect 12870 21734 12882 21786
rect 12934 21734 12946 21786
rect 12998 21734 13010 21786
rect 13062 21734 13074 21786
rect 13126 21734 18752 21786
rect 18804 21734 18816 21786
rect 18868 21734 18880 21786
rect 18932 21734 18944 21786
rect 18996 21734 19008 21786
rect 19060 21734 24686 21786
rect 24738 21734 24750 21786
rect 24802 21734 24814 21786
rect 24866 21734 24878 21786
rect 24930 21734 24942 21786
rect 24994 21734 25000 21786
rect 1104 21712 25000 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1360 21644 1808 21672
rect 1360 21632 1366 21644
rect 1670 21575 1676 21616
rect 1655 21569 1676 21575
rect 1394 21496 1400 21548
rect 1452 21496 1458 21548
rect 1655 21535 1667 21569
rect 1728 21564 1734 21616
rect 1780 21604 1808 21644
rect 2314 21632 2320 21684
rect 2372 21672 2378 21684
rect 2409 21675 2467 21681
rect 2409 21672 2421 21675
rect 2372 21644 2421 21672
rect 2372 21632 2378 21644
rect 2409 21641 2421 21644
rect 2455 21641 2467 21675
rect 2409 21635 2467 21641
rect 2590 21632 2596 21684
rect 2648 21672 2654 21684
rect 2961 21675 3019 21681
rect 2961 21672 2973 21675
rect 2648 21644 2973 21672
rect 2648 21632 2654 21644
rect 2961 21641 2973 21644
rect 3007 21672 3019 21675
rect 4062 21672 4068 21684
rect 3007 21644 4068 21672
rect 3007 21641 3019 21644
rect 2961 21635 3019 21641
rect 4062 21632 4068 21644
rect 4120 21632 4126 21684
rect 4614 21632 4620 21684
rect 4672 21632 4678 21684
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5721 21675 5779 21681
rect 5721 21672 5733 21675
rect 5132 21644 5733 21672
rect 5132 21632 5138 21644
rect 5721 21641 5733 21644
rect 5767 21641 5779 21675
rect 5721 21635 5779 21641
rect 6086 21632 6092 21684
rect 6144 21672 6150 21684
rect 8938 21672 8944 21684
rect 6144 21644 7696 21672
rect 6144 21632 6150 21644
rect 1780 21576 2820 21604
rect 1701 21538 1716 21564
rect 2792 21545 2820 21576
rect 2777 21539 2835 21545
rect 1701 21535 1713 21538
rect 1655 21529 1713 21535
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 4632 21536 4660 21632
rect 6362 21564 6368 21616
rect 6420 21604 6426 21616
rect 6549 21607 6607 21613
rect 6549 21604 6561 21607
rect 6420 21576 6561 21604
rect 6420 21564 6426 21576
rect 6549 21573 6561 21576
rect 6595 21573 6607 21607
rect 6549 21567 6607 21573
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 6825 21607 6883 21613
rect 6825 21604 6837 21607
rect 6696 21576 6837 21604
rect 6696 21564 6702 21576
rect 6825 21573 6837 21576
rect 6871 21573 6883 21607
rect 6825 21567 6883 21573
rect 6917 21607 6975 21613
rect 6917 21573 6929 21607
rect 6963 21604 6975 21607
rect 7374 21604 7380 21616
rect 6963 21576 7380 21604
rect 6963 21573 6975 21576
rect 6917 21567 6975 21573
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 7466 21564 7472 21616
rect 7524 21564 7530 21616
rect 7668 21613 7696 21644
rect 8404 21644 8944 21672
rect 8404 21616 8432 21644
rect 8938 21632 8944 21644
rect 8996 21632 9002 21684
rect 9122 21632 9128 21684
rect 9180 21672 9186 21684
rect 9585 21675 9643 21681
rect 9585 21672 9597 21675
rect 9180 21644 9597 21672
rect 9180 21632 9186 21644
rect 9585 21641 9597 21644
rect 9631 21641 9643 21675
rect 9585 21635 9643 21641
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9732 21644 9781 21672
rect 9732 21632 9738 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 10686 21632 10692 21684
rect 10744 21672 10750 21684
rect 10962 21672 10968 21684
rect 10744 21644 10968 21672
rect 10744 21632 10750 21644
rect 10962 21632 10968 21644
rect 11020 21632 11026 21684
rect 11974 21632 11980 21684
rect 12032 21672 12038 21684
rect 12805 21675 12863 21681
rect 12805 21672 12817 21675
rect 12032 21644 12817 21672
rect 12032 21632 12038 21644
rect 12805 21641 12817 21644
rect 12851 21641 12863 21675
rect 12805 21635 12863 21641
rect 14277 21675 14335 21681
rect 14277 21641 14289 21675
rect 14323 21672 14335 21675
rect 14734 21672 14740 21684
rect 14323 21644 14740 21672
rect 14323 21641 14335 21644
rect 14277 21635 14335 21641
rect 14734 21632 14740 21644
rect 14792 21632 14798 21684
rect 20254 21672 20260 21684
rect 14844 21644 20260 21672
rect 7653 21607 7711 21613
rect 7653 21573 7665 21607
rect 7699 21573 7711 21607
rect 7653 21567 7711 21573
rect 8386 21564 8392 21616
rect 8444 21564 8450 21616
rect 8481 21607 8539 21613
rect 8481 21573 8493 21607
rect 8527 21604 8539 21607
rect 11054 21604 11060 21616
rect 8527 21576 11060 21604
rect 8527 21573 8539 21576
rect 8481 21567 8539 21573
rect 11054 21564 11060 21576
rect 11112 21604 11118 21616
rect 12158 21604 12164 21616
rect 11112 21576 12164 21604
rect 11112 21564 11118 21576
rect 12158 21564 12164 21576
rect 12216 21564 12222 21616
rect 14844 21604 14872 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20864 21644 20913 21672
rect 20864 21632 20870 21644
rect 20901 21641 20913 21644
rect 20947 21641 20959 21675
rect 20901 21635 20959 21641
rect 13464 21576 14872 21604
rect 4709 21539 4767 21545
rect 4709 21536 4721 21539
rect 4632 21508 4721 21536
rect 3053 21499 3111 21505
rect 4709 21505 4721 21508
rect 4755 21505 4767 21539
rect 4709 21499 4767 21505
rect 4983 21539 5041 21545
rect 4983 21505 4995 21539
rect 5029 21536 5041 21539
rect 7190 21536 7196 21548
rect 5029 21508 7196 21536
rect 5029 21505 5041 21508
rect 4983 21499 5041 21505
rect 3068 21400 3096 21499
rect 7190 21496 7196 21508
rect 7248 21496 7254 21548
rect 7285 21539 7343 21545
rect 7285 21505 7297 21539
rect 7331 21536 7343 21539
rect 7484 21536 7512 21564
rect 7331 21508 7512 21536
rect 7331 21505 7343 21508
rect 7285 21499 7343 21505
rect 8754 21496 8760 21548
rect 8812 21496 8818 21548
rect 8846 21496 8852 21548
rect 8904 21496 8910 21548
rect 8938 21496 8944 21548
rect 8996 21536 9002 21548
rect 9217 21539 9275 21545
rect 9217 21536 9229 21539
rect 8996 21508 9229 21536
rect 8996 21496 9002 21508
rect 9217 21505 9229 21508
rect 9263 21505 9275 21539
rect 12035 21539 12093 21545
rect 12035 21536 12047 21539
rect 9217 21499 9275 21505
rect 9600 21508 12047 21536
rect 8484 21480 8536 21486
rect 9600 21480 9628 21508
rect 12035 21505 12047 21508
rect 12081 21536 12093 21539
rect 13464 21536 13492 21576
rect 15194 21564 15200 21616
rect 15252 21604 15258 21616
rect 16298 21604 16304 21616
rect 15252 21576 16304 21604
rect 15252 21564 15258 21576
rect 12081 21508 13492 21536
rect 12081 21505 12093 21508
rect 12035 21499 12093 21505
rect 13538 21496 13544 21548
rect 13596 21536 13602 21548
rect 15378 21545 15406 21576
rect 16298 21564 16304 21576
rect 16356 21564 16362 21616
rect 16758 21564 16764 21616
rect 16816 21564 16822 21616
rect 18598 21564 18604 21616
rect 18656 21604 18662 21616
rect 18656 21576 18920 21604
rect 18656 21564 18662 21576
rect 15363 21539 15421 21545
rect 13596 21508 13639 21536
rect 13596 21496 13602 21508
rect 15363 21505 15375 21539
rect 15409 21505 15421 21539
rect 15363 21499 15421 21505
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16776 21536 16804 21564
rect 16715 21508 16804 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 6730 21428 6736 21480
rect 6788 21428 6794 21480
rect 9582 21428 9588 21480
rect 9640 21428 9646 21480
rect 9858 21428 9864 21480
rect 9916 21468 9922 21480
rect 10594 21468 10600 21480
rect 9916 21440 10600 21468
rect 9916 21428 9922 21440
rect 10594 21428 10600 21440
rect 10652 21428 10658 21480
rect 11790 21428 11796 21480
rect 11848 21428 11854 21480
rect 13262 21428 13268 21480
rect 13320 21428 13326 21480
rect 15105 21471 15163 21477
rect 15105 21468 15117 21471
rect 14660 21440 15117 21468
rect 8484 21422 8536 21428
rect 2056 21372 3096 21400
rect 3237 21403 3295 21409
rect 1302 21292 1308 21344
rect 1360 21332 1366 21344
rect 2056 21332 2084 21372
rect 3237 21369 3249 21403
rect 3283 21400 3295 21403
rect 4614 21400 4620 21412
rect 3283 21372 4620 21400
rect 3283 21369 3295 21372
rect 3237 21363 3295 21369
rect 4614 21360 4620 21372
rect 4672 21360 4678 21412
rect 5626 21360 5632 21412
rect 5684 21400 5690 21412
rect 5902 21400 5908 21412
rect 5684 21372 5908 21400
rect 5684 21360 5690 21372
rect 5902 21360 5908 21372
rect 5960 21360 5966 21412
rect 7834 21360 7840 21412
rect 7892 21360 7898 21412
rect 10042 21360 10048 21412
rect 10100 21400 10106 21412
rect 10410 21400 10416 21412
rect 10100 21372 10416 21400
rect 10100 21360 10106 21372
rect 10410 21360 10416 21372
rect 10468 21400 10474 21412
rect 11808 21400 11836 21428
rect 10468 21372 11836 21400
rect 10468 21360 10474 21372
rect 1360 21304 2084 21332
rect 1360 21292 1366 21304
rect 4798 21292 4804 21344
rect 4856 21332 4862 21344
rect 5994 21332 6000 21344
rect 4856 21304 6000 21332
rect 4856 21292 4862 21304
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 10686 21332 10692 21344
rect 10376 21304 10692 21332
rect 10376 21292 10382 21304
rect 10686 21292 10692 21304
rect 10744 21292 10750 21344
rect 13280 21332 13308 21428
rect 14366 21332 14372 21344
rect 13280 21304 14372 21332
rect 14366 21292 14372 21304
rect 14424 21332 14430 21344
rect 14660 21332 14688 21440
rect 15105 21437 15117 21440
rect 15151 21437 15163 21471
rect 15105 21431 15163 21437
rect 16114 21428 16120 21480
rect 16172 21468 16178 21480
rect 16482 21468 16488 21480
rect 16172 21440 16488 21468
rect 16172 21428 16178 21440
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 16684 21400 16712 21499
rect 17586 21496 17592 21548
rect 17644 21496 17650 21548
rect 17862 21496 17868 21548
rect 17920 21496 17926 21548
rect 18892 21545 18920 21576
rect 19306 21576 19932 21604
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21536 18567 21539
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 18555 21508 18797 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 16758 21428 16764 21480
rect 16816 21468 16822 21480
rect 16853 21471 16911 21477
rect 16853 21468 16865 21471
rect 16816 21440 16865 21468
rect 16816 21428 16822 21440
rect 16853 21437 16865 21440
rect 16899 21468 16911 21471
rect 17034 21468 17040 21480
rect 16899 21440 17040 21468
rect 16899 21437 16911 21440
rect 16853 21431 16911 21437
rect 17034 21428 17040 21440
rect 17092 21428 17098 21480
rect 17678 21428 17684 21480
rect 17736 21477 17742 21480
rect 17736 21471 17764 21477
rect 17752 21437 17764 21471
rect 17736 21431 17764 21437
rect 17736 21428 17742 21431
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 19306 21468 19334 21576
rect 19518 21496 19524 21548
rect 19576 21496 19582 21548
rect 19794 21496 19800 21548
rect 19852 21496 19858 21548
rect 19904 21536 19932 21576
rect 20131 21539 20189 21545
rect 20131 21536 20143 21539
rect 19904 21508 20143 21536
rect 20131 21505 20143 21508
rect 20177 21505 20189 21539
rect 20916 21536 20944 21635
rect 20990 21632 20996 21684
rect 21048 21632 21054 21684
rect 21542 21632 21548 21684
rect 21600 21672 21606 21684
rect 22005 21675 22063 21681
rect 22005 21672 22017 21675
rect 21600 21644 22017 21672
rect 21600 21632 21606 21644
rect 22005 21641 22017 21644
rect 22051 21641 22063 21675
rect 22005 21635 22063 21641
rect 22278 21632 22284 21684
rect 22336 21672 22342 21684
rect 24397 21675 24455 21681
rect 22336 21644 24164 21672
rect 22336 21632 22342 21644
rect 21008 21604 21036 21632
rect 24136 21613 24164 21644
rect 24397 21641 24409 21675
rect 24443 21672 24455 21675
rect 24486 21672 24492 21684
rect 24443 21644 24492 21672
rect 24443 21641 24455 21644
rect 24397 21635 24455 21641
rect 24486 21632 24492 21644
rect 24544 21632 24550 21684
rect 24121 21607 24179 21613
rect 21008 21576 21404 21604
rect 21269 21539 21327 21545
rect 21269 21536 21281 21539
rect 20916 21508 21281 21536
rect 20131 21499 20189 21505
rect 21269 21505 21281 21508
rect 21315 21505 21327 21539
rect 21269 21499 21327 21505
rect 18104 21440 19334 21468
rect 19536 21468 19564 21496
rect 19889 21471 19947 21477
rect 19889 21468 19901 21471
rect 19536 21440 19901 21468
rect 18104 21428 18110 21440
rect 19889 21437 19901 21440
rect 19935 21437 19947 21471
rect 21376 21468 21404 21576
rect 24121 21573 24133 21607
rect 24167 21573 24179 21607
rect 24121 21567 24179 21573
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21508 21508 21833 21536
rect 21508 21496 21514 21508
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 21821 21499 21879 21505
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21536 23443 21539
rect 23474 21536 23480 21548
rect 23431 21508 23480 21536
rect 23431 21505 23443 21508
rect 23385 21499 23443 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 23569 21539 23627 21545
rect 23569 21505 23581 21539
rect 23615 21505 23627 21539
rect 23569 21499 23627 21505
rect 21545 21471 21603 21477
rect 21545 21468 21557 21471
rect 21376 21440 21557 21468
rect 19889 21431 19947 21437
rect 21545 21437 21557 21440
rect 21591 21437 21603 21471
rect 21545 21431 21603 21437
rect 23106 21428 23112 21480
rect 23164 21468 23170 21480
rect 23584 21468 23612 21499
rect 23658 21496 23664 21548
rect 23716 21496 23722 21548
rect 23164 21440 23612 21468
rect 23164 21428 23170 21440
rect 17126 21400 17132 21412
rect 16040 21372 16620 21400
rect 16684 21372 17132 21400
rect 14424 21304 14688 21332
rect 14424 21292 14430 21304
rect 15010 21292 15016 21344
rect 15068 21292 15074 21344
rect 15102 21292 15108 21344
rect 15160 21332 15166 21344
rect 16040 21332 16068 21372
rect 15160 21304 16068 21332
rect 15160 21292 15166 21304
rect 16114 21292 16120 21344
rect 16172 21292 16178 21344
rect 16592 21332 16620 21372
rect 17126 21360 17132 21372
rect 17184 21360 17190 21412
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 17313 21403 17371 21409
rect 17313 21400 17325 21403
rect 17276 21372 17325 21400
rect 17276 21360 17282 21372
rect 17313 21369 17325 21372
rect 17359 21369 17371 21403
rect 17313 21363 17371 21369
rect 18601 21403 18659 21409
rect 18601 21369 18613 21403
rect 18647 21400 18659 21403
rect 19334 21400 19340 21412
rect 18647 21372 19340 21400
rect 18647 21369 18659 21372
rect 18601 21363 18659 21369
rect 19334 21360 19340 21372
rect 19392 21360 19398 21412
rect 21453 21403 21511 21409
rect 21453 21369 21465 21403
rect 21499 21400 21511 21403
rect 23658 21400 23664 21412
rect 21499 21372 23664 21400
rect 21499 21369 21511 21372
rect 21453 21363 21511 21369
rect 23658 21360 23664 21372
rect 23716 21360 23722 21412
rect 17586 21332 17592 21344
rect 16592 21304 17592 21332
rect 17586 21292 17592 21304
rect 17644 21292 17650 21344
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 18969 21335 19027 21341
rect 18969 21332 18981 21335
rect 18840 21304 18981 21332
rect 18840 21292 18846 21304
rect 18969 21301 18981 21304
rect 19015 21301 19027 21335
rect 18969 21295 19027 21301
rect 19610 21292 19616 21344
rect 19668 21292 19674 21344
rect 21358 21292 21364 21344
rect 21416 21292 21422 21344
rect 23474 21292 23480 21344
rect 23532 21292 23538 21344
rect 23842 21292 23848 21344
rect 23900 21292 23906 21344
rect 1104 21242 24840 21264
rect 1104 21190 3917 21242
rect 3969 21190 3981 21242
rect 4033 21190 4045 21242
rect 4097 21190 4109 21242
rect 4161 21190 4173 21242
rect 4225 21190 9851 21242
rect 9903 21190 9915 21242
rect 9967 21190 9979 21242
rect 10031 21190 10043 21242
rect 10095 21190 10107 21242
rect 10159 21190 15785 21242
rect 15837 21190 15849 21242
rect 15901 21190 15913 21242
rect 15965 21190 15977 21242
rect 16029 21190 16041 21242
rect 16093 21190 21719 21242
rect 21771 21190 21783 21242
rect 21835 21190 21847 21242
rect 21899 21190 21911 21242
rect 21963 21190 21975 21242
rect 22027 21190 24840 21242
rect 1104 21168 24840 21190
rect 1394 21088 1400 21140
rect 1452 21088 1458 21140
rect 2501 21131 2559 21137
rect 2501 21097 2513 21131
rect 2547 21128 2559 21131
rect 8386 21128 8392 21140
rect 2547 21100 8392 21128
rect 2547 21097 2559 21100
rect 2501 21091 2559 21097
rect 8386 21088 8392 21100
rect 8444 21088 8450 21140
rect 8478 21088 8484 21140
rect 8536 21088 8542 21140
rect 8846 21088 8852 21140
rect 8904 21128 8910 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 8904 21100 9965 21128
rect 8904 21088 8910 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 14826 21128 14832 21140
rect 9953 21091 10011 21097
rect 10258 21100 14832 21128
rect 1412 21060 1440 21088
rect 2777 21063 2835 21069
rect 1412 21032 2728 21060
rect 1210 20952 1216 21004
rect 1268 20992 1274 21004
rect 1268 20964 2360 20992
rect 1268 20952 1274 20964
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 1673 20927 1731 20933
rect 1673 20893 1685 20927
rect 1719 20924 1731 20927
rect 2130 20924 2136 20936
rect 1719 20896 2136 20924
rect 1719 20893 1731 20896
rect 1673 20887 1731 20893
rect 2130 20884 2136 20896
rect 2188 20884 2194 20936
rect 2332 20933 2360 20964
rect 2317 20927 2375 20933
rect 2317 20893 2329 20927
rect 2363 20893 2375 20927
rect 2317 20887 2375 20893
rect 2593 20927 2651 20933
rect 2593 20893 2605 20927
rect 2639 20893 2651 20927
rect 2593 20887 2651 20893
rect 1302 20816 1308 20868
rect 1360 20856 1366 20868
rect 2608 20856 2636 20887
rect 1360 20828 2636 20856
rect 2700 20856 2728 21032
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 2866 21060 2872 21072
rect 2823 21032 2872 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 2866 21020 2872 21032
rect 2924 21020 2930 21072
rect 4706 21020 4712 21072
rect 4764 21020 4770 21072
rect 8202 21020 8208 21072
rect 8260 21060 8266 21072
rect 8260 21032 8892 21060
rect 8260 21020 8266 21032
rect 4724 20992 4752 21020
rect 8864 21004 8892 21032
rect 5902 20992 5908 21004
rect 4724 20964 5908 20992
rect 5902 20952 5908 20964
rect 5960 20952 5966 21004
rect 8478 20952 8484 21004
rect 8536 20992 8542 21004
rect 8662 20992 8668 21004
rect 8536 20964 8668 20992
rect 8536 20952 8542 20964
rect 8662 20952 8668 20964
rect 8720 20952 8726 21004
rect 8846 20952 8852 21004
rect 8904 20952 8910 21004
rect 2774 20884 2780 20936
rect 2832 20924 2838 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 2832 20896 3801 20924
rect 2832 20884 2838 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4063 20927 4121 20933
rect 4063 20893 4075 20927
rect 4109 20924 4121 20927
rect 4154 20924 4160 20936
rect 4109 20896 4160 20924
rect 4109 20893 4121 20896
rect 4063 20887 4121 20893
rect 4154 20884 4160 20896
rect 4212 20884 4218 20936
rect 4430 20884 4436 20936
rect 4488 20924 4494 20936
rect 5258 20924 5264 20936
rect 4488 20896 5264 20924
rect 4488 20884 4494 20896
rect 5258 20884 5264 20896
rect 5316 20884 5322 20936
rect 7469 20927 7527 20933
rect 7469 20893 7481 20927
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 7711 20927 7769 20933
rect 7711 20893 7723 20927
rect 7757 20924 7769 20927
rect 7834 20924 7840 20936
rect 7757 20896 7840 20924
rect 7757 20893 7769 20896
rect 7711 20887 7769 20893
rect 7484 20856 7512 20887
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8312 20896 8953 20924
rect 8312 20868 8340 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 9183 20927 9241 20933
rect 9183 20924 9195 20927
rect 8941 20887 8999 20893
rect 9048 20896 9195 20924
rect 8294 20856 8300 20868
rect 2700 20828 8300 20856
rect 1360 20816 1366 20828
rect 8294 20816 8300 20828
rect 8352 20816 8358 20868
rect 9048 20856 9076 20896
rect 9183 20893 9195 20896
rect 9229 20893 9241 20927
rect 9183 20887 9241 20893
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 10258 20924 10286 21100
rect 14826 21088 14832 21100
rect 14884 21088 14890 21140
rect 15010 21088 15016 21140
rect 15068 21088 15074 21140
rect 15378 21088 15384 21140
rect 15436 21128 15442 21140
rect 15436 21100 17632 21128
rect 15436 21088 15442 21100
rect 15028 21060 15056 21088
rect 17604 21060 17632 21100
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 17957 21131 18015 21137
rect 17957 21128 17969 21131
rect 17920 21100 17969 21128
rect 17920 21088 17926 21100
rect 17957 21097 17969 21100
rect 18003 21097 18015 21131
rect 17957 21091 18015 21097
rect 19610 21088 19616 21140
rect 19668 21088 19674 21140
rect 20441 21131 20499 21137
rect 20441 21097 20453 21131
rect 20487 21128 20499 21131
rect 21358 21128 21364 21140
rect 20487 21100 21364 21128
rect 20487 21097 20499 21100
rect 20441 21091 20499 21097
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 24210 21128 24216 21140
rect 22066 21100 24216 21128
rect 15028 21032 15516 21060
rect 17604 21032 19564 21060
rect 10318 20952 10324 21004
rect 10376 20952 10382 21004
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 13412 20964 14749 20992
rect 13412 20952 13418 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 14737 20955 14795 20961
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 15488 20992 15516 21032
rect 15657 20995 15715 21001
rect 15657 20992 15669 20995
rect 15488 20964 15669 20992
rect 15657 20961 15669 20964
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 15933 20995 15991 21001
rect 15933 20961 15945 20995
rect 15979 20992 15991 20995
rect 16114 20992 16120 21004
rect 15979 20964 16120 20992
rect 15979 20961 15991 20964
rect 15933 20955 15991 20961
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 16298 20952 16304 21004
rect 16356 20992 16362 21004
rect 16482 20992 16488 21004
rect 16356 20964 16488 20992
rect 16356 20952 16362 20964
rect 16482 20952 16488 20964
rect 16540 20992 16546 21004
rect 16945 20995 17003 21001
rect 16945 20992 16957 20995
rect 16540 20964 16957 20992
rect 16540 20952 16546 20964
rect 16945 20961 16957 20964
rect 16991 20961 17003 20995
rect 18782 20992 18788 21004
rect 16945 20955 17003 20961
rect 18708 20964 18788 20992
rect 10594 20933 10600 20936
rect 9640 20896 10286 20924
rect 10563 20927 10600 20933
rect 9640 20884 9646 20896
rect 10563 20893 10575 20927
rect 10563 20887 10600 20893
rect 10594 20884 10600 20887
rect 10652 20884 10658 20936
rect 11698 20884 11704 20936
rect 11756 20884 11762 20936
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 11974 20924 11980 20936
rect 11848 20896 11980 20924
rect 11848 20884 11854 20896
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12219 20927 12277 20933
rect 12219 20924 12231 20927
rect 12084 20896 12231 20924
rect 8588 20828 9076 20856
rect 1946 20748 1952 20800
rect 2004 20788 2010 20800
rect 2958 20788 2964 20800
rect 2004 20760 2964 20788
rect 2004 20748 2010 20760
rect 2958 20748 2964 20760
rect 3016 20748 3022 20800
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 4801 20791 4859 20797
rect 4801 20788 4813 20791
rect 4120 20760 4813 20788
rect 4120 20748 4126 20760
rect 4801 20757 4813 20760
rect 4847 20757 4859 20791
rect 4801 20751 4859 20757
rect 5074 20748 5080 20800
rect 5132 20788 5138 20800
rect 7650 20788 7656 20800
rect 5132 20760 7656 20788
rect 5132 20748 5138 20760
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 8110 20748 8116 20800
rect 8168 20788 8174 20800
rect 8588 20788 8616 20828
rect 9398 20816 9404 20868
rect 9456 20816 9462 20868
rect 11716 20856 11744 20884
rect 12084 20856 12112 20896
rect 12219 20893 12231 20896
rect 12265 20924 12277 20927
rect 12342 20924 12348 20936
rect 12265 20896 12348 20924
rect 12265 20893 12277 20896
rect 12219 20887 12277 20893
rect 12342 20884 12348 20896
rect 12400 20884 12406 20936
rect 13262 20884 13268 20936
rect 13320 20924 13326 20936
rect 14921 20927 14979 20933
rect 14921 20924 14933 20927
rect 13320 20896 14933 20924
rect 13320 20884 13326 20896
rect 14921 20893 14933 20896
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 15746 20884 15752 20936
rect 15804 20933 15810 20936
rect 18708 20933 18736 20964
rect 18782 20952 18788 20964
rect 18840 20952 18846 21004
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20992 18935 20995
rect 18923 20964 19012 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 15804 20927 15832 20933
rect 15820 20893 15832 20927
rect 17187 20927 17245 20933
rect 17187 20924 17199 20927
rect 15804 20887 15832 20893
rect 17052 20896 17199 20924
rect 15804 20884 15810 20887
rect 11716 20828 12112 20856
rect 16666 20816 16672 20868
rect 16724 20856 16730 20868
rect 17052 20856 17080 20896
rect 17187 20893 17199 20896
rect 17233 20893 17245 20927
rect 17187 20887 17245 20893
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20893 18751 20927
rect 18984 20924 19012 20964
rect 19334 20952 19340 21004
rect 19392 20992 19398 21004
rect 19392 20964 19472 20992
rect 19392 20952 19398 20964
rect 19150 20924 19156 20936
rect 18984 20896 19156 20924
rect 18693 20887 18751 20893
rect 19150 20884 19156 20896
rect 19208 20924 19214 20936
rect 19444 20933 19472 20964
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 19208 20896 19257 20924
rect 19208 20884 19214 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 16724 20828 17080 20856
rect 18969 20859 19027 20865
rect 16724 20816 16730 20828
rect 18969 20825 18981 20859
rect 19015 20825 19027 20859
rect 18969 20819 19027 20825
rect 19061 20859 19119 20865
rect 19061 20825 19073 20859
rect 19107 20856 19119 20859
rect 19337 20859 19395 20865
rect 19337 20856 19349 20859
rect 19107 20828 19349 20856
rect 19107 20825 19119 20828
rect 19061 20819 19119 20825
rect 19337 20825 19349 20828
rect 19383 20825 19395 20859
rect 19536 20856 19564 21032
rect 19628 20924 19656 21088
rect 20714 21020 20720 21072
rect 20772 21020 20778 21072
rect 20254 20952 20260 21004
rect 20312 20992 20318 21004
rect 22066 20992 22094 21100
rect 24210 21088 24216 21100
rect 24268 21088 24274 21140
rect 20312 20964 22094 20992
rect 20312 20952 20318 20964
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 22557 20995 22615 21001
rect 22557 20992 22569 20995
rect 22428 20964 22569 20992
rect 22428 20952 22434 20964
rect 22557 20961 22569 20964
rect 22603 20961 22615 20995
rect 22557 20955 22615 20961
rect 20349 20927 20407 20933
rect 20349 20924 20361 20927
rect 19628 20896 20361 20924
rect 20349 20893 20361 20896
rect 20395 20893 20407 20927
rect 20349 20887 20407 20893
rect 20898 20884 20904 20936
rect 20956 20884 20962 20936
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22813 20927 22871 20933
rect 22813 20924 22825 20927
rect 22152 20896 22825 20924
rect 22152 20884 22158 20896
rect 22813 20893 22825 20896
rect 22859 20893 22871 20927
rect 22813 20887 22871 20893
rect 24026 20884 24032 20936
rect 24084 20884 24090 20936
rect 22646 20856 22652 20868
rect 19536 20828 22652 20856
rect 19337 20819 19395 20825
rect 8168 20760 8616 20788
rect 8168 20748 8174 20760
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 9416 20788 9444 20816
rect 8720 20760 9444 20788
rect 8720 20748 8726 20760
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11333 20791 11391 20797
rect 11333 20788 11345 20791
rect 11020 20760 11345 20788
rect 11020 20748 11026 20760
rect 11333 20757 11345 20760
rect 11379 20757 11391 20791
rect 11333 20751 11391 20757
rect 12710 20748 12716 20800
rect 12768 20788 12774 20800
rect 12989 20791 13047 20797
rect 12989 20788 13001 20791
rect 12768 20760 13001 20788
rect 12768 20748 12774 20760
rect 12989 20757 13001 20760
rect 13035 20757 13047 20791
rect 12989 20751 13047 20757
rect 14458 20748 14464 20800
rect 14516 20788 14522 20800
rect 15746 20788 15752 20800
rect 14516 20760 15752 20788
rect 14516 20748 14522 20760
rect 15746 20748 15752 20760
rect 15804 20748 15810 20800
rect 16574 20748 16580 20800
rect 16632 20748 16638 20800
rect 18984 20788 19012 20819
rect 22646 20816 22652 20828
rect 22704 20816 22710 20868
rect 19702 20788 19708 20800
rect 18984 20760 19708 20788
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 23290 20748 23296 20800
rect 23348 20788 23354 20800
rect 23937 20791 23995 20797
rect 23937 20788 23949 20791
rect 23348 20760 23949 20788
rect 23348 20748 23354 20760
rect 23937 20757 23949 20760
rect 23983 20757 23995 20791
rect 23937 20751 23995 20757
rect 24121 20791 24179 20797
rect 24121 20757 24133 20791
rect 24167 20788 24179 20791
rect 24210 20788 24216 20800
rect 24167 20760 24216 20788
rect 24167 20757 24179 20760
rect 24121 20751 24179 20757
rect 24210 20748 24216 20760
rect 24268 20748 24274 20800
rect 1104 20698 25000 20720
rect 1104 20646 6884 20698
rect 6936 20646 6948 20698
rect 7000 20646 7012 20698
rect 7064 20646 7076 20698
rect 7128 20646 7140 20698
rect 7192 20646 12818 20698
rect 12870 20646 12882 20698
rect 12934 20646 12946 20698
rect 12998 20646 13010 20698
rect 13062 20646 13074 20698
rect 13126 20646 18752 20698
rect 18804 20646 18816 20698
rect 18868 20646 18880 20698
rect 18932 20646 18944 20698
rect 18996 20646 19008 20698
rect 19060 20646 24686 20698
rect 24738 20646 24750 20698
rect 24802 20646 24814 20698
rect 24866 20646 24878 20698
rect 24930 20646 24942 20698
rect 24994 20646 25000 20698
rect 1104 20624 25000 20646
rect 3786 20544 3792 20596
rect 3844 20584 3850 20596
rect 7834 20584 7840 20596
rect 3844 20556 7840 20584
rect 3844 20544 3850 20556
rect 7834 20544 7840 20556
rect 7892 20544 7898 20596
rect 8846 20544 8852 20596
rect 8904 20584 8910 20596
rect 9214 20584 9220 20596
rect 8904 20556 9220 20584
rect 8904 20544 8910 20556
rect 9214 20544 9220 20556
rect 9272 20544 9278 20596
rect 10410 20584 10416 20596
rect 9876 20556 10416 20584
rect 5258 20516 5264 20528
rect 4816 20488 5264 20516
rect 1671 20451 1729 20457
rect 1671 20417 1683 20451
rect 1717 20448 1729 20451
rect 2590 20448 2596 20460
rect 1717 20420 2596 20448
rect 1717 20417 1729 20420
rect 1671 20411 1729 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 3878 20408 3884 20460
rect 3936 20457 3942 20460
rect 3936 20451 3964 20457
rect 3952 20417 3964 20451
rect 3936 20411 3964 20417
rect 3936 20408 3942 20411
rect 4062 20408 4068 20460
rect 4120 20408 4126 20460
rect 4816 20457 4844 20488
rect 5258 20476 5264 20488
rect 5316 20516 5322 20528
rect 5316 20488 6592 20516
rect 5316 20476 5322 20488
rect 6564 20460 6592 20488
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 5075 20451 5133 20457
rect 5075 20417 5087 20451
rect 5121 20448 5133 20451
rect 5121 20420 6500 20448
rect 5121 20417 5133 20420
rect 5075 20411 5133 20417
rect 1394 20340 1400 20392
rect 1452 20340 1458 20392
rect 2869 20383 2927 20389
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 2958 20380 2964 20392
rect 2915 20352 2964 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 3053 20383 3111 20389
rect 3053 20349 3065 20383
rect 3099 20349 3111 20383
rect 3053 20343 3111 20349
rect 3789 20383 3847 20389
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 4246 20380 4252 20392
rect 3835 20352 4252 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 3068 20312 3096 20343
rect 4246 20340 4252 20352
rect 4304 20340 4310 20392
rect 6472 20380 6500 20420
rect 6546 20408 6552 20460
rect 6604 20408 6610 20460
rect 9876 20448 9904 20556
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 11238 20584 11244 20596
rect 10704 20556 11244 20584
rect 9953 20519 10011 20525
rect 9953 20485 9965 20519
rect 9999 20516 10011 20519
rect 10502 20516 10508 20528
rect 9999 20488 10508 20516
rect 9999 20485 10011 20488
rect 9953 20479 10011 20485
rect 10502 20476 10508 20488
rect 10560 20476 10566 20528
rect 10704 20525 10732 20556
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 13262 20584 13268 20596
rect 12360 20556 13268 20584
rect 10689 20519 10747 20525
rect 10689 20485 10701 20519
rect 10735 20485 10747 20519
rect 10689 20479 10747 20485
rect 11057 20519 11115 20525
rect 11057 20485 11069 20519
rect 11103 20516 11115 20519
rect 11330 20516 11336 20528
rect 11103 20488 11336 20516
rect 11103 20485 11115 20488
rect 11057 20479 11115 20485
rect 11330 20476 11336 20488
rect 11388 20516 11394 20528
rect 11388 20488 11560 20516
rect 11388 20476 11394 20488
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9876 20420 10241 20448
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10321 20451 10379 20457
rect 10321 20417 10333 20451
rect 10367 20448 10379 20451
rect 10594 20448 10600 20460
rect 10367 20420 10600 20448
rect 10367 20417 10379 20420
rect 10321 20411 10379 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 11422 20408 11428 20460
rect 11480 20408 11486 20460
rect 10968 20392 11020 20398
rect 8662 20380 8668 20392
rect 6472 20352 8668 20380
rect 8662 20340 8668 20352
rect 8720 20340 8726 20392
rect 10968 20334 11020 20340
rect 2332 20284 3096 20312
rect 1854 20204 1860 20256
rect 1912 20244 1918 20256
rect 2332 20244 2360 20284
rect 3510 20272 3516 20324
rect 3568 20272 3574 20324
rect 11440 20312 11468 20408
rect 11532 20380 11560 20488
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 12360 20457 12388 20556
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 15378 20544 15384 20596
rect 15436 20544 15442 20596
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 16206 20584 16212 20596
rect 15528 20556 16212 20584
rect 15528 20544 15534 20556
rect 16206 20544 16212 20556
rect 16264 20584 16270 20596
rect 18046 20584 18052 20596
rect 16264 20556 18052 20584
rect 16264 20544 16270 20556
rect 18046 20544 18052 20556
rect 18104 20544 18110 20596
rect 18785 20587 18843 20593
rect 18785 20553 18797 20587
rect 18831 20584 18843 20587
rect 19150 20584 19156 20596
rect 18831 20556 19156 20584
rect 18831 20553 18843 20556
rect 18785 20547 18843 20553
rect 19150 20544 19156 20556
rect 19208 20544 19214 20596
rect 22094 20544 22100 20596
rect 22152 20544 22158 20596
rect 23566 20544 23572 20596
rect 23624 20584 23630 20596
rect 23753 20587 23811 20593
rect 23753 20584 23765 20587
rect 23624 20556 23765 20584
rect 23624 20544 23630 20556
rect 23753 20553 23765 20556
rect 23799 20553 23811 20587
rect 23753 20547 23811 20553
rect 14734 20476 14740 20528
rect 14792 20516 14798 20528
rect 19610 20516 19616 20528
rect 14792 20488 19616 20516
rect 14792 20476 14798 20488
rect 19610 20476 19616 20488
rect 19668 20476 19674 20528
rect 22112 20516 22140 20544
rect 22112 20488 22692 20516
rect 12345 20451 12403 20457
rect 12345 20448 12357 20451
rect 11756 20420 12357 20448
rect 11756 20408 11762 20420
rect 12345 20417 12357 20420
rect 12391 20417 12403 20451
rect 12345 20411 12403 20417
rect 13354 20408 13360 20460
rect 13412 20457 13418 20460
rect 13412 20451 13440 20457
rect 13428 20417 13440 20451
rect 13412 20411 13440 20417
rect 13412 20408 13418 20411
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 14366 20408 14372 20460
rect 14424 20408 14430 20460
rect 14642 20457 14648 20460
rect 14611 20451 14648 20457
rect 14611 20417 14623 20451
rect 14611 20411 14648 20417
rect 14642 20408 14648 20411
rect 14700 20408 14706 20460
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 16356 20420 17785 20448
rect 16356 20408 16362 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18047 20451 18105 20457
rect 18047 20448 18059 20451
rect 18012 20420 18059 20448
rect 18012 20408 18018 20420
rect 18047 20417 18059 20420
rect 18093 20417 18105 20451
rect 18047 20411 18105 20417
rect 18506 20408 18512 20460
rect 18564 20448 18570 20460
rect 19150 20448 19156 20460
rect 18564 20420 19156 20448
rect 18564 20408 18570 20420
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22373 20451 22431 20457
rect 22373 20448 22385 20451
rect 22152 20420 22385 20448
rect 22152 20408 22158 20420
rect 22373 20417 22385 20420
rect 22419 20417 22431 20451
rect 22373 20411 22431 20417
rect 22554 20408 22560 20460
rect 22612 20408 22618 20460
rect 22664 20457 22692 20488
rect 22830 20476 22836 20528
rect 22888 20516 22894 20528
rect 22888 20488 22968 20516
rect 22888 20476 22894 20488
rect 22940 20478 22968 20488
rect 22999 20481 23057 20487
rect 22999 20478 23011 20481
rect 22649 20451 22707 20457
rect 22649 20417 22661 20451
rect 22695 20417 22707 20451
rect 22940 20450 23011 20478
rect 22999 20447 23011 20450
rect 23045 20447 23057 20481
rect 22999 20441 23057 20447
rect 23768 20448 23796 20547
rect 24121 20451 24179 20457
rect 24121 20448 24133 20451
rect 23768 20420 24133 20448
rect 22649 20411 22707 20417
rect 24121 20417 24133 20420
rect 24167 20417 24179 20451
rect 24121 20411 24179 20417
rect 24210 20408 24216 20460
rect 24268 20408 24274 20460
rect 12529 20383 12587 20389
rect 12529 20380 12541 20383
rect 11532 20352 12541 20380
rect 12529 20349 12541 20352
rect 12575 20380 12587 20383
rect 12618 20380 12624 20392
rect 12575 20352 12624 20380
rect 12575 20349 12587 20352
rect 12529 20343 12587 20349
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 12989 20383 13047 20389
rect 12989 20380 13001 20383
rect 12768 20352 13001 20380
rect 12768 20340 12774 20352
rect 12989 20349 13001 20352
rect 13035 20349 13047 20383
rect 13265 20383 13323 20389
rect 13265 20380 13277 20383
rect 12989 20343 13047 20349
rect 13096 20352 13277 20380
rect 13096 20312 13124 20352
rect 13265 20349 13277 20352
rect 13311 20380 13323 20383
rect 13311 20352 14412 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 11440 20284 13124 20312
rect 1912 20216 2360 20244
rect 1912 20204 1918 20216
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 4706 20204 4712 20256
rect 4764 20204 4770 20256
rect 5810 20204 5816 20256
rect 5868 20204 5874 20256
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 9398 20244 9404 20256
rect 6696 20216 9404 20244
rect 6696 20204 6702 20216
rect 9398 20204 9404 20216
rect 9456 20204 9462 20256
rect 11238 20204 11244 20256
rect 11296 20204 11302 20256
rect 14182 20204 14188 20256
rect 14240 20204 14246 20256
rect 14384 20244 14412 20352
rect 15378 20340 15384 20392
rect 15436 20380 15442 20392
rect 15746 20380 15752 20392
rect 15436 20352 15752 20380
rect 15436 20340 15442 20352
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 22572 20380 22600 20408
rect 22741 20383 22799 20389
rect 22741 20380 22753 20383
rect 22572 20352 22753 20380
rect 22741 20349 22753 20352
rect 22787 20349 22799 20383
rect 22741 20343 22799 20349
rect 23474 20340 23480 20392
rect 23532 20380 23538 20392
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 23532 20352 24409 20380
rect 23532 20340 23538 20352
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17678 20312 17684 20324
rect 17000 20284 17684 20312
rect 17000 20272 17006 20284
rect 17678 20272 17684 20284
rect 17736 20272 17742 20324
rect 22189 20315 22247 20321
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 22646 20312 22652 20324
rect 22235 20284 22652 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 22646 20272 22652 20284
rect 22704 20272 22710 20324
rect 24026 20312 24032 20324
rect 23400 20284 24032 20312
rect 16114 20244 16120 20256
rect 14384 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20244 16178 20256
rect 16666 20244 16672 20256
rect 16172 20216 16672 20244
rect 16172 20204 16178 20216
rect 16666 20204 16672 20216
rect 16724 20204 16730 20256
rect 22465 20247 22523 20253
rect 22465 20213 22477 20247
rect 22511 20244 22523 20247
rect 23400 20244 23428 20284
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 22511 20216 23428 20244
rect 22511 20213 22523 20216
rect 22465 20207 22523 20213
rect 24210 20204 24216 20256
rect 24268 20244 24274 20256
rect 24305 20247 24363 20253
rect 24305 20244 24317 20247
rect 24268 20216 24317 20244
rect 24268 20204 24274 20216
rect 24305 20213 24317 20216
rect 24351 20213 24363 20247
rect 24305 20207 24363 20213
rect 1104 20154 24840 20176
rect 1104 20102 3917 20154
rect 3969 20102 3981 20154
rect 4033 20102 4045 20154
rect 4097 20102 4109 20154
rect 4161 20102 4173 20154
rect 4225 20102 9851 20154
rect 9903 20102 9915 20154
rect 9967 20102 9979 20154
rect 10031 20102 10043 20154
rect 10095 20102 10107 20154
rect 10159 20102 15785 20154
rect 15837 20102 15849 20154
rect 15901 20102 15913 20154
rect 15965 20102 15977 20154
rect 16029 20102 16041 20154
rect 16093 20102 21719 20154
rect 21771 20102 21783 20154
rect 21835 20102 21847 20154
rect 21899 20102 21911 20154
rect 21963 20102 21975 20154
rect 22027 20102 24840 20154
rect 1104 20080 24840 20102
rect 1578 20000 1584 20052
rect 1636 20000 1642 20052
rect 2774 20040 2780 20052
rect 2332 20012 2780 20040
rect 2222 19864 2228 19916
rect 2280 19904 2286 19916
rect 2332 19913 2360 20012
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 3329 20043 3387 20049
rect 3329 20009 3341 20043
rect 3375 20040 3387 20043
rect 3510 20040 3516 20052
rect 3375 20012 3516 20040
rect 3375 20009 3387 20012
rect 3329 20003 3387 20009
rect 3510 20000 3516 20012
rect 3568 20000 3574 20052
rect 3973 20043 4031 20049
rect 3973 20009 3985 20043
rect 4019 20040 4031 20043
rect 5166 20040 5172 20052
rect 4019 20012 5172 20040
rect 4019 20009 4031 20012
rect 3973 20003 4031 20009
rect 5166 20000 5172 20012
rect 5224 20000 5230 20052
rect 7653 20043 7711 20049
rect 7653 20009 7665 20043
rect 7699 20009 7711 20043
rect 7653 20003 7711 20009
rect 7668 19916 7696 20003
rect 10594 20000 10600 20052
rect 10652 20040 10658 20052
rect 11149 20043 11207 20049
rect 11149 20040 11161 20043
rect 10652 20012 11161 20040
rect 10652 20000 10658 20012
rect 11149 20009 11161 20012
rect 11195 20009 11207 20043
rect 11149 20003 11207 20009
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 13354 20040 13360 20052
rect 12032 20012 13360 20040
rect 12032 20000 12038 20012
rect 2317 19907 2375 19913
rect 2317 19904 2329 19907
rect 2280 19876 2329 19904
rect 2280 19864 2286 19876
rect 2317 19873 2329 19876
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 5810 19864 5816 19916
rect 5868 19864 5874 19916
rect 6546 19864 6552 19916
rect 6604 19904 6610 19916
rect 6641 19907 6699 19913
rect 6641 19904 6653 19907
rect 6604 19876 6653 19904
rect 6604 19864 6610 19876
rect 6641 19873 6653 19876
rect 6687 19873 6699 19907
rect 6641 19867 6699 19873
rect 7650 19864 7656 19916
rect 7708 19864 7714 19916
rect 12544 19913 12572 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 13538 20000 13544 20052
rect 13596 20000 13602 20052
rect 13998 20000 14004 20052
rect 14056 20040 14062 20052
rect 16298 20040 16304 20052
rect 14056 20012 16304 20040
rect 14056 20000 14062 20012
rect 16298 20000 16304 20012
rect 16356 20000 16362 20052
rect 16574 20000 16580 20052
rect 16632 20040 16638 20052
rect 16632 20012 20760 20040
rect 16632 20000 16638 20012
rect 17770 19932 17776 19984
rect 17828 19932 17834 19984
rect 12529 19907 12587 19913
rect 12529 19873 12541 19907
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 14240 19876 15853 19904
rect 14240 19864 14246 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 16298 19864 16304 19916
rect 16356 19864 16362 19916
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16577 19907 16635 19913
rect 16577 19904 16589 19907
rect 16448 19876 16589 19904
rect 16448 19864 16454 19876
rect 16577 19873 16589 19876
rect 16623 19873 16635 19907
rect 17034 19904 17040 19916
rect 16577 19867 16635 19873
rect 16730 19876 17040 19904
rect 750 19796 756 19848
rect 808 19836 814 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 808 19808 1501 19836
rect 808 19796 814 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 2590 19836 2596 19848
rect 2551 19808 2596 19836
rect 1489 19799 1547 19805
rect 2590 19796 2596 19808
rect 2648 19796 2654 19848
rect 3789 19839 3847 19845
rect 3789 19836 3801 19839
rect 2746 19808 3801 19836
rect 1302 19728 1308 19780
rect 1360 19768 1366 19780
rect 2746 19768 2774 19808
rect 3789 19805 3801 19808
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 4893 19839 4951 19845
rect 4893 19805 4905 19839
rect 4939 19836 4951 19839
rect 4939 19808 5304 19836
rect 4939 19805 4951 19808
rect 4893 19799 4951 19805
rect 1360 19740 2774 19768
rect 1360 19728 1366 19740
rect 4430 19728 4436 19780
rect 4488 19768 4494 19780
rect 5123 19771 5181 19777
rect 5123 19768 5135 19771
rect 4488 19740 5135 19768
rect 4488 19728 4494 19740
rect 5123 19737 5135 19740
rect 5169 19737 5181 19771
rect 5276 19768 5304 19808
rect 5350 19796 5356 19848
rect 5408 19836 5414 19848
rect 5408 19808 5672 19836
rect 5408 19796 5414 19808
rect 5445 19771 5503 19777
rect 5445 19768 5457 19771
rect 5276 19740 5457 19768
rect 5123 19731 5181 19737
rect 5445 19737 5457 19740
rect 5491 19737 5503 19771
rect 5445 19731 5503 19737
rect 5534 19728 5540 19780
rect 5592 19728 5598 19780
rect 5644 19768 5672 19808
rect 5902 19796 5908 19848
rect 5960 19796 5966 19848
rect 6915 19839 6973 19845
rect 6915 19805 6927 19839
rect 6961 19836 6973 19839
rect 8205 19839 8263 19845
rect 6961 19808 7328 19836
rect 6961 19805 6973 19808
rect 6915 19799 6973 19805
rect 6273 19771 6331 19777
rect 6273 19768 6285 19771
rect 5644 19740 6285 19768
rect 6273 19737 6285 19740
rect 6319 19737 6331 19771
rect 7300 19768 7328 19808
rect 8205 19805 8217 19839
rect 8251 19836 8263 19839
rect 8294 19836 8300 19848
rect 8251 19808 8300 19836
rect 8251 19805 8263 19808
rect 8205 19799 8263 19805
rect 8294 19796 8300 19808
rect 8352 19796 8358 19848
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 10042 19836 10048 19848
rect 8444 19808 10048 19836
rect 8444 19796 8450 19808
rect 10042 19796 10048 19808
rect 10100 19796 10106 19848
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 10318 19836 10324 19848
rect 10183 19808 10324 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 10411 19839 10469 19845
rect 10411 19805 10423 19839
rect 10457 19836 10469 19839
rect 10870 19836 10876 19848
rect 10457 19808 10876 19836
rect 10457 19805 10469 19808
rect 10411 19799 10469 19805
rect 10870 19796 10876 19808
rect 10928 19796 10934 19848
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11606 19836 11612 19848
rect 11296 19808 11612 19836
rect 11296 19796 11302 19808
rect 11606 19796 11612 19808
rect 11664 19796 11670 19848
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 12803 19839 12861 19845
rect 12803 19836 12815 19839
rect 12768 19808 12815 19836
rect 12768 19796 12774 19808
rect 12803 19805 12815 19808
rect 12849 19836 12861 19839
rect 13262 19836 13268 19848
rect 12849 19808 13268 19836
rect 12849 19805 12861 19808
rect 12803 19799 12861 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13446 19796 13452 19848
rect 13504 19836 13510 19848
rect 14642 19836 14648 19848
rect 13504 19808 14648 19836
rect 13504 19796 13510 19808
rect 14642 19796 14648 19808
rect 14700 19796 14706 19848
rect 16730 19845 16758 19876
rect 17034 19864 17040 19876
rect 17092 19864 17098 19916
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 16715 19839 16773 19845
rect 16715 19805 16727 19839
rect 16761 19805 16773 19839
rect 16715 19799 16773 19805
rect 7558 19768 7564 19780
rect 7300 19740 7564 19768
rect 6273 19731 6331 19737
rect 7558 19728 7564 19740
rect 7616 19728 7622 19780
rect 8938 19728 8944 19780
rect 8996 19768 9002 19780
rect 15102 19768 15108 19780
rect 8996 19740 15108 19768
rect 8996 19728 9002 19740
rect 15102 19728 15108 19740
rect 15160 19768 15166 19780
rect 15672 19768 15700 19799
rect 16850 19796 16856 19848
rect 16908 19796 16914 19848
rect 17788 19836 17816 19932
rect 20732 19904 20760 20012
rect 22094 20000 22100 20052
rect 22152 20000 22158 20052
rect 22554 20040 22560 20052
rect 22204 20012 22560 20040
rect 22204 19913 22232 20012
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 23937 20043 23995 20049
rect 23937 20009 23949 20043
rect 23983 20040 23995 20043
rect 24026 20040 24032 20052
rect 23983 20012 24032 20040
rect 23983 20009 23995 20012
rect 23937 20003 23995 20009
rect 24026 20000 24032 20012
rect 24084 20000 24090 20052
rect 22189 19907 22247 19913
rect 20732 19876 20852 19904
rect 19061 19839 19119 19845
rect 19061 19836 19073 19839
rect 17788 19808 19073 19836
rect 19061 19805 19073 19808
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 15160 19740 15700 19768
rect 19076 19768 19104 19799
rect 19242 19796 19248 19848
rect 19300 19836 19306 19848
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 19300 19808 20729 19836
rect 19300 19796 19306 19808
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 20824 19836 20852 19876
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 20973 19839 21031 19845
rect 20973 19836 20985 19839
rect 20824 19808 20985 19836
rect 20717 19799 20775 19805
rect 20973 19805 20985 19808
rect 21019 19836 21031 19839
rect 21266 19836 21272 19848
rect 21019 19808 21272 19836
rect 21019 19805 21031 19808
rect 20973 19799 21031 19805
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 21542 19796 21548 19848
rect 21600 19836 21606 19848
rect 22431 19839 22489 19845
rect 22431 19836 22443 19839
rect 21600 19808 22094 19836
rect 21600 19796 21606 19808
rect 19490 19771 19548 19777
rect 19490 19768 19502 19771
rect 19076 19740 19502 19768
rect 15160 19728 15166 19740
rect 19490 19737 19502 19740
rect 19536 19737 19548 19771
rect 22066 19768 22094 19808
rect 22296 19808 22443 19836
rect 22296 19768 22324 19808
rect 22431 19805 22443 19808
rect 22477 19805 22489 19839
rect 22431 19799 22489 19805
rect 23658 19796 23664 19848
rect 23716 19796 23722 19848
rect 23842 19768 23848 19780
rect 22066 19740 22324 19768
rect 23124 19740 23848 19768
rect 19490 19731 19548 19737
rect 6457 19703 6515 19709
rect 6457 19669 6469 19703
rect 6503 19700 6515 19703
rect 6730 19700 6736 19712
rect 6503 19672 6736 19700
rect 6503 19669 6515 19672
rect 6457 19663 6515 19669
rect 6730 19660 6736 19672
rect 6788 19660 6794 19712
rect 6822 19660 6828 19712
rect 6880 19700 6886 19712
rect 11698 19700 11704 19712
rect 6880 19672 11704 19700
rect 6880 19660 6886 19672
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 11974 19660 11980 19712
rect 12032 19700 12038 19712
rect 14274 19700 14280 19712
rect 12032 19672 14280 19700
rect 12032 19660 12038 19672
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 17310 19700 17316 19712
rect 16632 19672 17316 19700
rect 16632 19660 16638 19672
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 17954 19700 17960 19712
rect 17543 19672 17960 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 17954 19660 17960 19672
rect 18012 19660 18018 19712
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 18877 19703 18935 19709
rect 18877 19700 18889 19703
rect 18656 19672 18889 19700
rect 18656 19660 18662 19672
rect 18877 19669 18889 19672
rect 18923 19669 18935 19703
rect 18877 19663 18935 19669
rect 20622 19660 20628 19712
rect 20680 19660 20686 19712
rect 20806 19660 20812 19712
rect 20864 19700 20870 19712
rect 23124 19700 23152 19740
rect 23842 19728 23848 19740
rect 23900 19728 23906 19780
rect 20864 19672 23152 19700
rect 20864 19660 20870 19672
rect 23198 19660 23204 19712
rect 23256 19660 23262 19712
rect 1104 19610 25000 19632
rect 1104 19558 6884 19610
rect 6936 19558 6948 19610
rect 7000 19558 7012 19610
rect 7064 19558 7076 19610
rect 7128 19558 7140 19610
rect 7192 19558 12818 19610
rect 12870 19558 12882 19610
rect 12934 19558 12946 19610
rect 12998 19558 13010 19610
rect 13062 19558 13074 19610
rect 13126 19558 18752 19610
rect 18804 19558 18816 19610
rect 18868 19558 18880 19610
rect 18932 19558 18944 19610
rect 18996 19558 19008 19610
rect 19060 19558 24686 19610
rect 24738 19558 24750 19610
rect 24802 19558 24814 19610
rect 24866 19558 24878 19610
rect 24930 19558 24942 19610
rect 24994 19558 25000 19610
rect 1104 19536 25000 19558
rect 1578 19456 1584 19508
rect 1636 19456 1642 19508
rect 2038 19456 2044 19508
rect 2096 19496 2102 19508
rect 3053 19499 3111 19505
rect 3053 19496 3065 19499
rect 2096 19468 3065 19496
rect 2096 19456 2102 19468
rect 3053 19465 3065 19468
rect 3099 19465 3111 19499
rect 3053 19459 3111 19465
rect 3513 19499 3571 19505
rect 3513 19465 3525 19499
rect 3559 19496 3571 19499
rect 4614 19496 4620 19508
rect 3559 19468 4620 19496
rect 3559 19465 3571 19468
rect 3513 19459 3571 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 4706 19456 4712 19508
rect 4764 19456 4770 19508
rect 5258 19456 5264 19508
rect 5316 19456 5322 19508
rect 5534 19456 5540 19508
rect 5592 19496 5598 19508
rect 5905 19499 5963 19505
rect 5905 19496 5917 19499
rect 5592 19468 5917 19496
rect 5592 19456 5598 19468
rect 5905 19465 5917 19468
rect 5951 19465 5963 19499
rect 5905 19459 5963 19465
rect 6638 19456 6644 19508
rect 6696 19456 6702 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7466 19496 7472 19508
rect 7147 19468 7472 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7466 19456 7472 19468
rect 7524 19496 7530 19508
rect 7926 19496 7932 19508
rect 7524 19468 7932 19496
rect 7524 19456 7530 19468
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8294 19496 8300 19508
rect 8034 19468 8300 19496
rect 4724 19428 4752 19456
rect 5276 19428 5304 19456
rect 3252 19400 4752 19428
rect 4908 19400 5304 19428
rect 842 19320 848 19372
rect 900 19360 906 19372
rect 1397 19363 1455 19369
rect 1397 19360 1409 19363
rect 900 19332 1409 19360
rect 900 19320 906 19332
rect 1397 19329 1409 19332
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1947 19363 2005 19369
rect 1947 19329 1959 19363
rect 1993 19360 2005 19363
rect 2590 19360 2596 19372
rect 1993 19332 2596 19360
rect 1993 19329 2005 19332
rect 1947 19323 2005 19329
rect 2590 19320 2596 19332
rect 2648 19320 2654 19372
rect 3252 19369 3280 19400
rect 3237 19363 3295 19369
rect 3237 19329 3249 19363
rect 3283 19329 3295 19363
rect 3237 19323 3295 19329
rect 3326 19320 3332 19372
rect 3384 19320 3390 19372
rect 4908 19369 4936 19400
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 5167 19363 5225 19369
rect 5167 19329 5179 19363
rect 5213 19360 5225 19363
rect 6656 19360 6684 19456
rect 8034 19428 8062 19468
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 9122 19456 9128 19508
rect 9180 19496 9186 19508
rect 14182 19496 14188 19508
rect 9180 19468 14188 19496
rect 9180 19456 9186 19468
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14274 19456 14280 19508
rect 14332 19496 14338 19508
rect 14332 19468 16804 19496
rect 14332 19456 14338 19468
rect 7392 19400 8062 19428
rect 7392 19369 7420 19400
rect 8202 19388 8208 19440
rect 8260 19388 8266 19440
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 9766 19428 9772 19440
rect 8628 19400 9772 19428
rect 8628 19388 8634 19400
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 10042 19388 10048 19440
rect 10100 19428 10106 19440
rect 13998 19428 14004 19440
rect 10100 19400 14004 19428
rect 10100 19388 10106 19400
rect 5213 19332 6684 19360
rect 7377 19363 7435 19369
rect 5213 19329 5225 19332
rect 5167 19323 5225 19329
rect 7377 19329 7389 19363
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 7466 19320 7472 19372
rect 7524 19320 7530 19372
rect 7834 19360 7840 19372
rect 7795 19332 7840 19360
rect 7834 19320 7840 19332
rect 7892 19360 7898 19372
rect 8294 19360 8300 19372
rect 7892 19332 8300 19360
rect 7892 19320 7898 19332
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 8386 19320 8392 19372
rect 8444 19360 8450 19372
rect 8849 19363 8907 19369
rect 8849 19360 8861 19363
rect 8444 19332 8861 19360
rect 8444 19320 8450 19332
rect 8849 19329 8861 19332
rect 8895 19329 8907 19363
rect 8849 19323 8907 19329
rect 9123 19363 9181 19369
rect 9123 19329 9135 19363
rect 9169 19360 9181 19363
rect 10318 19360 10324 19372
rect 9169 19332 10324 19360
rect 9169 19329 9181 19332
rect 9123 19323 9181 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 11791 19363 11849 19369
rect 11791 19360 11803 19363
rect 11756 19332 11803 19360
rect 11756 19320 11762 19332
rect 11791 19329 11803 19332
rect 11837 19360 11849 19363
rect 12250 19360 12256 19372
rect 11837 19332 12256 19360
rect 11837 19329 11849 19332
rect 11791 19323 11849 19329
rect 12250 19320 12256 19332
rect 12308 19320 12314 19372
rect 13464 19369 13492 19400
rect 13998 19388 14004 19400
rect 14056 19388 14062 19440
rect 16114 19428 16120 19440
rect 14476 19400 16120 19428
rect 14476 19372 14504 19400
rect 16114 19388 16120 19400
rect 16172 19428 16178 19440
rect 16574 19428 16580 19440
rect 16172 19400 16580 19428
rect 16172 19388 16178 19400
rect 16574 19388 16580 19400
rect 16632 19428 16638 19440
rect 16776 19428 16804 19468
rect 16850 19456 16856 19508
rect 16908 19496 16914 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 16908 19468 17693 19496
rect 16908 19456 16914 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 20165 19499 20223 19505
rect 17681 19459 17739 19465
rect 17788 19468 19840 19496
rect 16632 19400 16712 19428
rect 16776 19400 16896 19428
rect 16632 19388 16638 19400
rect 13449 19363 13507 19369
rect 13449 19329 13461 19363
rect 13495 19329 13507 19363
rect 13722 19360 13728 19372
rect 13683 19332 13728 19360
rect 13449 19323 13507 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14458 19320 14464 19372
rect 14516 19320 14522 19372
rect 16390 19320 16396 19372
rect 16448 19320 16454 19372
rect 16684 19369 16712 19400
rect 16868 19390 16896 19400
rect 16927 19393 16985 19399
rect 16927 19390 16939 19393
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16868 19362 16939 19390
rect 16927 19359 16939 19362
rect 16973 19359 16985 19393
rect 17310 19388 17316 19440
rect 17368 19428 17374 19440
rect 17788 19428 17816 19468
rect 19518 19428 19524 19440
rect 17368 19400 17816 19428
rect 19168 19400 19524 19428
rect 17368 19388 17374 19400
rect 19168 19369 19196 19400
rect 19518 19388 19524 19400
rect 19576 19388 19582 19440
rect 19610 19388 19616 19440
rect 19668 19388 19674 19440
rect 16927 19353 16985 19359
rect 19153 19363 19211 19369
rect 16669 19323 16727 19329
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19395 19363 19453 19369
rect 19395 19329 19407 19363
rect 19441 19360 19453 19363
rect 19628 19360 19656 19388
rect 19812 19372 19840 19468
rect 20165 19465 20177 19499
rect 20211 19465 20223 19499
rect 20165 19459 20223 19465
rect 19441 19332 19656 19360
rect 19441 19329 19453 19332
rect 19395 19323 19453 19329
rect 19794 19320 19800 19372
rect 19852 19320 19858 19372
rect 20180 19360 20208 19459
rect 20806 19456 20812 19508
rect 20864 19456 20870 19508
rect 21177 19499 21235 19505
rect 21177 19465 21189 19499
rect 21223 19465 21235 19499
rect 21177 19459 21235 19465
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 22830 19496 22836 19508
rect 22419 19468 22836 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 21192 19428 21220 19459
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 23198 19456 23204 19508
rect 23256 19456 23262 19508
rect 23290 19456 23296 19508
rect 23348 19456 23354 19508
rect 23216 19428 23244 19456
rect 21192 19400 21864 19428
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 20180 19332 20545 19360
rect 20533 19329 20545 19332
rect 20579 19360 20591 19363
rect 20901 19363 20959 19369
rect 20901 19360 20913 19363
rect 20579 19332 20913 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20901 19329 20913 19332
rect 20947 19329 20959 19363
rect 20901 19323 20959 19329
rect 21082 19320 21088 19372
rect 21140 19320 21146 19372
rect 21266 19320 21272 19372
rect 21324 19360 21330 19372
rect 21836 19369 21864 19400
rect 22480 19400 23244 19428
rect 22480 19369 22508 19400
rect 21361 19363 21419 19369
rect 21361 19360 21373 19363
rect 21324 19332 21373 19360
rect 21324 19320 21330 19332
rect 21361 19329 21373 19332
rect 21407 19329 21419 19363
rect 21361 19323 21419 19329
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 21913 19363 21971 19369
rect 21913 19329 21925 19363
rect 21959 19360 21971 19363
rect 22097 19363 22155 19369
rect 21959 19332 22048 19360
rect 21959 19329 21971 19332
rect 21913 19323 21971 19329
rect 1670 19252 1676 19304
rect 1728 19252 1734 19304
rect 4246 19252 4252 19304
rect 4304 19292 4310 19304
rect 4304 19264 4382 19292
rect 4304 19252 4310 19264
rect 2332 19196 4292 19224
rect 198 19116 204 19168
rect 256 19156 262 19168
rect 2332 19156 2360 19196
rect 4264 19168 4292 19196
rect 256 19128 2360 19156
rect 256 19116 262 19128
rect 2682 19116 2688 19168
rect 2740 19116 2746 19168
rect 4246 19116 4252 19168
rect 4304 19116 4310 19168
rect 4354 19156 4382 19264
rect 7650 19252 7656 19304
rect 7708 19252 7714 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 11517 19295 11575 19301
rect 11517 19292 11529 19295
rect 11296 19264 11529 19292
rect 11296 19252 11302 19264
rect 11517 19261 11529 19264
rect 11563 19261 11575 19295
rect 16408 19292 16436 19320
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 16408 19264 16497 19292
rect 11517 19255 11575 19261
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20993 19295 21051 19301
rect 20993 19292 21005 19295
rect 20855 19264 21005 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20993 19261 21005 19264
rect 21039 19261 21051 19295
rect 22020 19292 22048 19332
rect 22097 19329 22109 19363
rect 22143 19360 22155 19363
rect 22465 19363 22523 19369
rect 22465 19360 22477 19363
rect 22143 19332 22477 19360
rect 22143 19329 22155 19332
rect 22097 19323 22155 19329
rect 22465 19329 22477 19332
rect 22511 19329 22523 19363
rect 22465 19323 22523 19329
rect 22646 19320 22652 19372
rect 22704 19320 22710 19372
rect 23106 19320 23112 19372
rect 23164 19360 23170 19372
rect 23308 19360 23336 19456
rect 23569 19431 23627 19437
rect 23569 19397 23581 19431
rect 23615 19428 23627 19431
rect 23934 19428 23940 19440
rect 23615 19400 23940 19428
rect 23615 19397 23627 19400
rect 23569 19391 23627 19397
rect 23934 19388 23940 19400
rect 23992 19388 23998 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23164 19332 23244 19360
rect 23308 19332 23397 19360
rect 23164 19320 23170 19332
rect 22189 19295 22247 19301
rect 22189 19292 22201 19295
rect 22020 19264 22201 19292
rect 20993 19255 21051 19261
rect 22189 19261 22201 19264
rect 22235 19261 22247 19295
rect 22189 19255 22247 19261
rect 22373 19295 22431 19301
rect 22373 19261 22385 19295
rect 22419 19292 22431 19295
rect 22557 19295 22615 19301
rect 22557 19292 22569 19295
rect 22419 19264 22569 19292
rect 22419 19261 22431 19264
rect 22373 19255 22431 19261
rect 22557 19261 22569 19264
rect 22603 19261 22615 19295
rect 22557 19255 22615 19261
rect 8389 19227 8447 19233
rect 8389 19193 8401 19227
rect 8435 19193 8447 19227
rect 20530 19224 20536 19236
rect 8389 19187 8447 19193
rect 9600 19196 11652 19224
rect 5350 19156 5356 19168
rect 4354 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 8404 19156 8432 19187
rect 9600 19156 9628 19196
rect 8404 19128 9628 19156
rect 9674 19116 9680 19168
rect 9732 19156 9738 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9732 19128 9873 19156
rect 9732 19116 9738 19128
rect 9861 19125 9873 19128
rect 9907 19125 9919 19159
rect 9861 19119 9919 19125
rect 9950 19116 9956 19168
rect 10008 19156 10014 19168
rect 10318 19156 10324 19168
rect 10008 19128 10324 19156
rect 10008 19116 10014 19128
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 11624 19156 11652 19196
rect 12406 19196 13584 19224
rect 12406 19156 12434 19196
rect 11624 19128 12434 19156
rect 12529 19159 12587 19165
rect 12529 19125 12541 19159
rect 12575 19156 12587 19159
rect 12710 19156 12716 19168
rect 12575 19128 12716 19156
rect 12575 19125 12587 19128
rect 12529 19119 12587 19125
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 13556 19156 13584 19196
rect 14384 19196 16804 19224
rect 14384 19156 14412 19196
rect 13556 19128 14412 19156
rect 14458 19116 14464 19168
rect 14516 19116 14522 19168
rect 14734 19116 14740 19168
rect 14792 19156 14798 19168
rect 15562 19156 15568 19168
rect 14792 19128 15568 19156
rect 14792 19116 14798 19128
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16776 19156 16804 19196
rect 20180 19196 20536 19224
rect 20180 19156 20208 19196
rect 20530 19184 20536 19196
rect 20588 19184 20594 19236
rect 21174 19184 21180 19236
rect 21232 19224 21238 19236
rect 23106 19224 23112 19236
rect 21232 19196 23112 19224
rect 21232 19184 21238 19196
rect 23106 19184 23112 19196
rect 23164 19184 23170 19236
rect 23216 19233 23244 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 24397 19295 24455 19301
rect 24397 19261 24409 19295
rect 24443 19292 24455 19295
rect 25130 19292 25136 19304
rect 24443 19264 25136 19292
rect 24443 19261 24455 19264
rect 24397 19255 24455 19261
rect 25130 19252 25136 19264
rect 25188 19252 25194 19304
rect 23201 19227 23259 19233
rect 23201 19193 23213 19227
rect 23247 19193 23259 19227
rect 23201 19187 23259 19193
rect 16776 19128 20208 19156
rect 20254 19116 20260 19168
rect 20312 19156 20318 19168
rect 20625 19159 20683 19165
rect 20625 19156 20637 19159
rect 20312 19128 20637 19156
rect 20312 19116 20318 19128
rect 20625 19125 20637 19128
rect 20671 19125 20683 19159
rect 20625 19119 20683 19125
rect 23842 19116 23848 19168
rect 23900 19116 23906 19168
rect 1104 19066 24840 19088
rect 1104 19014 3917 19066
rect 3969 19014 3981 19066
rect 4033 19014 4045 19066
rect 4097 19014 4109 19066
rect 4161 19014 4173 19066
rect 4225 19014 9851 19066
rect 9903 19014 9915 19066
rect 9967 19014 9979 19066
rect 10031 19014 10043 19066
rect 10095 19014 10107 19066
rect 10159 19014 15785 19066
rect 15837 19014 15849 19066
rect 15901 19014 15913 19066
rect 15965 19014 15977 19066
rect 16029 19014 16041 19066
rect 16093 19014 21719 19066
rect 21771 19014 21783 19066
rect 21835 19014 21847 19066
rect 21899 19014 21911 19066
rect 21963 19014 21975 19066
rect 22027 19014 24840 19066
rect 1104 18992 24840 19014
rect 1394 18912 1400 18964
rect 1452 18912 1458 18964
rect 4614 18952 4620 18964
rect 3252 18924 4620 18952
rect 1412 18816 1440 18912
rect 3252 18893 3280 18924
rect 4614 18912 4620 18924
rect 4672 18912 4678 18964
rect 7466 18912 7472 18964
rect 7524 18952 7530 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7524 18924 8125 18952
rect 7524 18912 7530 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 13814 18952 13820 18964
rect 10560 18924 13820 18952
rect 10560 18912 10566 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 16114 18912 16120 18964
rect 16172 18912 16178 18964
rect 16298 18912 16304 18964
rect 16356 18952 16362 18964
rect 17037 18955 17095 18961
rect 17037 18952 17049 18955
rect 16356 18924 17049 18952
rect 16356 18912 16362 18924
rect 17037 18921 17049 18924
rect 17083 18921 17095 18955
rect 17037 18915 17095 18921
rect 18598 18912 18604 18964
rect 18656 18912 18662 18964
rect 19705 18955 19763 18961
rect 19705 18921 19717 18955
rect 19751 18952 19763 18955
rect 20254 18952 20260 18964
rect 19751 18924 20260 18952
rect 19751 18921 19763 18924
rect 19705 18915 19763 18921
rect 20254 18912 20260 18924
rect 20312 18912 20318 18964
rect 21082 18912 21088 18964
rect 21140 18912 21146 18964
rect 3237 18887 3295 18893
rect 3237 18853 3249 18887
rect 3283 18853 3295 18887
rect 3237 18847 3295 18853
rect 4706 18844 4712 18896
rect 4764 18884 4770 18896
rect 4801 18887 4859 18893
rect 4801 18884 4813 18887
rect 4764 18856 4813 18884
rect 4764 18844 4770 18856
rect 4801 18853 4813 18856
rect 4847 18853 4859 18887
rect 4801 18847 4859 18853
rect 10413 18887 10471 18893
rect 10413 18853 10425 18887
rect 10459 18853 10471 18887
rect 10413 18847 10471 18853
rect 12084 18856 14320 18884
rect 8944 18828 8996 18834
rect 1578 18816 1584 18828
rect 1412 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 6638 18776 6644 18828
rect 6696 18816 6702 18828
rect 7101 18819 7159 18825
rect 7101 18816 7113 18819
rect 6696 18788 7113 18816
rect 6696 18776 6702 18788
rect 7101 18785 7113 18788
rect 7147 18785 7159 18819
rect 7101 18779 7159 18785
rect 8944 18770 8996 18776
rect 1855 18751 1913 18757
rect 1855 18717 1867 18751
rect 1901 18748 1913 18751
rect 2314 18748 2320 18760
rect 1901 18720 2320 18748
rect 1901 18717 1913 18720
rect 1855 18711 1913 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18748 3847 18751
rect 3835 18720 3924 18748
rect 4062 18747 4068 18760
rect 3835 18717 3847 18720
rect 3789 18711 3847 18717
rect 1302 18640 1308 18692
rect 1360 18680 1366 18692
rect 3053 18683 3111 18689
rect 3053 18680 3065 18683
rect 1360 18652 3065 18680
rect 1360 18640 1366 18652
rect 3053 18649 3065 18652
rect 3099 18649 3111 18683
rect 3053 18643 3111 18649
rect 3896 18624 3924 18720
rect 4047 18741 4068 18747
rect 4047 18707 4059 18741
rect 4120 18708 4126 18760
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 7375 18751 7433 18757
rect 7375 18748 7387 18751
rect 5868 18720 7387 18748
rect 5868 18708 5874 18720
rect 7375 18717 7387 18720
rect 7421 18717 7433 18751
rect 7375 18711 7433 18717
rect 8018 18708 8024 18760
rect 8076 18748 8082 18760
rect 9401 18751 9459 18757
rect 9401 18748 9413 18751
rect 8076 18738 8892 18748
rect 9048 18738 9413 18748
rect 8076 18720 9413 18738
rect 8076 18708 8082 18720
rect 8864 18710 9076 18720
rect 9401 18717 9413 18720
rect 9447 18717 9459 18751
rect 10428 18748 10456 18847
rect 12084 18828 12112 18856
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18816 14151 18819
rect 14182 18816 14188 18828
rect 14139 18788 14188 18816
rect 14139 18785 14151 18788
rect 14093 18779 14151 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 14292 18816 14320 18856
rect 14458 18844 14464 18896
rect 14516 18884 14522 18896
rect 14737 18887 14795 18893
rect 14737 18884 14749 18887
rect 14516 18856 14749 18884
rect 14516 18844 14522 18856
rect 14737 18853 14749 18856
rect 14783 18853 14795 18887
rect 16132 18884 16160 18912
rect 14737 18847 14795 18853
rect 16040 18856 16160 18884
rect 18616 18884 18644 18912
rect 19981 18887 20039 18893
rect 18616 18856 19656 18884
rect 15010 18816 15016 18828
rect 14292 18788 15016 18816
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 15102 18776 15108 18828
rect 15160 18825 15166 18828
rect 16040 18825 16068 18856
rect 15160 18819 15188 18825
rect 15176 18785 15188 18819
rect 15160 18779 15188 18785
rect 16025 18819 16083 18825
rect 16025 18785 16037 18819
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 15160 18776 15166 18779
rect 10428 18720 11192 18748
rect 9401 18711 9459 18717
rect 4093 18707 4105 18708
rect 4047 18701 4105 18707
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 9125 18683 9183 18689
rect 9125 18680 9137 18683
rect 8352 18652 9137 18680
rect 8352 18640 8358 18652
rect 9125 18649 9137 18652
rect 9171 18649 9183 18683
rect 9125 18643 9183 18649
rect 9490 18640 9496 18692
rect 9548 18640 9554 18692
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 10042 18640 10048 18692
rect 10100 18680 10106 18692
rect 10229 18683 10287 18689
rect 10229 18680 10241 18683
rect 10100 18652 10241 18680
rect 10100 18640 10106 18652
rect 10229 18649 10241 18652
rect 10275 18680 10287 18683
rect 10870 18680 10876 18692
rect 10275 18652 10876 18680
rect 10275 18649 10287 18652
rect 10229 18643 10287 18649
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 11164 18680 11192 18720
rect 11238 18708 11244 18760
rect 11296 18708 11302 18760
rect 11515 18751 11573 18757
rect 11515 18717 11527 18751
rect 11561 18748 11573 18751
rect 11606 18748 11612 18760
rect 11561 18720 11612 18748
rect 11561 18717 11573 18720
rect 11515 18711 11573 18717
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 14274 18708 14280 18760
rect 14332 18708 14338 18760
rect 15286 18708 15292 18760
rect 15344 18708 15350 18760
rect 16283 18721 16341 18727
rect 16283 18687 16295 18721
rect 16329 18718 16341 18721
rect 16329 18692 16344 18718
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 19628 18757 19656 18856
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 21100 18884 21128 18912
rect 23474 18884 23480 18896
rect 20027 18856 21128 18884
rect 22756 18856 23480 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 17589 18751 17647 18757
rect 17589 18748 17601 18751
rect 17184 18720 17601 18748
rect 17184 18708 17190 18720
rect 17589 18717 17601 18720
rect 17635 18717 17647 18751
rect 19613 18751 19671 18757
rect 17589 18711 17647 18717
rect 17847 18721 17905 18727
rect 16283 18681 16304 18687
rect 11164 18652 14320 18680
rect 934 18572 940 18624
rect 992 18612 998 18624
rect 1210 18612 1216 18624
rect 992 18584 1216 18612
rect 992 18572 998 18584
rect 1210 18572 1216 18584
rect 1268 18572 1274 18624
rect 2593 18615 2651 18621
rect 2593 18581 2605 18615
rect 2639 18612 2651 18615
rect 2866 18612 2872 18624
rect 2639 18584 2872 18612
rect 2639 18581 2651 18584
rect 2593 18575 2651 18581
rect 2866 18572 2872 18584
rect 2924 18572 2930 18624
rect 3878 18572 3884 18624
rect 3936 18572 3942 18624
rect 3970 18572 3976 18624
rect 4028 18612 4034 18624
rect 8662 18612 8668 18624
rect 4028 18584 8668 18612
rect 4028 18572 4034 18584
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 10594 18612 10600 18624
rect 9640 18584 10600 18612
rect 9640 18572 9646 18584
rect 10594 18572 10600 18584
rect 10652 18612 10658 18624
rect 12066 18612 12072 18624
rect 10652 18584 12072 18612
rect 10652 18572 10658 18584
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12250 18572 12256 18624
rect 12308 18572 12314 18624
rect 14292 18612 14320 18652
rect 16298 18640 16304 18681
rect 16356 18640 16362 18692
rect 17847 18687 17859 18721
rect 17893 18718 17905 18721
rect 17893 18687 17906 18718
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18748 20223 18751
rect 20622 18748 20628 18760
rect 20211 18720 20628 18748
rect 20211 18717 20223 18720
rect 20165 18711 20223 18717
rect 20622 18708 20628 18720
rect 20680 18708 20686 18760
rect 22756 18757 22784 18856
rect 23474 18844 23480 18856
rect 23532 18844 23538 18896
rect 23569 18887 23627 18893
rect 23569 18853 23581 18887
rect 23615 18884 23627 18887
rect 25130 18884 25136 18896
rect 23615 18856 25136 18884
rect 23615 18853 23627 18856
rect 23569 18847 23627 18853
rect 25130 18844 25136 18856
rect 25188 18844 25194 18896
rect 22833 18819 22891 18825
rect 22833 18785 22845 18819
rect 22879 18816 22891 18819
rect 23658 18816 23664 18828
rect 22879 18788 23664 18816
rect 22879 18785 22891 18788
rect 22833 18779 22891 18785
rect 23658 18776 23664 18788
rect 23716 18776 23722 18828
rect 24302 18816 24308 18828
rect 23860 18788 24308 18816
rect 22741 18751 22799 18757
rect 22741 18717 22753 18751
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23201 18751 23259 18757
rect 23201 18748 23213 18751
rect 23124 18720 23213 18748
rect 17847 18681 17906 18687
rect 17878 18680 17906 18681
rect 17878 18652 19334 18680
rect 14826 18612 14832 18624
rect 14292 18584 14832 18612
rect 14826 18572 14832 18584
rect 14884 18572 14890 18624
rect 15930 18572 15936 18624
rect 15988 18572 15994 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18380 18584 18613 18612
rect 18380 18572 18386 18584
rect 18601 18581 18613 18584
rect 18647 18581 18659 18615
rect 19306 18612 19334 18652
rect 23124 18624 23152 18720
rect 23201 18717 23213 18720
rect 23247 18717 23259 18751
rect 23201 18711 23259 18717
rect 23382 18708 23388 18760
rect 23440 18708 23446 18760
rect 23860 18757 23888 18788
rect 24302 18776 24308 18788
rect 24360 18776 24366 18828
rect 23845 18751 23903 18757
rect 23845 18717 23857 18751
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 24213 18751 24271 18757
rect 24213 18717 24225 18751
rect 24259 18748 24271 18751
rect 25498 18748 25504 18760
rect 24259 18720 25504 18748
rect 24259 18717 24271 18720
rect 24213 18711 24271 18717
rect 25498 18708 25504 18720
rect 25556 18708 25562 18760
rect 20898 18612 20904 18624
rect 19306 18584 20904 18612
rect 18601 18575 18659 18581
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 23014 18572 23020 18624
rect 23072 18572 23078 18624
rect 23106 18572 23112 18624
rect 23164 18572 23170 18624
rect 1104 18522 25000 18544
rect 1104 18470 6884 18522
rect 6936 18470 6948 18522
rect 7000 18470 7012 18522
rect 7064 18470 7076 18522
rect 7128 18470 7140 18522
rect 7192 18470 12818 18522
rect 12870 18470 12882 18522
rect 12934 18470 12946 18522
rect 12998 18470 13010 18522
rect 13062 18470 13074 18522
rect 13126 18470 18752 18522
rect 18804 18470 18816 18522
rect 18868 18470 18880 18522
rect 18932 18470 18944 18522
rect 18996 18470 19008 18522
rect 19060 18470 24686 18522
rect 24738 18470 24750 18522
rect 24802 18470 24814 18522
rect 24866 18470 24878 18522
rect 24930 18470 24942 18522
rect 24994 18470 25000 18522
rect 1104 18448 25000 18470
rect 1857 18411 1915 18417
rect 1857 18377 1869 18411
rect 1903 18408 1915 18411
rect 1946 18408 1952 18420
rect 1903 18380 1952 18408
rect 1903 18377 1915 18380
rect 1857 18371 1915 18377
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2130 18368 2136 18420
rect 2188 18408 2194 18420
rect 3970 18408 3976 18420
rect 2188 18380 3976 18408
rect 2188 18368 2194 18380
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4246 18368 4252 18420
rect 4304 18408 4310 18420
rect 5537 18411 5595 18417
rect 5537 18408 5549 18411
rect 4304 18380 5549 18408
rect 4304 18368 4310 18380
rect 5537 18377 5549 18380
rect 5583 18377 5595 18411
rect 8294 18408 8300 18420
rect 5537 18371 5595 18377
rect 8036 18380 8300 18408
rect 1210 18300 1216 18352
rect 1268 18340 1274 18352
rect 3513 18343 3571 18349
rect 3513 18340 3525 18343
rect 1268 18312 3525 18340
rect 1268 18300 1274 18312
rect 3513 18309 3525 18312
rect 3559 18309 3571 18343
rect 5810 18340 5816 18352
rect 3513 18303 3571 18309
rect 4356 18312 5816 18340
rect 1670 18232 1676 18284
rect 1728 18232 1734 18284
rect 1762 18232 1768 18284
rect 1820 18232 1826 18284
rect 2314 18272 2320 18284
rect 2275 18244 2320 18272
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 4246 18232 4252 18284
rect 4304 18282 4310 18284
rect 4356 18282 4384 18312
rect 5810 18300 5816 18312
rect 5868 18300 5874 18352
rect 4304 18254 4384 18282
rect 4304 18244 4347 18254
rect 4304 18232 4310 18244
rect 5166 18232 5172 18284
rect 5224 18272 5230 18284
rect 5445 18275 5503 18281
rect 5445 18272 5457 18275
rect 5224 18244 5457 18272
rect 5224 18232 5230 18244
rect 5445 18241 5457 18244
rect 5491 18241 5503 18275
rect 8036 18272 8064 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8938 18368 8944 18420
rect 8996 18408 9002 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 8996 18380 9229 18408
rect 8996 18368 9002 18380
rect 9217 18377 9229 18380
rect 9263 18377 9275 18411
rect 9217 18371 9275 18377
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 15197 18411 15255 18417
rect 9548 18380 15148 18408
rect 9548 18368 9554 18380
rect 8110 18300 8116 18352
rect 8168 18340 8174 18352
rect 8168 18312 8614 18340
rect 8168 18300 8174 18312
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 8036 18244 8217 18272
rect 5445 18235 5503 18241
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 8478 18272 8484 18284
rect 8439 18244 8484 18272
rect 8205 18235 8263 18241
rect 8478 18232 8484 18244
rect 8536 18232 8542 18284
rect 8586 18272 8614 18312
rect 8754 18300 8760 18352
rect 8812 18340 8818 18352
rect 9582 18340 9588 18352
rect 8812 18312 9588 18340
rect 8812 18300 8818 18312
rect 9582 18300 9588 18312
rect 9640 18300 9646 18352
rect 10686 18340 10692 18352
rect 9876 18312 10692 18340
rect 9876 18311 9904 18312
rect 9843 18305 9904 18311
rect 9843 18272 9855 18305
rect 8586 18271 9855 18272
rect 9889 18271 9904 18305
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 11701 18343 11759 18349
rect 11701 18309 11713 18343
rect 11747 18340 11759 18343
rect 11790 18340 11796 18352
rect 11747 18312 11796 18340
rect 11747 18309 11759 18312
rect 11701 18303 11759 18309
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 12618 18300 12624 18352
rect 12676 18340 12682 18352
rect 12805 18343 12863 18349
rect 12805 18340 12817 18343
rect 12676 18312 12817 18340
rect 12676 18300 12682 18312
rect 12805 18309 12817 18312
rect 12851 18309 12863 18343
rect 13814 18340 13820 18352
rect 12805 18303 12863 18309
rect 13096 18312 13820 18340
rect 8586 18244 9904 18271
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11379 18244 11989 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12216 18244 12449 18272
rect 12216 18232 12222 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 1688 18204 1716 18232
rect 12716 18216 12768 18222
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1688 18176 2053 18204
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 3970 18164 3976 18216
rect 4028 18164 4034 18216
rect 9582 18164 9588 18216
rect 9640 18164 9646 18216
rect 12716 18158 12768 18164
rect 13096 18148 13124 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 15120 18340 15148 18380
rect 15197 18377 15209 18411
rect 15243 18408 15255 18411
rect 15286 18408 15292 18420
rect 15243 18380 15292 18408
rect 15243 18377 15255 18380
rect 15197 18371 15255 18377
rect 15286 18368 15292 18380
rect 15344 18368 15350 18420
rect 15396 18380 18828 18408
rect 15396 18340 15424 18380
rect 15120 18312 15424 18340
rect 18800 18340 18828 18380
rect 21358 18368 21364 18420
rect 21416 18408 21422 18420
rect 21416 18380 24164 18408
rect 21416 18368 21422 18380
rect 22802 18343 22860 18349
rect 22802 18340 22814 18343
rect 18800 18312 22814 18340
rect 22802 18309 22814 18312
rect 22848 18340 22860 18343
rect 23106 18340 23112 18352
rect 22848 18312 23112 18340
rect 22848 18309 22860 18312
rect 22802 18303 22860 18309
rect 23106 18300 23112 18312
rect 23164 18300 23170 18352
rect 24136 18349 24164 18380
rect 24121 18343 24179 18349
rect 24121 18309 24133 18343
rect 24167 18309 24179 18343
rect 24121 18303 24179 18309
rect 13998 18232 14004 18284
rect 14056 18272 14062 18284
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 14056 18244 14197 18272
rect 14056 18232 14062 18244
rect 14185 18241 14197 18244
rect 14231 18241 14243 18275
rect 14458 18272 14464 18284
rect 14419 18244 14464 18272
rect 14185 18235 14243 18241
rect 14458 18232 14464 18244
rect 14516 18232 14522 18284
rect 17129 18275 17187 18281
rect 17129 18241 17141 18275
rect 17175 18272 17187 18275
rect 17218 18272 17224 18284
rect 17175 18244 17224 18272
rect 17175 18241 17187 18244
rect 17129 18235 17187 18241
rect 17218 18232 17224 18244
rect 17276 18232 17282 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17494 18272 17500 18284
rect 17359 18244 17500 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 11330 18136 11336 18148
rect 4908 18108 8340 18136
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18037 3111 18071
rect 3053 18031 3111 18037
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4908 18068 4936 18108
rect 3651 18040 4936 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4982 18028 4988 18080
rect 5040 18028 5046 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 7282 18068 7288 18080
rect 5408 18040 7288 18068
rect 5408 18028 5414 18040
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 8312 18068 8340 18108
rect 10428 18108 11336 18136
rect 10428 18068 10456 18108
rect 11330 18096 11336 18108
rect 11388 18096 11394 18148
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18136 13047 18139
rect 13078 18136 13084 18148
rect 13035 18108 13084 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 13078 18096 13084 18108
rect 13136 18096 13142 18148
rect 17328 18136 17356 18235
rect 17494 18232 17500 18244
rect 17552 18232 17558 18284
rect 18322 18232 18328 18284
rect 18380 18232 18386 18284
rect 20990 18232 20996 18284
rect 21048 18232 21054 18284
rect 18046 18164 18052 18216
rect 18104 18164 18110 18216
rect 18187 18207 18245 18213
rect 18187 18173 18199 18207
rect 18233 18204 18245 18207
rect 21008 18204 21036 18232
rect 18233 18176 21036 18204
rect 18233 18173 18245 18176
rect 18187 18167 18245 18173
rect 14844 18108 17356 18136
rect 17773 18139 17831 18145
rect 8312 18040 10456 18068
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10597 18071 10655 18077
rect 10597 18068 10609 18071
rect 10560 18040 10609 18068
rect 10560 18028 10566 18040
rect 10597 18037 10609 18040
rect 10643 18037 10655 18071
rect 10597 18031 10655 18037
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 14844 18068 14872 18108
rect 17773 18105 17785 18139
rect 17819 18136 17831 18139
rect 17862 18136 17868 18148
rect 17819 18108 17868 18136
rect 17819 18105 17831 18108
rect 17773 18099 17831 18105
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 14332 18040 14872 18068
rect 14332 18028 14338 18040
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 18708 18068 18736 18176
rect 21266 18164 21272 18216
rect 21324 18204 21330 18216
rect 22370 18204 22376 18216
rect 21324 18176 22376 18204
rect 21324 18164 21330 18176
rect 22370 18164 22376 18176
rect 22428 18204 22434 18216
rect 22557 18207 22615 18213
rect 22557 18204 22569 18207
rect 22428 18176 22569 18204
rect 22428 18164 22434 18176
rect 22557 18173 22569 18176
rect 22603 18173 22615 18207
rect 22557 18167 22615 18173
rect 16172 18040 18736 18068
rect 18969 18071 19027 18077
rect 16172 18028 16178 18040
rect 18969 18037 18981 18071
rect 19015 18068 19027 18071
rect 19426 18068 19432 18080
rect 19015 18040 19432 18068
rect 19015 18037 19027 18040
rect 18969 18031 19027 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 23566 18028 23572 18080
rect 23624 18068 23630 18080
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23624 18040 23949 18068
rect 23624 18028 23630 18040
rect 23937 18037 23949 18040
rect 23983 18037 23995 18071
rect 23937 18031 23995 18037
rect 24394 18028 24400 18080
rect 24452 18028 24458 18080
rect 1104 17978 24840 18000
rect 1104 17926 3917 17978
rect 3969 17926 3981 17978
rect 4033 17926 4045 17978
rect 4097 17926 4109 17978
rect 4161 17926 4173 17978
rect 4225 17926 9851 17978
rect 9903 17926 9915 17978
rect 9967 17926 9979 17978
rect 10031 17926 10043 17978
rect 10095 17926 10107 17978
rect 10159 17926 15785 17978
rect 15837 17926 15849 17978
rect 15901 17926 15913 17978
rect 15965 17926 15977 17978
rect 16029 17926 16041 17978
rect 16093 17926 21719 17978
rect 21771 17926 21783 17978
rect 21835 17926 21847 17978
rect 21899 17926 21911 17978
rect 21963 17926 21975 17978
rect 22027 17926 24840 17978
rect 1104 17904 24840 17926
rect 2682 17864 2688 17876
rect 2424 17836 2688 17864
rect 2424 17805 2452 17836
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 3694 17864 3700 17876
rect 2832 17836 3700 17864
rect 2832 17824 2838 17836
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 4706 17864 4712 17876
rect 4448 17836 4712 17864
rect 2409 17799 2467 17805
rect 2409 17765 2421 17799
rect 2455 17765 2467 17799
rect 3602 17796 3608 17808
rect 2409 17759 2467 17765
rect 3436 17768 3608 17796
rect 1949 17731 2007 17737
rect 1949 17697 1961 17731
rect 1995 17728 2007 17731
rect 3436 17728 3464 17768
rect 3602 17756 3608 17768
rect 3660 17796 3666 17808
rect 4448 17805 4476 17836
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 14274 17864 14280 17876
rect 5644 17836 14280 17864
rect 4433 17799 4491 17805
rect 3660 17768 3924 17796
rect 3660 17756 3666 17768
rect 1995 17700 3464 17728
rect 1995 17697 2007 17700
rect 1949 17691 2007 17697
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3568 17700 3801 17728
rect 3568 17688 3574 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3896 17728 3924 17768
rect 4433 17765 4445 17799
rect 4479 17765 4491 17799
rect 4433 17759 4491 17765
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 3896 17700 4721 17728
rect 3789 17691 3847 17697
rect 4709 17697 4721 17700
rect 4755 17697 4767 17731
rect 5350 17728 5356 17740
rect 4709 17691 4767 17697
rect 4862 17700 5356 17728
rect 1394 17620 1400 17672
rect 1452 17620 1458 17672
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1811 17632 1992 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 1964 17604 1992 17632
rect 2682 17620 2688 17672
rect 2740 17620 2746 17672
rect 2774 17620 2780 17672
rect 2832 17669 2838 17672
rect 2832 17663 2860 17669
rect 2848 17629 2860 17663
rect 2832 17623 2860 17629
rect 2832 17620 2838 17623
rect 2958 17620 2964 17672
rect 3016 17620 3022 17672
rect 3970 17620 3976 17672
rect 4028 17620 4034 17672
rect 4862 17669 4890 17700
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 4847 17663 4905 17669
rect 4847 17629 4859 17663
rect 4893 17629 4905 17663
rect 4847 17623 4905 17629
rect 4982 17620 4988 17672
rect 5040 17620 5046 17672
rect 1946 17552 1952 17604
rect 2004 17552 2010 17604
rect 5644 17592 5672 17836
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 18141 17867 18199 17873
rect 18141 17864 18153 17867
rect 17920 17836 18153 17864
rect 17920 17824 17926 17836
rect 18141 17833 18153 17836
rect 18187 17833 18199 17867
rect 18141 17827 18199 17833
rect 22554 17824 22560 17876
rect 22612 17864 22618 17876
rect 22612 17836 22784 17864
rect 22612 17824 22618 17836
rect 5994 17756 6000 17808
rect 6052 17756 6058 17808
rect 10413 17799 10471 17805
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 10502 17796 10508 17808
rect 10459 17768 10508 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 18693 17799 18751 17805
rect 18693 17796 18705 17799
rect 18104 17768 18705 17796
rect 18104 17756 18110 17768
rect 18693 17765 18705 17768
rect 18739 17765 18751 17799
rect 18693 17759 18751 17765
rect 22097 17799 22155 17805
rect 22097 17765 22109 17799
rect 22143 17796 22155 17799
rect 22143 17768 22692 17796
rect 22143 17765 22155 17768
rect 22097 17759 22155 17765
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 3528 17564 4016 17592
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 3528 17524 3556 17564
rect 1627 17496 3556 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 3602 17484 3608 17536
rect 3660 17484 3666 17536
rect 3988 17524 4016 17564
rect 5552 17564 5672 17592
rect 5736 17700 6101 17728
rect 5736 17592 5764 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 9858 17688 9864 17740
rect 9916 17728 9922 17740
rect 10806 17731 10864 17737
rect 10806 17728 10818 17731
rect 9916 17700 10818 17728
rect 9916 17688 9922 17700
rect 10806 17697 10818 17700
rect 10852 17697 10864 17731
rect 10806 17691 10864 17697
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11388 17700 12265 17728
rect 11388 17688 11394 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 12710 17688 12716 17740
rect 12768 17688 12774 17740
rect 12989 17731 13047 17737
rect 12989 17697 13001 17731
rect 13035 17728 13047 17731
rect 14277 17731 14335 17737
rect 14277 17728 14289 17731
rect 13035 17700 14289 17728
rect 13035 17697 13047 17700
rect 12989 17691 13047 17697
rect 14277 17697 14289 17700
rect 14323 17697 14335 17731
rect 14277 17691 14335 17697
rect 5810 17620 5816 17672
rect 5868 17660 5874 17672
rect 6363 17663 6421 17669
rect 6363 17660 6375 17663
rect 5868 17632 6375 17660
rect 5868 17620 5874 17632
rect 6363 17629 6375 17632
rect 6409 17660 6421 17663
rect 6730 17660 6736 17672
rect 6409 17632 6736 17660
rect 6409 17629 6421 17632
rect 6363 17623 6421 17629
rect 6730 17620 6736 17632
rect 6788 17620 6794 17672
rect 7282 17620 7288 17672
rect 7340 17660 7346 17672
rect 9953 17663 10011 17669
rect 9953 17660 9965 17663
rect 7340 17632 9965 17660
rect 7340 17620 7346 17632
rect 9953 17629 9965 17632
rect 9999 17660 10011 17663
rect 10134 17660 10140 17672
rect 9999 17632 10140 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 10962 17620 10968 17672
rect 11020 17620 11026 17672
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17660 11667 17663
rect 11701 17663 11759 17669
rect 11701 17660 11713 17663
rect 11655 17632 11713 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 11701 17629 11713 17632
rect 11747 17629 11759 17663
rect 11882 17660 11888 17672
rect 11701 17623 11759 17629
rect 11808 17632 11888 17660
rect 5902 17592 5908 17604
rect 5736 17564 5908 17592
rect 5552 17524 5580 17564
rect 5902 17552 5908 17564
rect 5960 17592 5966 17604
rect 5960 17564 9996 17592
rect 5960 17552 5966 17564
rect 3988 17496 5580 17524
rect 5629 17527 5687 17533
rect 5629 17493 5641 17527
rect 5675 17524 5687 17527
rect 5810 17524 5816 17536
rect 5675 17496 5816 17524
rect 5675 17493 5687 17496
rect 5629 17487 5687 17493
rect 5810 17484 5816 17496
rect 5868 17484 5874 17536
rect 7101 17527 7159 17533
rect 7101 17493 7113 17527
rect 7147 17524 7159 17527
rect 7466 17524 7472 17536
rect 7147 17496 7472 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 9306 17484 9312 17536
rect 9364 17524 9370 17536
rect 9858 17524 9864 17536
rect 9364 17496 9864 17524
rect 9364 17484 9370 17496
rect 9858 17484 9864 17496
rect 9916 17484 9922 17536
rect 9968 17524 9996 17564
rect 10502 17524 10508 17536
rect 9968 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11808 17524 11836 17632
rect 11882 17620 11888 17632
rect 11940 17620 11946 17672
rect 12069 17663 12127 17669
rect 12069 17629 12081 17663
rect 12115 17660 12127 17663
rect 12158 17660 12164 17672
rect 12115 17632 12164 17660
rect 12115 17629 12127 17632
rect 12069 17623 12127 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 13078 17620 13084 17672
rect 13136 17669 13142 17672
rect 13136 17663 13164 17669
rect 13152 17629 13164 17663
rect 13136 17623 13164 17629
rect 13136 17620 13142 17623
rect 13262 17620 13268 17672
rect 13320 17620 13326 17672
rect 17126 17660 17132 17672
rect 13832 17632 17132 17660
rect 10928 17496 11836 17524
rect 10928 17484 10934 17496
rect 11882 17484 11888 17536
rect 11940 17484 11946 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 13832 17524 13860 17632
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 17371 17663 17429 17669
rect 17371 17660 17383 17663
rect 17236 17632 17383 17660
rect 15470 17552 15476 17604
rect 15528 17592 15534 17604
rect 17236 17592 17264 17632
rect 17371 17629 17383 17632
rect 17417 17660 17429 17663
rect 17494 17660 17500 17672
rect 17417 17632 17500 17660
rect 17417 17629 17429 17632
rect 17371 17623 17429 17629
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19512 17663 19570 17669
rect 19512 17629 19524 17663
rect 19558 17629 19570 17663
rect 20717 17663 20775 17669
rect 20717 17660 20729 17663
rect 19512 17623 19570 17629
rect 19628 17632 20729 17660
rect 15528 17564 17264 17592
rect 15528 17552 15534 17564
rect 12492 17496 13860 17524
rect 13909 17527 13967 17533
rect 12492 17484 12498 17496
rect 13909 17493 13921 17527
rect 13955 17524 13967 17527
rect 18506 17524 18512 17536
rect 13955 17496 18512 17524
rect 13955 17493 13967 17496
rect 13909 17487 13967 17493
rect 18506 17484 18512 17496
rect 18564 17484 18570 17536
rect 19260 17524 19288 17623
rect 19426 17552 19432 17604
rect 19484 17592 19490 17604
rect 19536 17592 19564 17623
rect 19484 17564 19564 17592
rect 19484 17552 19490 17564
rect 19628 17536 19656 17632
rect 20717 17629 20729 17632
rect 20763 17660 20775 17663
rect 21266 17660 21272 17672
rect 20763 17632 21272 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 22186 17620 22192 17672
rect 22244 17620 22250 17672
rect 22664 17669 22692 17768
rect 22756 17737 22784 17836
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 23753 17867 23811 17873
rect 23753 17864 23765 17867
rect 23532 17836 23765 17864
rect 23532 17824 23538 17836
rect 23753 17833 23765 17836
rect 23799 17833 23811 17867
rect 23753 17827 23811 17833
rect 22741 17731 22799 17737
rect 22741 17697 22753 17731
rect 22787 17697 22799 17731
rect 22741 17691 22799 17697
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 23032 17639 23244 17660
rect 22649 17623 22707 17629
rect 22999 17633 23244 17639
rect 20973 17595 21031 17601
rect 20973 17592 20985 17595
rect 20916 17564 20985 17592
rect 19610 17524 19616 17536
rect 19260 17496 19616 17524
rect 19610 17484 19616 17496
rect 19668 17484 19674 17536
rect 20622 17484 20628 17536
rect 20680 17484 20686 17536
rect 20714 17484 20720 17536
rect 20772 17524 20778 17536
rect 20916 17524 20944 17564
rect 20973 17561 20985 17564
rect 21019 17561 21031 17595
rect 22999 17599 23011 17633
rect 23045 17632 23244 17633
rect 23045 17602 23060 17632
rect 23045 17599 23057 17602
rect 22999 17593 23057 17599
rect 20973 17555 21031 17561
rect 22066 17564 22324 17592
rect 20772 17496 20944 17524
rect 20772 17484 20778 17496
rect 21634 17484 21640 17536
rect 21692 17524 21698 17536
rect 22066 17524 22094 17564
rect 22296 17533 22324 17564
rect 23216 17536 23244 17632
rect 24302 17620 24308 17672
rect 24360 17660 24366 17672
rect 24578 17660 24584 17672
rect 24360 17632 24584 17660
rect 24360 17620 24366 17632
rect 24578 17620 24584 17632
rect 24636 17620 24642 17672
rect 21692 17496 22094 17524
rect 22281 17527 22339 17533
rect 21692 17484 21698 17496
rect 22281 17493 22293 17527
rect 22327 17493 22339 17527
rect 22281 17487 22339 17493
rect 22462 17484 22468 17536
rect 22520 17484 22526 17536
rect 23198 17484 23204 17536
rect 23256 17484 23262 17536
rect 1104 17434 25000 17456
rect 1104 17382 6884 17434
rect 6936 17382 6948 17434
rect 7000 17382 7012 17434
rect 7064 17382 7076 17434
rect 7128 17382 7140 17434
rect 7192 17382 12818 17434
rect 12870 17382 12882 17434
rect 12934 17382 12946 17434
rect 12998 17382 13010 17434
rect 13062 17382 13074 17434
rect 13126 17382 18752 17434
rect 18804 17382 18816 17434
rect 18868 17382 18880 17434
rect 18932 17382 18944 17434
rect 18996 17382 19008 17434
rect 19060 17382 24686 17434
rect 24738 17382 24750 17434
rect 24802 17382 24814 17434
rect 24866 17382 24878 17434
rect 24930 17382 24942 17434
rect 24994 17382 25000 17434
rect 1104 17360 25000 17382
rect 3602 17320 3608 17332
rect 1596 17292 3608 17320
rect 1596 17193 1624 17292
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 4246 17280 4252 17332
rect 4304 17280 4310 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6420 17292 7604 17320
rect 6420 17280 6426 17292
rect 4264 17252 4292 17280
rect 5350 17252 5356 17264
rect 4264 17224 5356 17252
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 1719 17156 1992 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 1964 17128 1992 17156
rect 2866 17144 2872 17196
rect 2924 17144 2930 17196
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17184 3847 17187
rect 4798 17184 4804 17196
rect 3835 17156 4804 17184
rect 3835 17153 3847 17156
rect 3789 17147 3847 17153
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5150 17193 5178 17224
rect 5350 17212 5356 17224
rect 5408 17212 5414 17264
rect 6454 17212 6460 17264
rect 6512 17212 6518 17264
rect 6546 17212 6552 17264
rect 6604 17212 6610 17264
rect 6917 17255 6975 17261
rect 6917 17221 6929 17255
rect 6963 17252 6975 17255
rect 7466 17252 7472 17264
rect 6963 17224 7472 17252
rect 6963 17221 6975 17224
rect 6917 17215 6975 17221
rect 7466 17212 7472 17224
rect 7524 17212 7530 17264
rect 7576 17252 7604 17292
rect 7650 17280 7656 17332
rect 7708 17280 7714 17332
rect 10502 17280 10508 17332
rect 10560 17320 10566 17332
rect 10560 17292 10916 17320
rect 10560 17280 10566 17292
rect 9582 17252 9588 17264
rect 7576 17224 7770 17252
rect 5135 17187 5193 17193
rect 5135 17153 5147 17187
rect 5181 17153 5193 17187
rect 5135 17147 5193 17153
rect 5902 17144 5908 17196
rect 5960 17144 5966 17196
rect 6472 17184 6500 17212
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6472 17156 6837 17184
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7650 17184 7656 17196
rect 7331 17156 7656 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 1854 17076 1860 17128
rect 1912 17076 1918 17128
rect 1946 17076 1952 17128
rect 2004 17076 2010 17128
rect 2317 17119 2375 17125
rect 2317 17085 2329 17119
rect 2363 17116 2375 17119
rect 2406 17116 2412 17128
rect 2363 17088 2412 17116
rect 2363 17085 2375 17088
rect 2317 17079 2375 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 2590 17076 2596 17128
rect 2648 17076 2654 17128
rect 2731 17119 2789 17125
rect 2731 17085 2743 17119
rect 2777 17116 2789 17119
rect 4430 17116 4436 17128
rect 2777 17088 4436 17116
rect 2777 17085 2789 17088
rect 2731 17079 2789 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 4893 17119 4951 17125
rect 4893 17085 4905 17119
rect 4939 17085 4951 17119
rect 5920 17116 5948 17144
rect 4893 17079 4951 17085
rect 5552 17088 5948 17116
rect 1397 16983 1455 16989
rect 1397 16949 1409 16983
rect 1443 16980 1455 16983
rect 1578 16980 1584 16992
rect 1443 16952 1584 16980
rect 1443 16949 1455 16952
rect 1397 16943 1455 16949
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 3510 16940 3516 16992
rect 3568 16940 3574 16992
rect 3605 16983 3663 16989
rect 3605 16949 3617 16983
rect 3651 16980 3663 16983
rect 3786 16980 3792 16992
rect 3651 16952 3792 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 3786 16940 3792 16952
rect 3844 16940 3850 16992
rect 4908 16980 4936 17079
rect 5552 16980 5580 17088
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 6380 17048 6408 17102
rect 5951 17020 6408 17048
rect 7742 17048 7770 17224
rect 8680 17224 9588 17252
rect 8680 17196 8708 17224
rect 9582 17212 9588 17224
rect 9640 17252 9646 17264
rect 10888 17252 10916 17292
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 11057 17323 11115 17329
rect 11057 17320 11069 17323
rect 11020 17292 11069 17320
rect 11020 17280 11026 17292
rect 11057 17289 11069 17292
rect 11103 17289 11115 17323
rect 11057 17283 11115 17289
rect 13262 17280 13268 17332
rect 13320 17320 13326 17332
rect 13633 17323 13691 17329
rect 13633 17320 13645 17323
rect 13320 17292 13645 17320
rect 13320 17280 13326 17292
rect 13633 17289 13645 17292
rect 13679 17289 13691 17323
rect 13633 17283 13691 17289
rect 19426 17280 19432 17332
rect 19484 17280 19490 17332
rect 19521 17323 19579 17329
rect 19521 17289 19533 17323
rect 19567 17289 19579 17323
rect 19521 17283 19579 17289
rect 11238 17252 11244 17264
rect 9640 17224 10849 17252
rect 10888 17224 11244 17252
rect 9640 17212 9646 17224
rect 8662 17144 8668 17196
rect 8720 17144 8726 17196
rect 10060 17193 10088 17224
rect 10045 17187 10103 17193
rect 10045 17153 10057 17187
rect 10091 17153 10103 17187
rect 10045 17147 10103 17153
rect 10226 17144 10232 17196
rect 10284 17184 10290 17196
rect 10319 17187 10377 17193
rect 10319 17184 10331 17187
rect 10284 17156 10331 17184
rect 10284 17144 10290 17156
rect 10319 17153 10331 17156
rect 10365 17184 10377 17187
rect 10410 17184 10416 17196
rect 10365 17156 10416 17184
rect 10365 17153 10377 17156
rect 10319 17147 10377 17153
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 10821 17116 10849 17224
rect 11238 17212 11244 17224
rect 11296 17212 11302 17264
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 13538 17252 13544 17264
rect 12216 17224 12480 17252
rect 12216 17212 12222 17224
rect 12452 17196 12480 17224
rect 12910 17224 13544 17252
rect 12250 17144 12256 17196
rect 12308 17144 12314 17196
rect 12434 17144 12440 17196
rect 12492 17184 12498 17196
rect 12910 17193 12938 17224
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 14550 17212 14556 17264
rect 14608 17252 14614 17264
rect 14608 17224 16954 17252
rect 14608 17212 14614 17224
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12492 17156 12633 17184
rect 12492 17144 12498 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12895 17187 12953 17193
rect 12895 17153 12907 17187
rect 12941 17153 12953 17187
rect 12895 17147 12953 17153
rect 13722 17144 13728 17196
rect 13780 17184 13786 17196
rect 15439 17187 15497 17193
rect 15439 17184 15451 17187
rect 13780 17156 15451 17184
rect 13780 17144 13786 17156
rect 15439 17153 15451 17156
rect 15485 17184 15497 17187
rect 16574 17184 16580 17196
rect 15485 17156 16580 17184
rect 15485 17153 15497 17156
rect 15439 17147 15497 17153
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 16926 17193 16954 17224
rect 16911 17187 16969 17193
rect 16911 17153 16923 17187
rect 16957 17184 16969 17187
rect 17034 17184 17040 17196
rect 16957 17156 17040 17184
rect 16957 17153 16969 17156
rect 16911 17147 16969 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 19444 17184 19472 17280
rect 19536 17252 19564 17283
rect 20622 17280 20628 17332
rect 20680 17280 20686 17332
rect 20993 17323 21051 17329
rect 20993 17289 21005 17323
rect 21039 17320 21051 17323
rect 22186 17320 22192 17332
rect 21039 17292 22192 17320
rect 21039 17289 21051 17292
rect 20993 17283 21051 17289
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22462 17280 22468 17332
rect 22520 17280 22526 17332
rect 23014 17280 23020 17332
rect 23072 17280 23078 17332
rect 23569 17323 23627 17329
rect 23569 17289 23581 17323
rect 23615 17320 23627 17323
rect 25130 17320 25136 17332
rect 23615 17292 25136 17320
rect 23615 17289 23627 17292
rect 23569 17283 23627 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 19536 17224 20116 17252
rect 20088 17193 20116 17224
rect 19705 17187 19763 17193
rect 19705 17184 19717 17187
rect 19444 17156 19717 17184
rect 19705 17153 19717 17156
rect 19751 17153 19763 17187
rect 19705 17147 19763 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17153 20131 17187
rect 20640 17184 20668 17280
rect 21082 17212 21088 17264
rect 21140 17252 21146 17264
rect 22480 17252 22508 17280
rect 21140 17224 21579 17252
rect 21140 17212 21146 17224
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20640 17156 20729 17184
rect 20073 17147 20131 17153
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 10821 17088 12678 17116
rect 7834 17048 7840 17060
rect 7742 17020 7840 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 11882 17008 11888 17060
rect 11940 17008 11946 17060
rect 4908 16952 5580 16980
rect 10502 16940 10508 16992
rect 10560 16980 10566 16992
rect 11900 16980 11928 17008
rect 10560 16952 11928 16980
rect 10560 16940 10566 16952
rect 12434 16940 12440 16992
rect 12492 16940 12498 16992
rect 12650 16980 12678 17088
rect 14384 17088 15209 17116
rect 14384 16980 14412 17088
rect 15197 17085 15209 17088
rect 15243 17085 15255 17119
rect 16482 17116 16488 17128
rect 15197 17079 15255 17085
rect 15856 17088 16488 17116
rect 12650 16952 14412 16980
rect 14458 16940 14464 16992
rect 14516 16940 14522 16992
rect 15212 16980 15240 17079
rect 15856 16980 15884 17088
rect 16482 17076 16488 17088
rect 16540 17116 16546 17128
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16540 17088 16681 17116
rect 16540 17076 16546 17088
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 19886 17076 19892 17128
rect 19944 17116 19950 17128
rect 20438 17116 20444 17128
rect 19944 17088 20444 17116
rect 19944 17076 19950 17088
rect 20438 17076 20444 17088
rect 20496 17076 20502 17128
rect 20530 17076 20536 17128
rect 20588 17076 20594 17128
rect 20548 17048 20576 17076
rect 21192 17048 21220 17147
rect 21468 17060 21496 17147
rect 21551 17116 21579 17224
rect 21652 17224 22508 17252
rect 23032 17252 23060 17280
rect 23032 17224 24348 17252
rect 21652 17193 21680 17224
rect 21637 17187 21695 17193
rect 21637 17153 21649 17187
rect 21683 17153 21695 17187
rect 22063 17187 22121 17193
rect 22063 17184 22075 17187
rect 21637 17147 21695 17153
rect 21744 17156 22075 17184
rect 21744 17116 21772 17156
rect 22063 17153 22075 17156
rect 22109 17153 22121 17187
rect 22063 17147 22121 17153
rect 22830 17144 22836 17196
rect 22888 17184 22894 17196
rect 23385 17187 23443 17193
rect 23385 17184 23397 17187
rect 22888 17156 23397 17184
rect 22888 17144 22894 17156
rect 23385 17153 23397 17156
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 24320 17193 24348 17224
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17153 24363 17187
rect 24305 17147 24363 17153
rect 21551 17088 21772 17116
rect 21818 17076 21824 17128
rect 21876 17076 21882 17128
rect 20548 17020 21220 17048
rect 21450 17008 21456 17060
rect 21508 17048 21514 17060
rect 21508 17020 21956 17048
rect 21508 17008 21514 17020
rect 15212 16952 15884 16980
rect 16206 16940 16212 16992
rect 16264 16940 16270 16992
rect 17678 16940 17684 16992
rect 17736 16940 17742 16992
rect 20162 16940 20168 16992
rect 20220 16940 20226 16992
rect 20533 16983 20591 16989
rect 20533 16949 20545 16983
rect 20579 16980 20591 16983
rect 20714 16980 20720 16992
rect 20579 16952 20720 16980
rect 20579 16949 20591 16952
rect 20533 16943 20591 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 21542 16940 21548 16992
rect 21600 16940 21606 16992
rect 21928 16980 21956 17020
rect 22833 16983 22891 16989
rect 22833 16980 22845 16983
rect 21928 16952 22845 16980
rect 22833 16949 22845 16952
rect 22879 16949 22891 16983
rect 22833 16943 22891 16949
rect 24118 16940 24124 16992
rect 24176 16940 24182 16992
rect 24394 16940 24400 16992
rect 24452 16940 24458 16992
rect 1104 16890 24840 16912
rect 1104 16838 3917 16890
rect 3969 16838 3981 16890
rect 4033 16838 4045 16890
rect 4097 16838 4109 16890
rect 4161 16838 4173 16890
rect 4225 16838 9851 16890
rect 9903 16838 9915 16890
rect 9967 16838 9979 16890
rect 10031 16838 10043 16890
rect 10095 16838 10107 16890
rect 10159 16838 15785 16890
rect 15837 16838 15849 16890
rect 15901 16838 15913 16890
rect 15965 16838 15977 16890
rect 16029 16838 16041 16890
rect 16093 16838 21719 16890
rect 21771 16838 21783 16890
rect 21835 16838 21847 16890
rect 21899 16838 21911 16890
rect 21963 16838 21975 16890
rect 22027 16838 24840 16890
rect 1104 16816 24840 16838
rect 1026 16736 1032 16788
rect 1084 16776 1090 16788
rect 1949 16779 2007 16785
rect 1949 16776 1961 16779
rect 1084 16748 1961 16776
rect 1084 16736 1090 16748
rect 1949 16745 1961 16748
rect 1995 16745 2007 16779
rect 1949 16739 2007 16745
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3973 16779 4031 16785
rect 3973 16776 3985 16779
rect 3384 16748 3985 16776
rect 3384 16736 3390 16748
rect 3973 16745 3985 16748
rect 4019 16745 4031 16779
rect 3973 16739 4031 16745
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 4856 16748 8769 16776
rect 4856 16736 4862 16748
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 15565 16779 15623 16785
rect 8757 16739 8815 16745
rect 12636 16748 13308 16776
rect 5994 16708 6000 16720
rect 492 16680 6000 16708
rect 492 16652 520 16680
rect 5994 16668 6000 16680
rect 6052 16708 6058 16720
rect 6052 16680 7696 16708
rect 6052 16668 6058 16680
rect 474 16600 480 16652
rect 532 16600 538 16652
rect 2424 16612 3372 16640
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 2424 16581 2452 16612
rect 3344 16584 3372 16612
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 7466 16640 7472 16652
rect 6972 16612 7472 16640
rect 6972 16600 6978 16612
rect 7466 16600 7472 16612
rect 7524 16600 7530 16652
rect 7558 16600 7564 16652
rect 7616 16600 7622 16652
rect 7668 16640 7696 16680
rect 9766 16668 9772 16720
rect 9824 16708 9830 16720
rect 11054 16708 11060 16720
rect 9824 16680 11060 16708
rect 9824 16668 9830 16680
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 7954 16643 8012 16649
rect 7954 16640 7966 16643
rect 7668 16612 7966 16640
rect 7954 16609 7966 16612
rect 8000 16609 8012 16643
rect 7954 16603 8012 16609
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16640 8171 16643
rect 8478 16640 8484 16652
rect 8159 16612 8484 16640
rect 8159 16609 8171 16612
rect 8113 16603 8171 16609
rect 8478 16600 8484 16612
rect 8536 16600 8542 16652
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 12636 16649 12664 16748
rect 12621 16643 12679 16649
rect 12621 16640 12633 16643
rect 11296 16612 12633 16640
rect 11296 16600 11302 16612
rect 12621 16609 12633 16612
rect 12667 16609 12679 16643
rect 12621 16603 12679 16609
rect 13280 16584 13308 16748
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 16114 16776 16120 16788
rect 15611 16748 16120 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 16114 16736 16120 16748
rect 16172 16736 16178 16788
rect 16206 16736 16212 16788
rect 16264 16776 16270 16788
rect 16264 16748 16436 16776
rect 16264 16736 16270 16748
rect 16408 16717 16436 16748
rect 17678 16736 17684 16788
rect 17736 16736 17742 16788
rect 19886 16736 19892 16788
rect 19944 16736 19950 16788
rect 20162 16736 20168 16788
rect 20220 16776 20226 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20220 16748 21281 16776
rect 20220 16736 20226 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 21450 16736 21456 16788
rect 21508 16736 21514 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 21600 16748 22140 16776
rect 21600 16736 21606 16748
rect 13633 16711 13691 16717
rect 13633 16677 13645 16711
rect 13679 16677 13691 16711
rect 13633 16671 13691 16677
rect 16393 16711 16451 16717
rect 16393 16677 16405 16711
rect 16439 16677 16451 16711
rect 16393 16671 16451 16677
rect 13648 16640 13676 16671
rect 13648 16612 14122 16640
rect 15562 16600 15568 16652
rect 15620 16640 15626 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15620 16612 15761 16640
rect 15620 16600 15626 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 15930 16600 15936 16652
rect 15988 16600 15994 16652
rect 16022 16600 16028 16652
rect 16080 16640 16086 16652
rect 16758 16640 16764 16652
rect 16816 16649 16822 16652
rect 16816 16643 16844 16649
rect 16080 16612 16764 16640
rect 16080 16600 16086 16612
rect 16758 16600 16764 16612
rect 16832 16609 16844 16643
rect 16816 16603 16844 16609
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 17696 16640 17724 16736
rect 19904 16708 19932 16736
rect 19812 16680 19932 16708
rect 21468 16708 21496 16736
rect 21468 16680 21588 16708
rect 19812 16649 19840 16680
rect 16991 16612 17724 16640
rect 19797 16643 19855 16649
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 16816 16600 16822 16603
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 21266 16640 21272 16652
rect 20588 16612 21272 16640
rect 20588 16600 20594 16612
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21450 16600 21456 16652
rect 21508 16600 21514 16652
rect 2409 16575 2467 16581
rect 1872 16544 2360 16572
rect 1872 16513 1900 16544
rect 1857 16507 1915 16513
rect 1857 16473 1869 16507
rect 1903 16473 1915 16507
rect 1857 16467 1915 16473
rect 2130 16464 2136 16516
rect 2188 16464 2194 16516
rect 2332 16504 2360 16544
rect 2409 16541 2421 16575
rect 2455 16541 2467 16575
rect 2409 16535 2467 16541
rect 2884 16544 3280 16572
rect 2884 16504 2912 16544
rect 2332 16476 2912 16504
rect 2958 16464 2964 16516
rect 3016 16464 3022 16516
rect 3252 16504 3280 16544
rect 3326 16532 3332 16584
rect 3384 16532 3390 16584
rect 3602 16532 3608 16584
rect 3660 16532 3666 16584
rect 7101 16575 7159 16581
rect 3712 16544 6316 16572
rect 3712 16504 3740 16544
rect 3252 16476 3740 16504
rect 3786 16464 3792 16516
rect 3844 16504 3850 16516
rect 3881 16507 3939 16513
rect 3881 16504 3893 16507
rect 3844 16476 3893 16504
rect 3844 16464 3850 16476
rect 3881 16473 3893 16476
rect 3927 16473 3939 16507
rect 3881 16467 3939 16473
rect 1581 16439 1639 16445
rect 1581 16405 1593 16439
rect 1627 16436 1639 16439
rect 2148 16436 2176 16464
rect 1627 16408 2176 16436
rect 1627 16405 1639 16408
rect 1581 16399 1639 16405
rect 2682 16396 2688 16448
rect 2740 16396 2746 16448
rect 3050 16396 3056 16448
rect 3108 16396 3114 16448
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3384 16408 3433 16436
rect 3384 16396 3390 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 5534 16436 5540 16448
rect 4304 16408 5540 16436
rect 4304 16396 4310 16408
rect 5534 16396 5540 16408
rect 5592 16396 5598 16448
rect 6288 16436 6316 16544
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7282 16572 7288 16584
rect 7147 16544 7288 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7834 16532 7840 16584
rect 7892 16532 7898 16584
rect 12526 16572 12532 16584
rect 12268 16544 12532 16572
rect 12268 16516 12296 16544
rect 12526 16532 12532 16544
rect 12584 16572 12590 16584
rect 12863 16575 12921 16581
rect 12863 16572 12875 16575
rect 12584 16544 12875 16572
rect 12584 16532 12590 16544
rect 12863 16541 12875 16544
rect 12909 16541 12921 16575
rect 12863 16535 12921 16541
rect 13262 16532 13268 16584
rect 13320 16532 13326 16584
rect 14458 16532 14464 16584
rect 14516 16572 14522 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14516 16544 14565 16572
rect 14516 16532 14522 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16572 15071 16575
rect 15059 16544 15976 16572
rect 15059 16541 15071 16544
rect 15013 16535 15071 16541
rect 15948 16516 15976 16544
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 17589 16575 17647 16581
rect 17589 16541 17601 16575
rect 17635 16572 17647 16575
rect 17681 16575 17739 16581
rect 17681 16572 17693 16575
rect 17635 16544 17693 16572
rect 17635 16541 17647 16544
rect 17589 16535 17647 16541
rect 17681 16541 17693 16544
rect 17727 16541 17739 16575
rect 17681 16535 17739 16541
rect 17862 16532 17868 16584
rect 17920 16572 17926 16584
rect 18598 16572 18604 16584
rect 17920 16544 18604 16572
rect 17920 16532 17926 16544
rect 18598 16532 18604 16544
rect 18656 16572 18662 16584
rect 21177 16575 21235 16581
rect 18656 16565 20098 16572
rect 18656 16544 20051 16565
rect 18656 16532 18662 16544
rect 20039 16531 20051 16544
rect 20085 16534 20098 16565
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 21560 16572 21588 16680
rect 21634 16668 21640 16720
rect 21692 16708 21698 16720
rect 22005 16711 22063 16717
rect 22005 16708 22017 16711
rect 21692 16680 22017 16708
rect 21692 16668 21698 16680
rect 22005 16677 22017 16680
rect 22051 16677 22063 16711
rect 22005 16671 22063 16677
rect 22112 16640 22140 16748
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 22112 16612 22201 16640
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 22189 16603 22247 16609
rect 22296 16612 23704 16640
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21560 16544 21925 16572
rect 21177 16535 21235 16541
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 22296 16572 22324 16612
rect 21913 16535 21971 16541
rect 22204 16544 22324 16572
rect 20085 16531 20097 16534
rect 20039 16525 20097 16531
rect 12250 16464 12256 16516
rect 12308 16464 12314 16516
rect 12406 16476 14596 16504
rect 12406 16436 12434 16476
rect 6288 16408 12434 16436
rect 14090 16396 14096 16448
rect 14148 16436 14154 16448
rect 14277 16439 14335 16445
rect 14277 16436 14289 16439
rect 14148 16408 14289 16436
rect 14148 16396 14154 16408
rect 14277 16405 14289 16408
rect 14323 16405 14335 16439
rect 14568 16436 14596 16476
rect 14642 16464 14648 16516
rect 14700 16464 14706 16516
rect 15120 16476 15700 16504
rect 15120 16436 15148 16476
rect 14568 16408 15148 16436
rect 14277 16399 14335 16405
rect 15378 16396 15384 16448
rect 15436 16396 15442 16448
rect 15672 16436 15700 16476
rect 15930 16464 15936 16516
rect 15988 16464 15994 16516
rect 17865 16439 17923 16445
rect 17865 16436 17877 16439
rect 15672 16408 17877 16436
rect 17865 16405 17877 16408
rect 17911 16405 17923 16439
rect 17865 16399 17923 16405
rect 20809 16439 20867 16445
rect 20809 16405 20821 16439
rect 20855 16436 20867 16439
rect 20990 16436 20996 16448
rect 20855 16408 20996 16436
rect 20855 16405 20867 16408
rect 20809 16399 20867 16405
rect 20990 16396 20996 16408
rect 21048 16436 21054 16448
rect 21192 16436 21220 16535
rect 22204 16513 22232 16544
rect 22922 16532 22928 16584
rect 22980 16532 22986 16584
rect 23477 16575 23535 16581
rect 23477 16541 23489 16575
rect 23523 16572 23535 16575
rect 23566 16572 23572 16584
rect 23523 16544 23572 16572
rect 23523 16541 23535 16544
rect 23477 16535 23535 16541
rect 23566 16532 23572 16544
rect 23624 16532 23630 16584
rect 23676 16581 23704 16612
rect 23934 16600 23940 16652
rect 23992 16600 23998 16652
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16541 23719 16575
rect 23661 16535 23719 16541
rect 22189 16507 22247 16513
rect 22189 16473 22201 16507
rect 22235 16473 22247 16507
rect 22189 16467 22247 16473
rect 21048 16408 21220 16436
rect 21453 16439 21511 16445
rect 21048 16396 21054 16408
rect 21453 16405 21465 16439
rect 21499 16436 21511 16439
rect 21634 16436 21640 16448
rect 21499 16408 21640 16436
rect 21499 16405 21511 16408
rect 21453 16399 21511 16405
rect 21634 16396 21640 16408
rect 21692 16396 21698 16448
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22554 16436 22560 16448
rect 22152 16408 22560 16436
rect 22152 16396 22158 16408
rect 22554 16396 22560 16408
rect 22612 16396 22618 16448
rect 22940 16436 22968 16532
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22940 16408 23305 16436
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 1104 16346 25000 16368
rect 1104 16294 6884 16346
rect 6936 16294 6948 16346
rect 7000 16294 7012 16346
rect 7064 16294 7076 16346
rect 7128 16294 7140 16346
rect 7192 16294 12818 16346
rect 12870 16294 12882 16346
rect 12934 16294 12946 16346
rect 12998 16294 13010 16346
rect 13062 16294 13074 16346
rect 13126 16294 18752 16346
rect 18804 16294 18816 16346
rect 18868 16294 18880 16346
rect 18932 16294 18944 16346
rect 18996 16294 19008 16346
rect 19060 16294 24686 16346
rect 24738 16294 24750 16346
rect 24802 16294 24814 16346
rect 24866 16294 24878 16346
rect 24930 16294 24942 16346
rect 24994 16294 25000 16346
rect 1104 16272 25000 16294
rect 1762 16192 1768 16244
rect 1820 16192 1826 16244
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2958 16232 2964 16244
rect 2188 16204 2964 16232
rect 2188 16192 2194 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 3660 16204 5365 16232
rect 3660 16192 3666 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 7576 16204 8156 16232
rect 1673 16167 1731 16173
rect 1673 16133 1685 16167
rect 1719 16164 1731 16167
rect 2038 16164 2044 16176
rect 1719 16136 2044 16164
rect 1719 16133 1731 16136
rect 1673 16127 1731 16133
rect 2038 16124 2044 16136
rect 2096 16124 2102 16176
rect 2222 16124 2228 16176
rect 2280 16124 2286 16176
rect 3326 16164 3332 16176
rect 2424 16136 3332 16164
rect 2424 16135 2452 16136
rect 2391 16129 2452 16135
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2240 16096 2268 16124
rect 2179 16068 2268 16096
rect 2391 16095 2403 16129
rect 2437 16098 2452 16129
rect 3326 16124 3332 16136
rect 3384 16124 3390 16176
rect 2437 16095 2449 16098
rect 2391 16089 2449 16095
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2148 15892 2176 16059
rect 2774 16056 2780 16108
rect 2832 16096 2838 16108
rect 3513 16099 3571 16105
rect 3513 16096 3525 16099
rect 2832 16068 3525 16096
rect 2832 16056 2838 16068
rect 3513 16065 3525 16068
rect 3559 16065 3571 16099
rect 3513 16059 3571 16065
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 4522 16056 4528 16108
rect 4580 16105 4586 16108
rect 4580 16099 4608 16105
rect 4596 16065 4608 16099
rect 7576 16096 7604 16204
rect 4580 16059 4608 16065
rect 7484 16068 7604 16096
rect 7727 16099 7785 16105
rect 4580 16056 4586 16059
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 3694 16028 3700 16040
rect 3016 16000 3700 16028
rect 3016 15988 3022 16000
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 4706 15988 4712 16040
rect 4764 15988 4770 16040
rect 4890 15988 4896 16040
rect 4948 16028 4954 16040
rect 7006 16028 7012 16040
rect 4948 16000 7012 16028
rect 4948 15988 4954 16000
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7484 16037 7512 16068
rect 7727 16065 7739 16099
rect 7773 16096 7785 16099
rect 7834 16096 7840 16108
rect 7773 16068 7840 16096
rect 7773 16065 7785 16068
rect 7727 16059 7785 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 8128 16096 8156 16204
rect 8386 16192 8392 16244
rect 8444 16192 8450 16244
rect 8478 16192 8484 16244
rect 8536 16192 8542 16244
rect 8956 16204 12354 16232
rect 8404 16164 8432 16192
rect 8956 16164 8984 16204
rect 8404 16136 8984 16164
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 9088 16136 10732 16164
rect 9088 16124 9094 16136
rect 8662 16096 8668 16108
rect 8128 16068 8668 16096
rect 8662 16056 8668 16068
rect 8720 16096 8726 16108
rect 8849 16099 8907 16105
rect 8849 16096 8861 16099
rect 8720 16068 8861 16096
rect 8720 16056 8726 16068
rect 8849 16065 8861 16068
rect 8895 16065 8907 16099
rect 8849 16059 8907 16065
rect 9123 16099 9181 16105
rect 9123 16065 9135 16099
rect 9169 16096 9181 16099
rect 9766 16096 9772 16108
rect 9169 16068 9772 16096
rect 9169 16065 9181 16068
rect 9123 16059 9181 16065
rect 9766 16056 9772 16068
rect 9824 16056 9830 16108
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 15997 7527 16031
rect 7469 15991 7527 15997
rect 3145 15963 3203 15969
rect 3145 15929 3157 15963
rect 3191 15960 3203 15963
rect 4157 15963 4215 15969
rect 4157 15960 4169 15963
rect 3191 15932 4169 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 4157 15929 4169 15932
rect 4203 15929 4215 15963
rect 4157 15923 4215 15929
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 6638 15960 6644 15972
rect 5500 15932 6644 15960
rect 5500 15920 5506 15932
rect 6638 15920 6644 15932
rect 6696 15920 6702 15972
rect 6822 15920 6828 15972
rect 6880 15960 6886 15972
rect 7484 15960 7512 15991
rect 10413 15963 10471 15969
rect 10413 15960 10425 15963
rect 6880 15932 7512 15960
rect 9508 15932 10425 15960
rect 6880 15920 6886 15932
rect 3694 15892 3700 15904
rect 2148 15864 3700 15892
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 4614 15852 4620 15904
rect 4672 15892 4678 15904
rect 9508 15892 9536 15932
rect 10413 15929 10425 15932
rect 10459 15929 10471 15963
rect 10413 15923 10471 15929
rect 4672 15864 9536 15892
rect 4672 15852 4678 15864
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 9861 15895 9919 15901
rect 9861 15892 9873 15895
rect 9732 15864 9873 15892
rect 9732 15852 9738 15864
rect 9861 15861 9873 15864
rect 9907 15861 9919 15895
rect 10704 15892 10732 16136
rect 12158 16124 12164 16176
rect 12216 16124 12222 16176
rect 12326 16135 12354 16204
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 12768 16204 13093 16232
rect 12768 16192 12774 16204
rect 13081 16201 13093 16204
rect 13127 16201 13139 16235
rect 13081 16195 13139 16201
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 15381 16235 15439 16241
rect 15381 16232 15393 16235
rect 14700 16204 15393 16232
rect 14700 16192 14706 16204
rect 15381 16201 15393 16204
rect 15427 16201 15439 16235
rect 15381 16195 15439 16201
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 17218 16232 17224 16244
rect 15988 16204 17224 16232
rect 15988 16192 15994 16204
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 19245 16235 19303 16241
rect 19245 16201 19257 16235
rect 19291 16201 19303 16235
rect 19245 16195 19303 16201
rect 12326 16129 12385 16135
rect 10778 16056 10784 16108
rect 10836 16096 10842 16108
rect 11238 16096 11244 16108
rect 10836 16068 11244 16096
rect 10836 16056 10842 16068
rect 11238 16056 11244 16068
rect 11296 16096 11302 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 11296 16068 12081 16096
rect 11296 16056 11302 16068
rect 12069 16065 12081 16068
rect 12115 16096 12127 16099
rect 12176 16096 12204 16124
rect 12326 16098 12339 16129
rect 12115 16068 12204 16096
rect 12327 16095 12339 16098
rect 12373 16096 12385 16129
rect 16022 16124 16028 16176
rect 16080 16164 16086 16176
rect 16298 16164 16304 16176
rect 16080 16136 16304 16164
rect 16080 16124 16086 16136
rect 16298 16124 16304 16136
rect 16356 16124 16362 16176
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 18110 16167 18168 16173
rect 18110 16164 18122 16167
rect 18012 16136 18122 16164
rect 18012 16124 18018 16136
rect 18110 16133 18122 16136
rect 18156 16133 18168 16167
rect 19260 16164 19288 16195
rect 20714 16192 20720 16244
rect 20772 16192 20778 16244
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 21450 16232 21456 16244
rect 20855 16204 21456 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 21450 16192 21456 16204
rect 21508 16192 21514 16244
rect 23474 16192 23480 16244
rect 23532 16192 23538 16244
rect 23842 16192 23848 16244
rect 23900 16232 23906 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 23900 16204 24317 16232
rect 23900 16192 23906 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 19260 16136 19840 16164
rect 18110 16127 18168 16133
rect 12710 16096 12716 16108
rect 12373 16095 12716 16096
rect 12327 16089 12716 16095
rect 12342 16068 12716 16089
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 13814 16056 13820 16108
rect 13872 16096 13878 16108
rect 14642 16105 14648 16108
rect 14611 16099 14648 16105
rect 14611 16096 14623 16099
rect 13872 16068 14623 16096
rect 13872 16056 13878 16068
rect 14611 16065 14623 16068
rect 14611 16059 14648 16065
rect 14642 16056 14648 16059
rect 14700 16056 14706 16108
rect 18874 16056 18880 16108
rect 18932 16096 18938 16108
rect 19812 16105 19840 16136
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 18932 16068 19349 16096
rect 18932 16056 18938 16068
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19337 16059 19395 16065
rect 19797 16099 19855 16105
rect 19797 16065 19809 16099
rect 19843 16065 19855 16099
rect 19797 16059 19855 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20732 16096 20760 16192
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20732 16068 20821 16096
rect 20625 16059 20683 16065
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 13262 15988 13268 16040
rect 13320 16028 13326 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 13320 16000 14381 16028
rect 13320 15988 13326 16000
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 17218 15988 17224 16040
rect 17276 16028 17282 16040
rect 17862 16028 17868 16040
rect 17276 16000 17868 16028
rect 17276 15988 17282 16000
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 20640 16028 20668 16059
rect 20990 16056 20996 16108
rect 21048 16056 21054 16108
rect 22891 16099 22949 16105
rect 22891 16096 22903 16099
rect 22066 16068 22903 16096
rect 21008 16028 21036 16056
rect 20640 16000 21036 16028
rect 19794 15920 19800 15972
rect 19852 15960 19858 15972
rect 20990 15960 20996 15972
rect 19852 15932 20996 15960
rect 19852 15920 19858 15932
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 15102 15892 15108 15904
rect 10704 15864 15108 15892
rect 9861 15855 9919 15861
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 19518 15892 19524 15904
rect 19475 15864 19524 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 19613 15895 19671 15901
rect 19613 15861 19625 15895
rect 19659 15892 19671 15895
rect 19978 15892 19984 15904
rect 19659 15864 19984 15892
rect 19659 15861 19671 15864
rect 19613 15855 19671 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 22066 15892 22094 16068
rect 22891 16065 22903 16068
rect 22937 16065 22949 16099
rect 23492 16096 23520 16192
rect 24029 16099 24087 16105
rect 24029 16096 24041 16099
rect 23492 16068 24041 16096
rect 22891 16059 22949 16065
rect 24029 16065 24041 16068
rect 24075 16065 24087 16099
rect 24029 16059 24087 16065
rect 24121 16099 24179 16105
rect 24121 16065 24133 16099
rect 24167 16096 24179 16099
rect 24394 16096 24400 16108
rect 24167 16068 24400 16096
rect 24167 16065 24179 16068
rect 24121 16059 24179 16065
rect 24394 16056 24400 16068
rect 24452 16056 24458 16108
rect 22554 15988 22560 16040
rect 22612 16028 22618 16040
rect 22649 16031 22707 16037
rect 22649 16028 22661 16031
rect 22612 16000 22661 16028
rect 22612 15988 22618 16000
rect 22649 15997 22661 16000
rect 22695 15997 22707 16031
rect 22649 15991 22707 15997
rect 23658 15988 23664 16040
rect 23716 16028 23722 16040
rect 24305 16031 24363 16037
rect 24305 16028 24317 16031
rect 23716 16000 24317 16028
rect 23716 15988 23722 16000
rect 24305 15997 24317 16000
rect 24351 15997 24363 16031
rect 24305 15991 24363 15997
rect 20220 15864 22094 15892
rect 20220 15852 20226 15864
rect 23658 15852 23664 15904
rect 23716 15852 23722 15904
rect 1104 15802 24840 15824
rect 1104 15750 3917 15802
rect 3969 15750 3981 15802
rect 4033 15750 4045 15802
rect 4097 15750 4109 15802
rect 4161 15750 4173 15802
rect 4225 15750 9851 15802
rect 9903 15750 9915 15802
rect 9967 15750 9979 15802
rect 10031 15750 10043 15802
rect 10095 15750 10107 15802
rect 10159 15750 15785 15802
rect 15837 15750 15849 15802
rect 15901 15750 15913 15802
rect 15965 15750 15977 15802
rect 16029 15750 16041 15802
rect 16093 15750 21719 15802
rect 21771 15750 21783 15802
rect 21835 15750 21847 15802
rect 21899 15750 21911 15802
rect 21963 15750 21975 15802
rect 22027 15750 24840 15802
rect 1104 15728 24840 15750
rect 2866 15648 2872 15700
rect 2924 15648 2930 15700
rect 4614 15688 4620 15700
rect 3344 15660 4620 15688
rect 3234 15484 3240 15496
rect 2240 15456 3240 15484
rect 2240 15425 2268 15456
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 1857 15419 1915 15425
rect 1857 15385 1869 15419
rect 1903 15416 1915 15419
rect 2225 15419 2283 15425
rect 2225 15416 2237 15419
rect 1903 15388 2237 15416
rect 1903 15385 1915 15388
rect 1857 15379 1915 15385
rect 2225 15385 2237 15388
rect 2271 15385 2283 15419
rect 2225 15379 2283 15385
rect 2777 15419 2835 15425
rect 2777 15385 2789 15419
rect 2823 15416 2835 15419
rect 3344 15416 3372 15660
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 4801 15691 4859 15697
rect 4801 15688 4813 15691
rect 4764 15660 4813 15688
rect 4764 15648 4770 15660
rect 4801 15657 4813 15660
rect 4847 15657 4859 15691
rect 4801 15651 4859 15657
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7837 15691 7895 15697
rect 7837 15688 7849 15691
rect 7616 15660 7849 15688
rect 7616 15648 7622 15660
rect 7837 15657 7849 15660
rect 7883 15657 7895 15691
rect 7837 15651 7895 15657
rect 9674 15648 9680 15700
rect 9732 15648 9738 15700
rect 10594 15648 10600 15700
rect 10652 15688 10658 15700
rect 10781 15691 10839 15697
rect 10781 15688 10793 15691
rect 10652 15660 10793 15688
rect 10652 15648 10658 15660
rect 10781 15657 10793 15660
rect 10827 15657 10839 15691
rect 10781 15651 10839 15657
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 16758 15688 16764 15700
rect 12400 15660 16764 15688
rect 12400 15648 12406 15660
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 18325 15691 18383 15697
rect 18325 15657 18337 15691
rect 18371 15688 18383 15691
rect 18874 15688 18880 15700
rect 18371 15660 18880 15688
rect 18371 15657 18383 15660
rect 18325 15651 18383 15657
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 23842 15688 23848 15700
rect 19352 15660 19932 15688
rect 9585 15623 9643 15629
rect 9585 15589 9597 15623
rect 9631 15620 9643 15623
rect 9692 15620 9720 15648
rect 19352 15620 19380 15660
rect 9631 15592 9720 15620
rect 18248 15592 19380 15620
rect 9631 15589 9643 15592
rect 9585 15583 9643 15589
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 3789 15555 3847 15561
rect 3789 15552 3801 15555
rect 3752 15524 3801 15552
rect 3752 15512 3758 15524
rect 3789 15521 3801 15524
rect 3835 15521 3847 15555
rect 3789 15515 3847 15521
rect 5442 15512 5448 15564
rect 5500 15512 5506 15564
rect 6362 15512 6368 15564
rect 6420 15552 6426 15564
rect 6822 15552 6828 15564
rect 6420 15524 6828 15552
rect 6420 15512 6426 15524
rect 6822 15512 6828 15524
rect 6880 15512 6886 15564
rect 8941 15555 8999 15561
rect 8941 15521 8953 15555
rect 8987 15552 8999 15555
rect 9030 15552 9036 15564
rect 8987 15524 9036 15552
rect 8987 15521 8999 15524
rect 8941 15515 8999 15521
rect 9030 15512 9036 15524
rect 9088 15552 9094 15564
rect 9306 15552 9312 15564
rect 9088 15524 9312 15552
rect 9088 15512 9094 15524
rect 9306 15512 9312 15524
rect 9364 15512 9370 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9978 15555 10036 15561
rect 9978 15552 9990 15555
rect 9732 15524 9990 15552
rect 9732 15512 9738 15524
rect 9978 15521 9990 15524
rect 10024 15521 10036 15555
rect 9978 15515 10036 15521
rect 13354 15512 13360 15564
rect 13412 15552 13418 15564
rect 18248 15552 18276 15592
rect 13412 15524 18276 15552
rect 13412 15512 13418 15524
rect 19904 15496 19932 15660
rect 21652 15660 23848 15688
rect 21652 15632 21680 15660
rect 23842 15648 23848 15660
rect 23900 15648 23906 15700
rect 24118 15648 24124 15700
rect 24176 15648 24182 15700
rect 21634 15580 21640 15632
rect 21692 15580 21698 15632
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 21192 15524 22385 15552
rect 21192 15496 21220 15524
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 22373 15515 22431 15521
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 2823 15388 3372 15416
rect 3436 15416 3464 15447
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 4031 15487 4089 15493
rect 4031 15484 4043 15487
rect 3568 15456 4043 15484
rect 3568 15444 3574 15456
rect 4031 15453 4043 15456
rect 4077 15453 4089 15487
rect 4031 15447 4089 15453
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 5350 15484 5356 15496
rect 4212 15456 5356 15484
rect 4212 15444 4218 15456
rect 5350 15444 5356 15456
rect 5408 15484 5414 15496
rect 5687 15487 5745 15493
rect 5687 15484 5699 15487
rect 5408 15456 5699 15484
rect 5408 15444 5414 15456
rect 5687 15453 5699 15456
rect 5733 15453 5745 15487
rect 5687 15447 5745 15453
rect 6196 15456 6682 15484
rect 6196 15416 6224 15456
rect 3436 15388 6224 15416
rect 2823 15385 2835 15388
rect 2777 15379 2835 15385
rect 2314 15308 2320 15360
rect 2372 15308 2378 15360
rect 3234 15308 3240 15360
rect 3292 15308 3298 15360
rect 3694 15308 3700 15360
rect 3752 15348 3758 15360
rect 6362 15348 6368 15360
rect 3752 15320 6368 15348
rect 3752 15308 3758 15320
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6457 15351 6515 15357
rect 6457 15317 6469 15351
rect 6503 15348 6515 15351
rect 6546 15348 6552 15360
rect 6503 15320 6552 15348
rect 6503 15317 6515 15320
rect 6457 15311 6515 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 6654 15348 6682 15456
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7099 15487 7157 15493
rect 7099 15484 7111 15487
rect 7064 15456 7111 15484
rect 7064 15444 7070 15456
rect 7099 15453 7111 15456
rect 7145 15453 7157 15487
rect 7099 15447 7157 15453
rect 9122 15444 9128 15496
rect 9180 15444 9186 15496
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 11147 15487 11205 15493
rect 11147 15453 11159 15487
rect 11193 15484 11205 15487
rect 11193 15456 11560 15484
rect 11193 15453 11205 15456
rect 11147 15447 11205 15453
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7742 15416 7748 15428
rect 7432 15388 7748 15416
rect 7432 15376 7438 15388
rect 7742 15376 7748 15388
rect 7800 15376 7806 15428
rect 10888 15416 10916 15447
rect 11238 15416 11244 15428
rect 10888 15388 11244 15416
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 11422 15376 11428 15428
rect 11480 15416 11486 15428
rect 11532 15416 11560 15456
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 16850 15484 16856 15496
rect 11664 15456 16856 15484
rect 11664 15444 11670 15456
rect 16850 15444 16856 15456
rect 16908 15444 16914 15496
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18012 15456 18521 15484
rect 18012 15444 18018 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19352 15477 19546 15484
rect 19352 15456 19499 15477
rect 11698 15416 11704 15428
rect 11480 15388 11704 15416
rect 11480 15376 11486 15388
rect 11698 15376 11704 15388
rect 11756 15416 11762 15428
rect 14090 15416 14096 15428
rect 11756 15388 14096 15416
rect 11756 15376 11762 15388
rect 14090 15376 14096 15388
rect 14148 15376 14154 15428
rect 19260 15416 19288 15447
rect 19352 15428 19380 15456
rect 19487 15443 19499 15456
rect 19533 15446 19546 15477
rect 19533 15443 19545 15446
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 20162 15484 20168 15496
rect 19944 15456 20168 15484
rect 19944 15444 19950 15456
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 21174 15444 21180 15496
rect 21232 15444 21238 15496
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22281 15487 22339 15493
rect 22281 15484 22293 15487
rect 22244 15456 22293 15484
rect 22244 15444 22250 15456
rect 22281 15453 22293 15456
rect 22327 15453 22339 15487
rect 22281 15447 22339 15453
rect 19487 15437 19545 15443
rect 17972 15388 19288 15416
rect 17972 15360 18000 15388
rect 19334 15376 19340 15428
rect 19392 15376 19398 15428
rect 22296 15416 22324 15447
rect 22462 15444 22468 15496
rect 22520 15484 22526 15496
rect 23937 15487 23995 15493
rect 23937 15484 23949 15487
rect 22520 15456 23949 15484
rect 22520 15444 22526 15456
rect 23937 15453 23949 15456
rect 23983 15453 23995 15487
rect 23937 15447 23995 15453
rect 22618 15419 22676 15425
rect 22618 15416 22630 15419
rect 22296 15388 22630 15416
rect 22618 15385 22630 15388
rect 22664 15385 22676 15419
rect 22618 15379 22676 15385
rect 10962 15348 10968 15360
rect 6654 15320 10968 15348
rect 10962 15308 10968 15320
rect 11020 15308 11026 15360
rect 11882 15308 11888 15360
rect 11940 15308 11946 15360
rect 13538 15308 13544 15360
rect 13596 15348 13602 15360
rect 15286 15348 15292 15360
rect 13596 15320 15292 15348
rect 13596 15308 13602 15320
rect 15286 15308 15292 15320
rect 15344 15308 15350 15360
rect 17954 15308 17960 15360
rect 18012 15308 18018 15360
rect 19794 15308 19800 15360
rect 19852 15348 19858 15360
rect 20257 15351 20315 15357
rect 20257 15348 20269 15351
rect 19852 15320 20269 15348
rect 19852 15308 19858 15320
rect 20257 15317 20269 15320
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 22097 15351 22155 15357
rect 22097 15317 22109 15351
rect 22143 15348 22155 15351
rect 22738 15348 22744 15360
rect 22143 15320 22744 15348
rect 22143 15317 22155 15320
rect 22097 15311 22155 15317
rect 22738 15308 22744 15320
rect 22796 15308 22802 15360
rect 23750 15308 23756 15360
rect 23808 15308 23814 15360
rect 1104 15258 25000 15280
rect 1104 15206 6884 15258
rect 6936 15206 6948 15258
rect 7000 15206 7012 15258
rect 7064 15206 7076 15258
rect 7128 15206 7140 15258
rect 7192 15206 12818 15258
rect 12870 15206 12882 15258
rect 12934 15206 12946 15258
rect 12998 15206 13010 15258
rect 13062 15206 13074 15258
rect 13126 15206 18752 15258
rect 18804 15206 18816 15258
rect 18868 15206 18880 15258
rect 18932 15206 18944 15258
rect 18996 15206 19008 15258
rect 19060 15206 24686 15258
rect 24738 15206 24750 15258
rect 24802 15206 24814 15258
rect 24866 15206 24878 15258
rect 24930 15206 24942 15258
rect 24994 15206 25000 15258
rect 1104 15184 25000 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 2130 15144 2136 15156
rect 1627 15116 2136 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 2130 15104 2136 15116
rect 2188 15104 2194 15156
rect 2746 15116 4384 15144
rect 2314 15076 2320 15088
rect 1872 15048 2320 15076
rect 1872 15020 1900 15048
rect 2314 15036 2320 15048
rect 2372 15076 2378 15088
rect 2746 15076 2774 15116
rect 2372 15048 2774 15076
rect 2372 15036 2378 15048
rect 3142 15036 3148 15088
rect 3200 15036 3206 15088
rect 3234 15036 3240 15088
rect 3292 15076 3298 15088
rect 3329 15079 3387 15085
rect 3329 15076 3341 15079
rect 3292 15048 3341 15076
rect 3292 15036 3298 15048
rect 3329 15045 3341 15048
rect 3375 15045 3387 15079
rect 3329 15039 3387 15045
rect 4154 15036 4160 15088
rect 4212 15036 4218 15088
rect 1762 14968 1768 15020
rect 1820 14968 1826 15020
rect 1854 14968 1860 15020
rect 1912 14968 1918 15020
rect 2131 15011 2189 15017
rect 2131 14977 2143 15011
rect 2177 15008 2189 15011
rect 3160 15008 3188 15036
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 2177 14980 3096 15008
rect 3160 14980 3893 15008
rect 2177 14977 2189 14980
rect 2131 14971 2189 14977
rect 3068 14940 3096 14980
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 3881 14971 3939 14977
rect 4172 14940 4200 15036
rect 4356 15017 4384 15116
rect 4614 15104 4620 15156
rect 4672 15104 4678 15156
rect 7282 15144 7288 15156
rect 6564 15116 7288 15144
rect 4632 15047 4660 15104
rect 6564 15076 6592 15116
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 9950 15144 9956 15156
rect 8904 15116 9956 15144
rect 8904 15104 8910 15116
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10229 15147 10287 15153
rect 10229 15144 10241 15147
rect 10192 15116 10241 15144
rect 10192 15104 10198 15116
rect 10229 15113 10241 15116
rect 10275 15113 10287 15147
rect 10229 15107 10287 15113
rect 10334 15116 12296 15144
rect 4599 15041 4660 15047
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 14977 4399 15011
rect 4599 15007 4611 15041
rect 4645 15010 4660 15041
rect 5000 15048 6592 15076
rect 5000 15020 5028 15048
rect 4645 15007 4657 15010
rect 4599 15001 4657 15007
rect 4341 14971 4399 14977
rect 4982 14968 4988 15020
rect 5040 14968 5046 15020
rect 6564 15017 6592 15048
rect 9306 15036 9312 15088
rect 9364 15036 9370 15088
rect 9674 15036 9680 15088
rect 9732 15076 9738 15088
rect 10334 15076 10362 15116
rect 9732 15048 10362 15076
rect 11701 15079 11759 15085
rect 9732 15036 9738 15048
rect 11701 15045 11713 15079
rect 11747 15076 11759 15079
rect 11790 15076 11796 15088
rect 11747 15048 11796 15076
rect 11747 15045 11759 15048
rect 11701 15039 11759 15045
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 12268 15076 12296 15116
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12805 15147 12863 15153
rect 12805 15144 12817 15147
rect 12676 15116 12817 15144
rect 12676 15104 12682 15116
rect 12805 15113 12817 15116
rect 12851 15113 12863 15147
rect 12805 15107 12863 15113
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13170 15144 13176 15156
rect 13035 15116 13176 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13004 15076 13032 15107
rect 13170 15104 13176 15116
rect 13228 15144 13234 15156
rect 13538 15144 13544 15156
rect 13228 15116 13544 15144
rect 13228 15104 13234 15116
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 14642 15104 14648 15156
rect 14700 15144 14706 15156
rect 16390 15144 16396 15156
rect 14700 15116 16396 15144
rect 14700 15104 14706 15116
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 17586 15144 17592 15156
rect 16500 15116 17592 15144
rect 12023 15048 12204 15076
rect 12268 15048 13032 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 7466 15017 7472 15020
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 7423 15011 7472 15017
rect 7423 14977 7435 15011
rect 7469 14977 7472 15011
rect 7423 14971 7472 14977
rect 7466 14968 7472 14971
rect 7524 14968 7530 15020
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 9324 15008 9352 15036
rect 9491 15011 9549 15017
rect 9491 15008 9503 15011
rect 9324 14980 9503 15008
rect 9491 14977 9503 14980
rect 9537 15008 9549 15011
rect 10226 15008 10232 15020
rect 9537 14980 10232 15008
rect 9537 14977 9549 14980
rect 9491 14971 9549 14977
rect 10226 14968 10232 14980
rect 10284 15008 10290 15020
rect 10870 15008 10876 15020
rect 10284 14980 10876 15008
rect 10284 14968 10290 14980
rect 10870 14968 10876 14980
rect 10928 14968 10934 15020
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 12176 15008 12204 15048
rect 14183 15021 14241 15027
rect 12342 15008 12348 15020
rect 12176 14980 12348 15008
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 15008 12495 15011
rect 13722 15008 13728 15020
rect 12483 14980 13728 15008
rect 12483 14977 12495 14980
rect 12437 14971 12495 14977
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 14090 14968 14096 15020
rect 14148 15008 14154 15020
rect 14183 15008 14195 15021
rect 14148 14987 14195 15008
rect 14229 15008 14241 15021
rect 16500 15008 16528 15116
rect 17586 15104 17592 15116
rect 17644 15144 17650 15156
rect 19334 15144 19340 15156
rect 17644 15116 19340 15144
rect 17644 15104 17650 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 22462 15144 22468 15156
rect 19751 15116 22468 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22738 15104 22744 15156
rect 22796 15104 22802 15156
rect 24210 15144 24216 15156
rect 23768 15116 24216 15144
rect 17218 15076 17224 15088
rect 17144 15048 17224 15076
rect 17144 15017 17172 15048
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 17396 15079 17454 15085
rect 17396 15045 17408 15079
rect 17442 15076 17454 15079
rect 17770 15076 17776 15088
rect 17442 15048 17776 15076
rect 17442 15045 17454 15048
rect 17396 15039 17454 15045
rect 17770 15036 17776 15048
rect 17828 15036 17834 15088
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 19610 15076 19616 15088
rect 17920 15048 19616 15076
rect 17920 15036 17926 15048
rect 19610 15036 19616 15048
rect 19668 15076 19674 15088
rect 21174 15076 21180 15088
rect 19668 15048 21180 15076
rect 19668 15036 19674 15048
rect 14229 14987 16528 15008
rect 14148 14980 16528 14987
rect 17129 15011 17187 15017
rect 14148 14968 14154 14980
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 18506 14968 18512 15020
rect 18564 14968 18570 15020
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 6362 14940 6368 14952
rect 3068 14912 4200 14940
rect 5000 14912 6368 14940
rect 2746 14844 4108 14872
rect 1302 14764 1308 14816
rect 1360 14804 1366 14816
rect 2746 14804 2774 14844
rect 1360 14776 2774 14804
rect 1360 14764 1366 14776
rect 2866 14764 2872 14816
rect 2924 14764 2930 14816
rect 3050 14764 3056 14816
rect 3108 14804 3114 14816
rect 3421 14807 3479 14813
rect 3421 14804 3433 14807
rect 3108 14776 3433 14804
rect 3108 14764 3114 14776
rect 3421 14773 3433 14776
rect 3467 14773 3479 14807
rect 3421 14767 3479 14773
rect 3970 14764 3976 14816
rect 4028 14764 4034 14816
rect 4080 14804 4108 14844
rect 4798 14804 4804 14816
rect 4080 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14804 4862 14816
rect 5000 14804 5028 14912
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 6914 14900 6920 14952
rect 6972 14940 6978 14952
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6972 14912 7021 14940
rect 6972 14900 6978 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 7009 14903 7067 14909
rect 7114 14912 7297 14940
rect 5074 14832 5080 14884
rect 5132 14872 5138 14884
rect 5132 14844 5488 14872
rect 5132 14832 5138 14844
rect 4856 14776 5028 14804
rect 4856 14764 4862 14776
rect 5350 14764 5356 14816
rect 5408 14764 5414 14816
rect 5460 14804 5488 14844
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 7114 14872 7142 14912
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 8680 14940 8708 14968
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 7800 14912 9229 14940
rect 7800 14900 7806 14912
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 11882 14900 11888 14952
rect 11940 14900 11946 14952
rect 13906 14900 13912 14952
rect 13964 14900 13970 14952
rect 5960 14844 7142 14872
rect 18524 14872 18552 14968
rect 19444 14940 19472 14971
rect 19518 14968 19524 15020
rect 19576 14968 19582 15020
rect 19794 15008 19800 15020
rect 19628 14980 19800 15008
rect 19628 14940 19656 14980
rect 19794 14968 19800 14980
rect 19852 14968 19858 15020
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 20272 15017 20300 15048
rect 21174 15036 21180 15048
rect 21232 15036 21238 15088
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20513 15011 20571 15017
rect 20513 15008 20525 15011
rect 20257 14971 20315 14977
rect 20364 14980 20525 15008
rect 19444 14912 19656 14940
rect 19705 14943 19763 14949
rect 19705 14909 19717 14943
rect 19751 14940 19763 14943
rect 19889 14943 19947 14949
rect 19889 14940 19901 14943
rect 19751 14912 19901 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 19889 14909 19901 14912
rect 19935 14909 19947 14943
rect 20364 14940 20392 14980
rect 20513 14977 20525 14980
rect 20559 14977 20571 15011
rect 20513 14971 20571 14977
rect 20806 14968 20812 15020
rect 20864 15008 20870 15020
rect 22063 15011 22121 15017
rect 22063 15008 22075 15011
rect 20864 14980 22075 15008
rect 20864 14968 20870 14980
rect 22063 14977 22075 14980
rect 22109 14977 22121 15011
rect 22756 15008 22784 15104
rect 23768 15085 23796 15116
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 23753 15079 23811 15085
rect 23753 15045 23765 15079
rect 23799 15045 23811 15079
rect 23753 15039 23811 15045
rect 23385 15011 23443 15017
rect 23385 15008 23397 15011
rect 22756 14980 23397 15008
rect 22063 14971 22121 14977
rect 23385 14977 23397 14980
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 24210 15008 24216 15020
rect 23716 14980 24216 15008
rect 23716 14968 23722 14980
rect 24210 14968 24216 14980
rect 24268 14968 24274 15020
rect 19889 14903 19947 14909
rect 20272 14912 20392 14940
rect 20272 14884 20300 14912
rect 21266 14900 21272 14952
rect 21324 14940 21330 14952
rect 21542 14940 21548 14952
rect 21324 14912 21548 14940
rect 21324 14900 21330 14912
rect 21542 14900 21548 14912
rect 21600 14940 21606 14952
rect 21821 14943 21879 14949
rect 21821 14940 21833 14943
rect 21600 14912 21833 14940
rect 21600 14900 21606 14912
rect 21821 14909 21833 14912
rect 21867 14909 21879 14943
rect 21821 14903 21879 14909
rect 22830 14900 22836 14952
rect 22888 14940 22894 14952
rect 24489 14943 24547 14949
rect 24489 14940 24501 14943
rect 22888 14912 24501 14940
rect 22888 14900 22894 14912
rect 24489 14909 24501 14912
rect 24535 14909 24547 14943
rect 24489 14903 24547 14909
rect 20254 14872 20260 14884
rect 18524 14844 20260 14872
rect 5960 14832 5966 14844
rect 20254 14832 20260 14844
rect 20312 14832 20318 14884
rect 23477 14875 23535 14881
rect 23477 14841 23489 14875
rect 23523 14872 23535 14875
rect 24305 14875 24363 14881
rect 24305 14872 24317 14875
rect 23523 14844 24317 14872
rect 23523 14841 23535 14844
rect 23477 14835 23535 14841
rect 24305 14841 24317 14844
rect 24351 14841 24363 14875
rect 24305 14835 24363 14841
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 5460 14776 8217 14804
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 11422 14804 11428 14816
rect 8720 14776 11428 14804
rect 8720 14764 8726 14776
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 14918 14764 14924 14816
rect 14976 14764 14982 14816
rect 18506 14764 18512 14816
rect 18564 14764 18570 14816
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14804 21695 14807
rect 22186 14804 22192 14816
rect 21683 14776 22192 14804
rect 21683 14773 21695 14776
rect 21637 14767 21695 14773
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 22833 14807 22891 14813
rect 22833 14804 22845 14807
rect 22612 14776 22845 14804
rect 22612 14764 22618 14776
rect 22833 14773 22845 14776
rect 22879 14773 22891 14807
rect 22833 14767 22891 14773
rect 24026 14764 24032 14816
rect 24084 14764 24090 14816
rect 24397 14807 24455 14813
rect 24397 14773 24409 14807
rect 24443 14804 24455 14807
rect 24443 14776 24900 14804
rect 24443 14773 24455 14776
rect 24397 14767 24455 14773
rect 1104 14714 24840 14736
rect 1104 14662 3917 14714
rect 3969 14662 3981 14714
rect 4033 14662 4045 14714
rect 4097 14662 4109 14714
rect 4161 14662 4173 14714
rect 4225 14662 9851 14714
rect 9903 14662 9915 14714
rect 9967 14662 9979 14714
rect 10031 14662 10043 14714
rect 10095 14662 10107 14714
rect 10159 14662 15785 14714
rect 15837 14662 15849 14714
rect 15901 14662 15913 14714
rect 15965 14662 15977 14714
rect 16029 14662 16041 14714
rect 16093 14662 21719 14714
rect 21771 14662 21783 14714
rect 21835 14662 21847 14714
rect 21899 14662 21911 14714
rect 21963 14662 21975 14714
rect 22027 14662 24840 14714
rect 1104 14640 24840 14662
rect 2866 14600 2872 14612
rect 2424 14572 2872 14600
rect 2424 14541 2452 14572
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 5074 14600 5080 14612
rect 4172 14572 5080 14600
rect 2409 14535 2467 14541
rect 2409 14501 2421 14535
rect 2455 14501 2467 14535
rect 2409 14495 2467 14501
rect 3510 14492 3516 14544
rect 3568 14532 3574 14544
rect 4065 14535 4123 14541
rect 4065 14532 4077 14535
rect 3568 14504 4077 14532
rect 3568 14492 3574 14504
rect 4065 14501 4077 14504
rect 4111 14501 4123 14535
rect 4065 14495 4123 14501
rect 2866 14473 2872 14476
rect 2823 14467 2872 14473
rect 2823 14433 2835 14467
rect 2869 14433 2872 14467
rect 2823 14427 2872 14433
rect 2866 14424 2872 14427
rect 2924 14464 2930 14476
rect 2924 14436 3924 14464
rect 2924 14424 2930 14436
rect 1302 14356 1308 14408
rect 1360 14396 1366 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1360 14368 1777 14396
rect 1360 14356 1366 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 1765 14359 1823 14365
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 2130 14396 2136 14408
rect 1995 14368 2136 14396
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 2130 14356 2136 14368
rect 2188 14356 2194 14408
rect 2682 14356 2688 14408
rect 2740 14356 2746 14408
rect 2958 14356 2964 14408
rect 3016 14356 3022 14408
rect 3896 14328 3924 14436
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4172 14396 4200 14572
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5902 14600 5908 14612
rect 5276 14572 5908 14600
rect 5276 14532 5304 14572
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 6564 14572 7512 14600
rect 6564 14544 6592 14572
rect 4448 14504 5304 14532
rect 4448 14476 4476 14504
rect 5350 14492 5356 14544
rect 5408 14532 5414 14544
rect 5537 14535 5595 14541
rect 5537 14532 5549 14535
rect 5408 14504 5549 14532
rect 5408 14492 5414 14504
rect 5537 14501 5549 14504
rect 5583 14501 5595 14535
rect 5537 14495 5595 14501
rect 6546 14492 6552 14544
rect 6604 14492 6610 14544
rect 6733 14535 6791 14541
rect 6733 14501 6745 14535
rect 6779 14532 6791 14535
rect 6822 14532 6828 14544
rect 6779 14504 6828 14532
rect 6779 14501 6791 14504
rect 6733 14495 6791 14501
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 7484 14532 7512 14572
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7616 14572 7849 14600
rect 7616 14560 7622 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 7837 14563 7895 14569
rect 10502 14560 10508 14612
rect 10560 14560 10566 14612
rect 12066 14560 12072 14612
rect 12124 14600 12130 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 12124 14572 12265 14600
rect 12124 14560 12130 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12253 14563 12311 14569
rect 12342 14560 12348 14612
rect 12400 14600 12406 14612
rect 12400 14572 13308 14600
rect 12400 14560 12406 14572
rect 10520 14532 10548 14560
rect 7484 14504 10548 14532
rect 4430 14424 4436 14476
rect 4488 14424 4494 14476
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 5442 14464 5448 14476
rect 4571 14436 5448 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 5442 14424 5448 14436
rect 5500 14424 5506 14476
rect 5902 14424 5908 14476
rect 5960 14473 5966 14476
rect 5960 14467 6009 14473
rect 5960 14433 5963 14467
rect 5997 14464 6009 14467
rect 5997 14436 6684 14464
rect 5997 14433 6009 14436
rect 5960 14427 6009 14433
rect 5960 14424 5966 14427
rect 4019 14368 4200 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4246 14356 4252 14408
rect 4304 14356 4310 14408
rect 4448 14328 4476 14424
rect 4614 14356 4620 14408
rect 4672 14356 4678 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 3436 14300 3832 14328
rect 3896 14300 4476 14328
rect 4632 14328 4660 14356
rect 4982 14328 4988 14340
rect 4632 14300 4988 14328
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 3436 14260 3464 14300
rect 2740 14232 3464 14260
rect 2740 14220 2746 14232
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 3804 14269 3832 14300
rect 4982 14288 4988 14300
rect 5040 14328 5046 14340
rect 5092 14328 5120 14359
rect 5810 14356 5816 14408
rect 5868 14356 5874 14408
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 5040 14300 5120 14328
rect 6656 14328 6684 14436
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8202 14464 8208 14476
rect 7616 14436 8208 14464
rect 7616 14424 7622 14436
rect 8202 14424 8208 14436
rect 8260 14424 8266 14476
rect 11238 14424 11244 14476
rect 11296 14424 11302 14476
rect 6730 14356 6736 14408
rect 6788 14396 6794 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6788 14368 6837 14396
rect 6788 14356 6794 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7006 14356 7012 14408
rect 7064 14396 7070 14408
rect 7099 14399 7157 14405
rect 7099 14396 7111 14399
rect 7064 14368 7111 14396
rect 7064 14356 7070 14368
rect 7099 14365 7111 14368
rect 7145 14365 7157 14399
rect 7099 14359 7157 14365
rect 7466 14356 7472 14408
rect 7524 14356 7530 14408
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 11514 14396 11520 14408
rect 10928 14368 11520 14396
rect 10928 14356 10934 14368
rect 11514 14356 11520 14368
rect 11572 14356 11578 14408
rect 12618 14356 12624 14408
rect 12676 14356 12682 14408
rect 12863 14399 12921 14405
rect 12863 14365 12875 14399
rect 12909 14365 12921 14399
rect 13280 14396 13308 14572
rect 14918 14560 14924 14612
rect 14976 14560 14982 14612
rect 16574 14600 16580 14612
rect 15028 14572 16580 14600
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13630 14532 13636 14544
rect 13412 14504 13636 14532
rect 13412 14492 13418 14504
rect 13630 14492 13636 14504
rect 13688 14492 13694 14544
rect 14734 14492 14740 14544
rect 14792 14492 14798 14544
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 14461 14467 14519 14473
rect 14461 14464 14473 14467
rect 13780 14436 14473 14464
rect 13780 14424 13786 14436
rect 14461 14433 14473 14436
rect 14507 14433 14519 14467
rect 14752 14464 14780 14492
rect 14936 14473 14964 14560
rect 14461 14427 14519 14433
rect 14568 14436 14780 14464
rect 14921 14467 14979 14473
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13280 14368 14289 14396
rect 12863 14359 12921 14365
rect 14277 14365 14289 14368
rect 14323 14396 14335 14399
rect 14568 14396 14596 14436
rect 14921 14433 14933 14467
rect 14967 14433 14979 14467
rect 15028 14464 15056 14572
rect 16574 14560 16580 14572
rect 16632 14600 16638 14612
rect 16942 14600 16948 14612
rect 16632 14572 16948 14600
rect 16632 14560 16638 14572
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 18506 14560 18512 14612
rect 18564 14560 18570 14612
rect 20254 14560 20260 14612
rect 20312 14560 20318 14612
rect 21545 14603 21603 14609
rect 21545 14569 21557 14603
rect 21591 14600 21603 14603
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21591 14572 21925 14600
rect 21591 14569 21603 14572
rect 21545 14563 21603 14569
rect 21913 14569 21925 14572
rect 21959 14569 21971 14603
rect 24872 14600 24900 14776
rect 25498 14696 25504 14748
rect 25556 14696 25562 14748
rect 21913 14563 21971 14569
rect 23492 14572 24900 14600
rect 18141 14535 18199 14541
rect 16684 14504 16970 14532
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 15028 14436 15209 14464
rect 14921 14427 14979 14433
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15335 14467 15393 14473
rect 15335 14433 15347 14467
rect 15381 14464 15393 14467
rect 16114 14464 16120 14476
rect 15381 14436 16120 14464
rect 15381 14433 15393 14436
rect 15335 14427 15393 14433
rect 16114 14424 16120 14436
rect 16172 14464 16178 14476
rect 16684 14464 16712 14504
rect 16172 14436 16712 14464
rect 16172 14424 16178 14436
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 16942 14464 16970 14504
rect 18141 14501 18153 14535
rect 18187 14501 18199 14535
rect 18141 14495 18199 14501
rect 17218 14464 17224 14476
rect 17276 14473 17282 14476
rect 17276 14467 17304 14473
rect 16942 14436 17224 14464
rect 17218 14424 17224 14436
rect 17292 14433 17304 14467
rect 17276 14427 17304 14433
rect 17276 14424 17282 14427
rect 17770 14424 17776 14476
rect 17828 14464 17834 14476
rect 18049 14467 18107 14473
rect 18049 14464 18061 14467
rect 17828 14436 18061 14464
rect 17828 14424 17834 14436
rect 18049 14433 18061 14436
rect 18095 14433 18107 14467
rect 18156 14464 18184 14495
rect 18156 14436 18460 14464
rect 18049 14427 18107 14433
rect 14323 14368 14596 14396
rect 14323 14365 14335 14368
rect 14277 14359 14335 14365
rect 7484 14328 7512 14356
rect 11882 14328 11888 14340
rect 6656 14300 7512 14328
rect 8404 14300 11888 14328
rect 5040 14288 5046 14300
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 4338 14220 4344 14272
rect 4396 14260 4402 14272
rect 8404 14260 8432 14300
rect 11882 14288 11888 14300
rect 11940 14288 11946 14340
rect 12878 14328 12906 14359
rect 15470 14356 15476 14408
rect 15528 14356 15534 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14396 16267 14399
rect 16298 14396 16304 14408
rect 16255 14368 16304 14396
rect 16255 14365 16267 14368
rect 16209 14359 16267 14365
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16390 14356 16396 14408
rect 16448 14356 16454 14408
rect 17126 14356 17132 14408
rect 17184 14356 17190 14408
rect 17402 14356 17408 14408
rect 17460 14356 17466 14408
rect 18432 14405 18460 14436
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18524 14396 18552 14560
rect 18877 14399 18935 14405
rect 18877 14396 18889 14399
rect 18524 14368 18889 14396
rect 18417 14359 18475 14365
rect 18877 14365 18889 14368
rect 18923 14365 18935 14399
rect 20272 14396 20300 14560
rect 22462 14532 22468 14544
rect 21836 14504 22468 14532
rect 21836 14405 21864 14504
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 22557 14467 22615 14473
rect 22557 14464 22569 14467
rect 22143 14436 22569 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 22557 14433 22569 14436
rect 22603 14433 22615 14467
rect 22557 14427 22615 14433
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20272 14368 21097 14396
rect 18877 14359 18935 14365
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 12360 14300 12906 14328
rect 4396 14232 8432 14260
rect 4396 14220 4402 14232
rect 12066 14220 12072 14272
rect 12124 14260 12130 14272
rect 12360 14260 12388 14300
rect 16114 14288 16120 14340
rect 16172 14288 16178 14340
rect 12124 14232 12388 14260
rect 12124 14220 12130 14232
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13228 14232 13645 14260
rect 13228 14220 13234 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 17310 14220 17316 14272
rect 17368 14260 17374 14272
rect 17862 14260 17868 14272
rect 17368 14232 17868 14260
rect 17368 14220 17374 14232
rect 17862 14220 17868 14232
rect 17920 14260 17926 14272
rect 18340 14260 18368 14359
rect 21468 14328 21496 14359
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 22373 14399 22431 14405
rect 22373 14396 22385 14399
rect 22244 14368 22385 14396
rect 22244 14356 22250 14368
rect 22373 14365 22385 14368
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 23385 14399 23443 14405
rect 23385 14365 23397 14399
rect 23431 14396 23443 14399
rect 23492 14396 23520 14572
rect 23569 14535 23627 14541
rect 23569 14501 23581 14535
rect 23615 14532 23627 14535
rect 25130 14532 25136 14544
rect 23615 14504 25136 14532
rect 23615 14501 23627 14504
rect 23569 14495 23627 14501
rect 25130 14492 25136 14504
rect 25188 14492 25194 14544
rect 23750 14424 23756 14476
rect 23808 14424 23814 14476
rect 24121 14467 24179 14473
rect 24121 14433 24133 14467
rect 24167 14464 24179 14467
rect 25516 14464 25544 14696
rect 24167 14436 25544 14464
rect 24167 14433 24179 14436
rect 24121 14427 24179 14433
rect 23431 14368 23520 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 22664 14328 22692 14359
rect 23308 14328 23336 14359
rect 23768 14328 23796 14424
rect 23845 14399 23903 14405
rect 23845 14365 23857 14399
rect 23891 14396 23903 14399
rect 23891 14368 24164 14396
rect 23891 14365 23903 14368
rect 23845 14359 23903 14365
rect 24136 14340 24164 14368
rect 20916 14300 21496 14328
rect 22204 14300 22692 14328
rect 22756 14300 23244 14328
rect 23308 14300 23796 14328
rect 17920 14232 18368 14260
rect 17920 14220 17926 14232
rect 18506 14220 18512 14272
rect 18564 14220 18570 14272
rect 18693 14263 18751 14269
rect 18693 14229 18705 14263
rect 18739 14260 18751 14263
rect 19150 14260 19156 14272
rect 18739 14232 19156 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 20916 14269 20944 14300
rect 20901 14263 20959 14269
rect 20901 14229 20913 14263
rect 20947 14229 20959 14263
rect 20901 14223 20959 14229
rect 21634 14220 21640 14272
rect 21692 14260 21698 14272
rect 22204 14269 22232 14300
rect 22756 14272 22784 14300
rect 22097 14263 22155 14269
rect 22097 14260 22109 14263
rect 21692 14232 22109 14260
rect 21692 14220 21698 14232
rect 22097 14229 22109 14232
rect 22143 14229 22155 14263
rect 22097 14223 22155 14229
rect 22189 14263 22247 14269
rect 22189 14229 22201 14263
rect 22235 14229 22247 14263
rect 22189 14223 22247 14229
rect 22738 14220 22744 14272
rect 22796 14220 22802 14272
rect 23106 14220 23112 14272
rect 23164 14220 23170 14272
rect 23216 14260 23244 14300
rect 24118 14288 24124 14340
rect 24176 14288 24182 14340
rect 24210 14260 24216 14272
rect 23216 14232 24216 14260
rect 24210 14220 24216 14232
rect 24268 14220 24274 14272
rect 1104 14170 25000 14192
rect 1104 14118 6884 14170
rect 6936 14118 6948 14170
rect 7000 14118 7012 14170
rect 7064 14118 7076 14170
rect 7128 14118 7140 14170
rect 7192 14118 12818 14170
rect 12870 14118 12882 14170
rect 12934 14118 12946 14170
rect 12998 14118 13010 14170
rect 13062 14118 13074 14170
rect 13126 14118 18752 14170
rect 18804 14118 18816 14170
rect 18868 14118 18880 14170
rect 18932 14118 18944 14170
rect 18996 14118 19008 14170
rect 19060 14118 24686 14170
rect 24738 14118 24750 14170
rect 24802 14118 24814 14170
rect 24866 14118 24878 14170
rect 24930 14118 24942 14170
rect 24994 14118 25000 14170
rect 1104 14096 25000 14118
rect 1394 14016 1400 14068
rect 1452 14056 1458 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 1452 14028 1593 14056
rect 1452 14016 1458 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 1581 14019 1639 14025
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3237 14059 3295 14065
rect 3237 14056 3249 14059
rect 3016 14028 3249 14056
rect 3016 14016 3022 14028
rect 3237 14025 3249 14028
rect 3283 14025 3295 14059
rect 3237 14019 3295 14025
rect 5905 14059 5963 14065
rect 5905 14025 5917 14059
rect 5951 14056 5963 14059
rect 6086 14056 6092 14068
rect 5951 14028 6092 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 12158 14056 12164 14068
rect 6420 14028 12164 14056
rect 6420 14016 6426 14028
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 12618 14016 12624 14068
rect 12676 14056 12682 14068
rect 12802 14056 12808 14068
rect 12676 14028 12808 14056
rect 12676 14016 12682 14028
rect 12802 14016 12808 14028
rect 12860 14056 12866 14068
rect 13906 14056 13912 14068
rect 12860 14028 13912 14056
rect 12860 14016 12866 14028
rect 13906 14016 13912 14028
rect 13964 14056 13970 14068
rect 13964 14028 14136 14056
rect 13964 14016 13970 14028
rect 1489 13991 1547 13997
rect 1489 13957 1501 13991
rect 1535 13988 1547 13991
rect 6546 13988 6552 14000
rect 1535 13960 6552 13988
rect 1535 13957 1547 13960
rect 1489 13951 1547 13957
rect 6546 13948 6552 13960
rect 6604 13948 6610 14000
rect 7466 13948 7472 14000
rect 7524 13988 7530 14000
rect 11698 13988 11704 14000
rect 7524 13960 11704 13988
rect 7524 13948 7530 13960
rect 11698 13948 11704 13960
rect 11756 13948 11762 14000
rect 14108 13988 14136 14028
rect 14274 14016 14280 14068
rect 14332 14016 14338 14068
rect 15286 14016 15292 14068
rect 15344 14016 15350 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15528 14028 15669 14056
rect 15528 14016 15534 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 16816 14028 17356 14056
rect 16816 14016 16822 14028
rect 14108 13960 14688 13988
rect 1946 13880 1952 13932
rect 2004 13920 2010 13932
rect 2133 13923 2191 13929
rect 2133 13920 2145 13923
rect 2004 13892 2145 13920
rect 2004 13880 2010 13892
rect 2133 13889 2145 13892
rect 2179 13889 2191 13923
rect 2133 13883 2191 13889
rect 2406 13880 2412 13932
rect 2464 13920 2470 13932
rect 2499 13923 2557 13929
rect 2499 13920 2511 13923
rect 2464 13892 2511 13920
rect 2464 13880 2470 13892
rect 2499 13889 2511 13892
rect 2545 13889 2557 13923
rect 2499 13883 2557 13889
rect 3694 13880 3700 13932
rect 3752 13880 3758 13932
rect 4338 13880 4344 13932
rect 4396 13880 4402 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5167 13923 5225 13929
rect 5167 13920 5179 13923
rect 5132 13892 5179 13920
rect 5132 13880 5138 13892
rect 5167 13889 5179 13892
rect 5213 13920 5225 13923
rect 5258 13920 5264 13932
rect 5213 13892 5264 13920
rect 5213 13889 5225 13892
rect 5167 13883 5225 13889
rect 5258 13880 5264 13892
rect 5316 13880 5322 13932
rect 6730 13880 6736 13932
rect 6788 13920 6794 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6788 13892 6837 13920
rect 6788 13880 6794 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 7099 13923 7157 13929
rect 7099 13889 7111 13923
rect 7145 13920 7157 13923
rect 8110 13920 8116 13932
rect 7145 13892 8116 13920
rect 7145 13889 7157 13892
rect 7099 13883 7157 13889
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13821 2283 13855
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 2225 13815 2283 13821
rect 2884 13824 4905 13852
rect 2240 13784 2268 13815
rect 2240 13756 2360 13784
rect 2332 13728 2360 13756
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2884 13716 2912 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 4157 13787 4215 13793
rect 4157 13784 4169 13787
rect 3016 13756 4169 13784
rect 3016 13744 3022 13756
rect 4157 13753 4169 13756
rect 4203 13753 4215 13787
rect 4157 13747 4215 13753
rect 2372 13688 2912 13716
rect 2372 13676 2378 13688
rect 3786 13676 3792 13728
rect 3844 13676 3850 13728
rect 6840 13716 6868 13883
rect 8110 13880 8116 13892
rect 8168 13880 8174 13932
rect 8479 13923 8537 13929
rect 8479 13889 8491 13923
rect 8525 13920 8537 13923
rect 8846 13920 8852 13932
rect 8525 13892 8852 13920
rect 8525 13889 8537 13892
rect 8479 13883 8537 13889
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 9858 13929 9864 13932
rect 9827 13923 9864 13929
rect 9827 13889 9839 13923
rect 9827 13883 9864 13889
rect 9858 13880 9864 13883
rect 9916 13880 9922 13932
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 12483 13892 12848 13920
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7484 13824 8217 13852
rect 7484 13716 7512 13824
rect 8205 13821 8217 13824
rect 8251 13821 8263 13855
rect 9306 13852 9312 13864
rect 8205 13815 8263 13821
rect 8864 13824 9312 13852
rect 6840 13688 7512 13716
rect 7834 13676 7840 13728
rect 7892 13676 7898 13728
rect 8220 13716 8248 13815
rect 8864 13716 8892 13824
rect 9306 13812 9312 13824
rect 9364 13852 9370 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9364 13824 9597 13852
rect 9364 13812 9370 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 12618 13812 12624 13864
rect 12676 13812 12682 13864
rect 12820 13852 12848 13892
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 13495 13923 13553 13929
rect 13495 13889 13507 13923
rect 13541 13920 13553 13923
rect 13541 13898 13584 13920
rect 13541 13889 13544 13898
rect 13495 13883 13544 13889
rect 13081 13855 13139 13861
rect 12820 13824 13032 13852
rect 8938 13744 8944 13796
rect 8996 13784 9002 13796
rect 8996 13756 9674 13784
rect 8996 13744 9002 13756
rect 8220 13688 8892 13716
rect 9214 13676 9220 13728
rect 9272 13676 9278 13728
rect 9646 13716 9674 13756
rect 10410 13716 10416 13728
rect 9646 13688 10416 13716
rect 10410 13676 10416 13688
rect 10468 13676 10474 13728
rect 10502 13676 10508 13728
rect 10560 13716 10566 13728
rect 10597 13719 10655 13725
rect 10597 13716 10609 13719
rect 10560 13688 10609 13716
rect 10560 13676 10566 13688
rect 10597 13685 10609 13688
rect 10643 13685 10655 13719
rect 13004 13716 13032 13824
rect 13081 13821 13093 13855
rect 13127 13852 13139 13855
rect 13170 13852 13176 13864
rect 13127 13824 13176 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13538 13846 13544 13883
rect 13596 13846 13602 13898
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 14550 13852 14556 13864
rect 14016 13824 14556 13852
rect 14016 13716 14044 13824
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 14660 13861 14688 13960
rect 14903 13953 14961 13959
rect 14903 13919 14915 13953
rect 14949 13950 14961 13953
rect 14949 13932 14964 13950
rect 15194 13948 15200 14000
rect 15252 13948 15258 14000
rect 15304 13988 15332 14016
rect 17328 13988 17356 14028
rect 17402 14016 17408 14068
rect 17460 14056 17466 14068
rect 17681 14059 17739 14065
rect 17681 14056 17693 14059
rect 17460 14028 17693 14056
rect 17460 14016 17466 14028
rect 17681 14025 17693 14028
rect 17727 14025 17739 14059
rect 17681 14019 17739 14025
rect 17770 14016 17776 14068
rect 17828 14056 17834 14068
rect 20806 14056 20812 14068
rect 17828 14028 20812 14056
rect 17828 14016 17834 14028
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 22278 14016 22284 14068
rect 22336 14056 22342 14068
rect 23014 14056 23020 14068
rect 22336 14028 23020 14056
rect 22336 14016 22342 14028
rect 23014 14016 23020 14028
rect 23072 14016 23078 14068
rect 23106 14016 23112 14068
rect 23164 14016 23170 14068
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14025 23259 14059
rect 23201 14019 23259 14025
rect 18138 13988 18144 14000
rect 15304 13960 16954 13988
rect 17328 13960 18144 13988
rect 16926 13959 16954 13960
rect 16926 13953 16985 13959
rect 14903 13913 14924 13919
rect 14918 13880 14924 13913
rect 14976 13880 14982 13932
rect 15212 13920 15240 13948
rect 16114 13920 16120 13932
rect 15212 13892 16120 13920
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16482 13880 16488 13932
rect 16540 13920 16546 13932
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16540 13892 16681 13920
rect 16540 13880 16546 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16926 13922 16939 13953
rect 16927 13919 16939 13922
rect 16973 13920 16985 13953
rect 18138 13948 18144 13960
rect 18196 13988 18202 14000
rect 18196 13960 18334 13988
rect 18196 13948 18202 13960
rect 17402 13920 17408 13932
rect 16973 13919 17408 13920
rect 16927 13913 17408 13919
rect 16942 13892 17408 13913
rect 16669 13883 16727 13889
rect 14645 13855 14703 13861
rect 14645 13821 14657 13855
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14660 13784 14688 13815
rect 14568 13756 14688 13784
rect 14568 13728 14596 13756
rect 13004 13688 14044 13716
rect 10597 13679 10655 13685
rect 14550 13676 14556 13728
rect 14608 13676 14614 13728
rect 16684 13716 16712 13883
rect 17402 13880 17408 13892
rect 17460 13880 17466 13932
rect 18306 13929 18334 13960
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 19208 13960 19656 13988
rect 19208 13948 19214 13960
rect 19628 13929 19656 13960
rect 22830 13948 22836 14000
rect 22888 13948 22894 14000
rect 23124 13988 23152 14016
rect 22940 13960 23152 13988
rect 23216 13988 23244 14019
rect 23845 13991 23903 13997
rect 23845 13988 23857 13991
rect 23216 13960 23857 13988
rect 18291 13923 18349 13929
rect 18291 13889 18303 13923
rect 18337 13889 18349 13923
rect 19429 13923 19487 13929
rect 19429 13920 19441 13923
rect 18291 13883 18349 13889
rect 18892 13892 19441 13920
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 18012 13824 18061 13852
rect 18012 13812 18018 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18892 13796 18920 13892
rect 19429 13889 19441 13892
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 22462 13920 22468 13932
rect 20956 13892 22468 13920
rect 20956 13880 20962 13892
rect 22462 13880 22468 13892
rect 22520 13880 22526 13932
rect 22738 13880 22744 13932
rect 22796 13880 22802 13932
rect 22940 13929 22968 13960
rect 23845 13957 23857 13960
rect 23891 13957 23903 13991
rect 23845 13951 23903 13957
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13889 23075 13923
rect 23017 13883 23075 13889
rect 19150 13812 19156 13864
rect 19208 13852 19214 13864
rect 19521 13855 19579 13861
rect 19521 13852 19533 13855
rect 19208 13824 19533 13852
rect 19208 13812 19214 13824
rect 19521 13821 19533 13824
rect 19567 13821 19579 13855
rect 23032 13852 23060 13883
rect 23106 13880 23112 13932
rect 23164 13920 23170 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 23164 13892 23213 13920
rect 23164 13880 23170 13892
rect 23201 13889 23213 13892
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23290 13880 23296 13932
rect 23348 13920 23354 13932
rect 23477 13923 23535 13929
rect 23477 13920 23489 13923
rect 23348 13892 23489 13920
rect 23348 13880 23354 13892
rect 23477 13889 23489 13892
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 24121 13923 24179 13929
rect 24121 13889 24133 13923
rect 24167 13889 24179 13923
rect 24121 13883 24179 13889
rect 23382 13852 23388 13864
rect 23032 13824 23388 13852
rect 19521 13815 19579 13821
rect 23382 13812 23388 13824
rect 23440 13812 23446 13864
rect 18874 13744 18880 13796
rect 18932 13784 18938 13796
rect 19061 13787 19119 13793
rect 19061 13784 19073 13787
rect 18932 13756 19073 13784
rect 18932 13744 18938 13756
rect 19061 13753 19073 13756
rect 19107 13753 19119 13787
rect 19061 13747 19119 13753
rect 20438 13744 20444 13796
rect 20496 13784 20502 13796
rect 20496 13756 21404 13784
rect 20496 13744 20502 13756
rect 21266 13716 21272 13728
rect 16684 13688 21272 13716
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 21376 13716 21404 13756
rect 23474 13744 23480 13796
rect 23532 13744 23538 13796
rect 24136 13716 24164 13883
rect 21376 13688 24164 13716
rect 24394 13676 24400 13728
rect 24452 13676 24458 13728
rect 1104 13626 24840 13648
rect 1104 13574 3917 13626
rect 3969 13574 3981 13626
rect 4033 13574 4045 13626
rect 4097 13574 4109 13626
rect 4161 13574 4173 13626
rect 4225 13574 9851 13626
rect 9903 13574 9915 13626
rect 9967 13574 9979 13626
rect 10031 13574 10043 13626
rect 10095 13574 10107 13626
rect 10159 13574 15785 13626
rect 15837 13574 15849 13626
rect 15901 13574 15913 13626
rect 15965 13574 15977 13626
rect 16029 13574 16041 13626
rect 16093 13574 21719 13626
rect 21771 13574 21783 13626
rect 21835 13574 21847 13626
rect 21899 13574 21911 13626
rect 21963 13574 21975 13626
rect 22027 13574 24840 13626
rect 1104 13552 24840 13574
rect 1210 13472 1216 13524
rect 1268 13512 1274 13524
rect 2317 13515 2375 13521
rect 2317 13512 2329 13515
rect 1268 13484 2329 13512
rect 1268 13472 1274 13484
rect 2317 13481 2329 13484
rect 2363 13481 2375 13515
rect 2317 13475 2375 13481
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2832 13484 2881 13512
rect 2832 13472 2838 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 9122 13512 9128 13524
rect 2869 13475 2927 13481
rect 8220 13484 9128 13512
rect 8220 13456 8248 13484
rect 9122 13472 9128 13484
rect 9180 13512 9186 13524
rect 9180 13484 9674 13512
rect 9180 13472 9186 13484
rect 1670 13404 1676 13456
rect 1728 13404 1734 13456
rect 8202 13404 8208 13456
rect 8260 13404 8266 13456
rect 8386 13404 8392 13456
rect 8444 13444 8450 13456
rect 9309 13447 9367 13453
rect 9309 13444 9321 13447
rect 8444 13416 9321 13444
rect 8444 13404 8450 13416
rect 9309 13413 9321 13416
rect 9355 13413 9367 13447
rect 9309 13407 9367 13413
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 3234 13376 3240 13388
rect 2096 13348 3240 13376
rect 2096 13336 2102 13348
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 3344 13348 3556 13376
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13308 1547 13311
rect 3344 13308 3372 13348
rect 3528 13320 3556 13348
rect 3786 13336 3792 13388
rect 3844 13336 3850 13388
rect 7282 13336 7288 13388
rect 7340 13376 7346 13388
rect 8938 13376 8944 13388
rect 7340 13348 8944 13376
rect 7340 13336 7346 13348
rect 8938 13336 8944 13348
rect 8996 13336 9002 13388
rect 9646 13376 9674 13484
rect 10410 13472 10416 13524
rect 10468 13472 10474 13524
rect 10778 13512 10784 13524
rect 10520 13484 10784 13512
rect 9953 13379 10011 13385
rect 9953 13376 9965 13379
rect 9646 13348 9965 13376
rect 9953 13345 9965 13348
rect 9999 13376 10011 13379
rect 10134 13376 10140 13388
rect 9999 13348 10140 13376
rect 9999 13345 10011 13348
rect 9953 13339 10011 13345
rect 10134 13336 10140 13348
rect 10192 13336 10198 13388
rect 10428 13385 10456 13472
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13345 10471 13379
rect 10520 13376 10548 13484
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11422 13472 11428 13524
rect 11480 13512 11486 13524
rect 12710 13512 12716 13524
rect 11480 13484 12716 13512
rect 11480 13472 11486 13484
rect 12710 13472 12716 13484
rect 12768 13512 12774 13524
rect 12768 13484 13584 13512
rect 12768 13472 12774 13484
rect 10827 13379 10885 13385
rect 10520 13348 10732 13376
rect 10413 13339 10471 13345
rect 9493 13327 9551 13333
rect 9493 13320 9505 13327
rect 9539 13320 9551 13327
rect 1535 13280 3372 13308
rect 3421 13311 3479 13317
rect 1535 13277 1547 13280
rect 1489 13271 1547 13277
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 290 13200 296 13252
rect 348 13240 354 13252
rect 842 13240 848 13252
rect 348 13212 848 13240
rect 348 13200 354 13212
rect 842 13200 848 13212
rect 900 13200 906 13252
rect 1578 13200 1584 13252
rect 1636 13240 1642 13252
rect 2225 13243 2283 13249
rect 2225 13240 2237 13243
rect 1636 13212 2237 13240
rect 1636 13200 1642 13212
rect 2225 13209 2237 13212
rect 2271 13209 2283 13243
rect 2225 13203 2283 13209
rect 2774 13200 2780 13252
rect 2832 13200 2838 13252
rect 3436 13240 3464 13271
rect 3510 13268 3516 13320
rect 3568 13268 3574 13320
rect 4062 13317 4068 13320
rect 4047 13311 4068 13317
rect 4047 13277 4059 13311
rect 4047 13271 4068 13277
rect 4062 13268 4068 13271
rect 4120 13268 4126 13320
rect 4430 13268 4436 13320
rect 4488 13308 4494 13320
rect 5442 13308 5448 13320
rect 4488 13280 5448 13308
rect 4488 13268 4494 13280
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8076 13280 9444 13308
rect 8076 13268 8082 13280
rect 9416 13240 9444 13280
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 10704 13317 10732 13348
rect 10827 13345 10839 13379
rect 10873 13376 10885 13379
rect 10873 13348 11560 13376
rect 10873 13345 10885 13348
rect 10827 13339 10885 13345
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 9784 13240 9812 13271
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 9950 13240 9956 13252
rect 3436 13212 9352 13240
rect 9416 13212 9956 13240
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13172 3295 13175
rect 3786 13172 3792 13184
rect 3283 13144 3792 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 4430 13132 4436 13184
rect 4488 13172 4494 13184
rect 4801 13175 4859 13181
rect 4801 13172 4813 13175
rect 4488 13144 4813 13172
rect 4488 13132 4494 13144
rect 4801 13141 4813 13144
rect 4847 13141 4859 13175
rect 4801 13135 4859 13141
rect 5258 13132 5264 13184
rect 5316 13172 5322 13184
rect 8386 13172 8392 13184
rect 5316 13144 8392 13172
rect 5316 13132 5322 13144
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9324 13172 9352 13212
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 11532 13240 11560 13348
rect 12158 13336 12164 13388
rect 12216 13376 12222 13388
rect 12342 13376 12348 13388
rect 12216 13348 12348 13376
rect 12216 13336 12222 13348
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 13556 13376 13584 13484
rect 13630 13472 13636 13524
rect 13688 13472 13694 13524
rect 16485 13515 16543 13521
rect 15488 13484 16160 13512
rect 15488 13385 15516 13484
rect 15473 13379 15531 13385
rect 13556 13348 14136 13376
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 11664 13280 12633 13308
rect 11664 13268 11670 13280
rect 12621 13277 12633 13280
rect 12667 13308 12679 13311
rect 12802 13308 12808 13320
rect 12667 13280 12808 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 12895 13311 12953 13317
rect 12895 13277 12907 13311
rect 12941 13308 12953 13311
rect 13814 13308 13820 13320
rect 12941 13280 13820 13308
rect 12941 13277 12953 13280
rect 12895 13271 12953 13277
rect 13648 13252 13676 13280
rect 13814 13268 13820 13280
rect 13872 13268 13878 13320
rect 14108 13308 14136 13348
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 16132 13376 16160 13484
rect 16485 13481 16497 13515
rect 16531 13512 16543 13515
rect 16850 13512 16856 13524
rect 16531 13484 16856 13512
rect 16531 13481 16543 13484
rect 16485 13475 16543 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 18506 13472 18512 13524
rect 18564 13512 18570 13524
rect 18601 13515 18659 13521
rect 18601 13512 18613 13515
rect 18564 13484 18613 13512
rect 18564 13472 18570 13484
rect 18601 13481 18613 13484
rect 18647 13481 18659 13515
rect 18601 13475 18659 13481
rect 18693 13515 18751 13521
rect 18693 13481 18705 13515
rect 18739 13512 18751 13515
rect 20438 13512 20444 13524
rect 18739 13484 20444 13512
rect 18739 13481 18751 13484
rect 18693 13475 18751 13481
rect 20438 13472 20444 13484
rect 20496 13472 20502 13524
rect 22649 13515 22707 13521
rect 22649 13481 22661 13515
rect 22695 13512 22707 13515
rect 23198 13512 23204 13524
rect 22695 13484 23204 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 16942 13404 16948 13456
rect 17000 13444 17006 13456
rect 19518 13444 19524 13456
rect 17000 13416 19524 13444
rect 17000 13404 17006 13416
rect 19518 13404 19524 13416
rect 19576 13404 19582 13456
rect 19720 13416 20668 13444
rect 16482 13376 16488 13388
rect 16132 13348 16488 13376
rect 15473 13339 15531 13345
rect 16482 13336 16488 13348
rect 16540 13336 16546 13388
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13376 18843 13379
rect 18966 13376 18972 13388
rect 18831 13348 18972 13376
rect 18831 13345 18843 13348
rect 18785 13339 18843 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 15194 13308 15200 13320
rect 14108 13280 15200 13308
rect 15194 13268 15200 13280
rect 15252 13308 15258 13320
rect 15715 13311 15773 13317
rect 15715 13308 15727 13311
rect 15252 13280 15727 13308
rect 15252 13268 15258 13280
rect 15715 13277 15727 13280
rect 15761 13308 15773 13311
rect 17770 13308 17776 13320
rect 15761 13280 17776 13308
rect 15761 13277 15773 13280
rect 15715 13271 15773 13277
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 18874 13308 18880 13320
rect 18555 13280 18880 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 18874 13268 18880 13280
rect 18932 13268 18938 13320
rect 19720 13317 19748 13416
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 19904 13348 20453 13376
rect 19904 13317 19932 13348
rect 20441 13345 20453 13348
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19260 13280 19717 13308
rect 13538 13240 13544 13252
rect 11532 13212 13544 13240
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 13630 13200 13636 13252
rect 13688 13200 13694 13252
rect 19260 13184 19288 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 20346 13268 20352 13320
rect 20404 13268 20410 13320
rect 20640 13317 20668 13416
rect 22278 13404 22284 13456
rect 22336 13404 22342 13456
rect 22833 13379 22891 13385
rect 22833 13376 22845 13379
rect 21192 13348 22845 13376
rect 21192 13320 21220 13348
rect 22833 13345 22845 13348
rect 22879 13345 22891 13379
rect 22833 13339 22891 13345
rect 20625 13311 20683 13317
rect 20625 13277 20637 13311
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 20806 13268 20812 13320
rect 20864 13268 20870 13320
rect 21174 13268 21180 13320
rect 21232 13268 21238 13320
rect 22465 13311 22523 13317
rect 22465 13277 22477 13311
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 22581 13313 22639 13319
rect 22581 13279 22593 13313
rect 22627 13310 22639 13313
rect 22627 13308 22784 13310
rect 23474 13308 23480 13320
rect 22627 13282 23480 13308
rect 22627 13279 22639 13282
rect 22756 13280 23480 13282
rect 22581 13273 22639 13279
rect 20162 13200 20168 13252
rect 20220 13200 20226 13252
rect 20257 13243 20315 13249
rect 20257 13209 20269 13243
rect 20303 13240 20315 13243
rect 20717 13243 20775 13249
rect 20717 13240 20729 13243
rect 20303 13212 20729 13240
rect 20303 13209 20315 13212
rect 20257 13203 20315 13209
rect 20717 13209 20729 13212
rect 20763 13209 20775 13243
rect 22480 13240 22508 13271
rect 23474 13268 23480 13280
rect 23532 13268 23538 13320
rect 23100 13243 23158 13249
rect 22480 13212 22600 13240
rect 20717 13203 20775 13209
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 9324 13144 11621 13172
rect 11609 13141 11621 13144
rect 11655 13141 11667 13175
rect 11609 13135 11667 13141
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 21450 13172 21456 13184
rect 19392 13144 21456 13172
rect 19392 13132 19398 13144
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 22572 13172 22600 13212
rect 23100 13209 23112 13243
rect 23146 13240 23158 13243
rect 23198 13240 23204 13252
rect 23146 13212 23204 13240
rect 23146 13209 23158 13212
rect 23100 13203 23158 13209
rect 23198 13200 23204 13212
rect 23256 13200 23262 13252
rect 24213 13175 24271 13181
rect 24213 13172 24225 13175
rect 22572 13144 24225 13172
rect 24213 13141 24225 13144
rect 24259 13141 24271 13175
rect 24213 13135 24271 13141
rect 1104 13082 25000 13104
rect 1104 13030 6884 13082
rect 6936 13030 6948 13082
rect 7000 13030 7012 13082
rect 7064 13030 7076 13082
rect 7128 13030 7140 13082
rect 7192 13030 12818 13082
rect 12870 13030 12882 13082
rect 12934 13030 12946 13082
rect 12998 13030 13010 13082
rect 13062 13030 13074 13082
rect 13126 13030 18752 13082
rect 18804 13030 18816 13082
rect 18868 13030 18880 13082
rect 18932 13030 18944 13082
rect 18996 13030 19008 13082
rect 19060 13030 24686 13082
rect 24738 13030 24750 13082
rect 24802 13030 24814 13082
rect 24866 13030 24878 13082
rect 24930 13030 24942 13082
rect 24994 13030 25000 13082
rect 1104 13008 25000 13030
rect 1504 12940 3004 12968
rect 1504 12909 1532 12940
rect 2976 12912 3004 12940
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 4338 12968 4344 12980
rect 3844 12940 4344 12968
rect 3844 12928 3850 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 5810 12968 5816 12980
rect 5592 12940 5816 12968
rect 5592 12928 5598 12940
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6822 12968 6828 12980
rect 6052 12940 6828 12968
rect 6052 12928 6058 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 7926 12968 7932 12980
rect 7248 12940 7932 12968
rect 7248 12928 7254 12940
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9490 12928 9496 12980
rect 9548 12968 9554 12980
rect 9861 12971 9919 12977
rect 9861 12968 9873 12971
rect 9548 12940 9873 12968
rect 9548 12928 9554 12940
rect 9861 12937 9873 12940
rect 9907 12937 9919 12971
rect 9861 12931 9919 12937
rect 9950 12928 9956 12980
rect 10008 12928 10014 12980
rect 10226 12928 10232 12980
rect 10284 12968 10290 12980
rect 10870 12968 10876 12980
rect 10284 12940 10876 12968
rect 10284 12928 10290 12940
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 11020 12940 11069 12968
rect 11020 12928 11026 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 20162 12968 20168 12980
rect 11057 12931 11115 12937
rect 11164 12940 20168 12968
rect 1489 12903 1547 12909
rect 1489 12869 1501 12903
rect 1535 12869 1547 12903
rect 1489 12863 1547 12869
rect 1854 12860 1860 12912
rect 1912 12860 1918 12912
rect 2406 12900 2412 12912
rect 2332 12872 2412 12900
rect 2332 12841 2360 12872
rect 2406 12860 2412 12872
rect 2464 12860 2470 12912
rect 2958 12860 2964 12912
rect 3016 12860 3022 12912
rect 3878 12900 3884 12912
rect 3160 12872 3884 12900
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12801 2375 12835
rect 2317 12795 2375 12801
rect 2591 12835 2649 12841
rect 2591 12801 2603 12835
rect 2637 12832 2649 12835
rect 3160 12832 3188 12872
rect 3878 12860 3884 12872
rect 3936 12860 3942 12912
rect 7208 12900 7236 12928
rect 6196 12872 7236 12900
rect 9968 12900 9996 12928
rect 11164 12900 11192 12940
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 20864 12940 21373 12968
rect 20864 12928 20870 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 21361 12931 21419 12937
rect 22186 12928 22192 12980
rect 22244 12928 22250 12980
rect 22646 12928 22652 12980
rect 22704 12928 22710 12980
rect 23382 12928 23388 12980
rect 23440 12928 23446 12980
rect 9968 12872 11192 12900
rect 2637 12804 3188 12832
rect 2637 12801 2649 12804
rect 2591 12795 2649 12801
rect 2222 12656 2228 12708
rect 2280 12696 2286 12708
rect 2332 12696 2360 12795
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 3292 12804 3709 12832
rect 3292 12792 3298 12804
rect 3697 12801 3709 12804
rect 3743 12832 3755 12835
rect 3743 12804 4108 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4080 12776 4108 12804
rect 4706 12792 4712 12844
rect 4764 12841 4770 12844
rect 4764 12835 4792 12841
rect 4780 12801 4792 12835
rect 4764 12795 4792 12801
rect 4764 12792 4770 12795
rect 4890 12792 4896 12844
rect 4948 12792 4954 12844
rect 3050 12724 3056 12776
rect 3108 12764 3114 12776
rect 3326 12764 3332 12776
rect 3108 12736 3332 12764
rect 3108 12724 3114 12736
rect 3326 12724 3332 12736
rect 3384 12764 3390 12776
rect 3881 12767 3939 12773
rect 3881 12764 3893 12767
rect 3384 12736 3893 12764
rect 3384 12724 3390 12736
rect 3881 12733 3893 12736
rect 3927 12733 3939 12767
rect 3881 12727 3939 12733
rect 4062 12724 4068 12776
rect 4120 12724 4126 12776
rect 4341 12767 4399 12773
rect 4341 12733 4353 12767
rect 4387 12764 4399 12767
rect 4430 12764 4436 12776
rect 4387 12736 4436 12764
rect 4387 12733 4399 12736
rect 4341 12727 4399 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4614 12724 4620 12776
rect 4672 12764 4678 12776
rect 6196 12764 6224 12872
rect 12342 12860 12348 12912
rect 12400 12900 12406 12912
rect 13722 12900 13728 12912
rect 12400 12872 13728 12900
rect 12400 12860 12406 12872
rect 13722 12860 13728 12872
rect 13780 12860 13786 12912
rect 15010 12900 15016 12912
rect 14200 12872 15016 12900
rect 14200 12871 14228 12872
rect 14167 12865 14228 12871
rect 6270 12792 6276 12844
rect 6328 12832 6334 12844
rect 6607 12835 6665 12841
rect 6607 12832 6619 12835
rect 6328 12804 6619 12832
rect 6328 12792 6334 12804
rect 6607 12801 6619 12804
rect 6653 12832 6665 12835
rect 7282 12832 7288 12844
rect 6653 12804 7288 12832
rect 6653 12801 6665 12804
rect 6607 12795 6665 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 8018 12832 8024 12844
rect 7760 12804 8024 12832
rect 4672 12736 6224 12764
rect 6365 12767 6423 12773
rect 4672 12724 4678 12736
rect 6365 12733 6377 12767
rect 6411 12733 6423 12767
rect 6365 12727 6423 12733
rect 2280 12668 2360 12696
rect 3252 12668 3464 12696
rect 2280 12656 2286 12668
rect 2038 12588 2044 12640
rect 2096 12628 2102 12640
rect 3252 12628 3280 12668
rect 2096 12600 3280 12628
rect 2096 12588 2102 12600
rect 3326 12588 3332 12640
rect 3384 12588 3390 12640
rect 3436 12628 3464 12668
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 6380 12696 6408 12727
rect 6144 12668 6408 12696
rect 6144 12656 6150 12668
rect 7098 12656 7104 12708
rect 7156 12696 7162 12708
rect 7377 12699 7435 12705
rect 7377 12696 7389 12699
rect 7156 12668 7389 12696
rect 7156 12656 7162 12668
rect 7377 12665 7389 12668
rect 7423 12665 7435 12699
rect 7377 12659 7435 12665
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 3436 12600 5549 12628
rect 5537 12597 5549 12600
rect 5583 12597 5595 12631
rect 5537 12591 5595 12597
rect 6270 12588 6276 12640
rect 6328 12628 6334 12640
rect 7760 12628 7788 12804
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 9030 12792 9036 12844
rect 9088 12841 9094 12844
rect 9088 12835 9116 12841
rect 9104 12801 9116 12835
rect 9088 12795 9116 12801
rect 9088 12792 9094 12795
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 10319 12835 10377 12841
rect 10319 12801 10331 12835
rect 10365 12832 10377 12835
rect 10410 12832 10416 12844
rect 10365 12804 10416 12832
rect 10365 12801 10377 12804
rect 10319 12795 10377 12801
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 11606 12792 11612 12844
rect 11664 12792 11670 12844
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 11975 12835 12033 12841
rect 11975 12832 11987 12835
rect 11940 12804 11987 12832
rect 11940 12792 11946 12804
rect 11975 12801 11987 12804
rect 12021 12801 12033 12835
rect 14167 12832 14179 12865
rect 11975 12795 12033 12801
rect 12406 12831 14179 12832
rect 14213 12831 14228 12865
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 17034 12871 17040 12912
rect 17019 12865 17040 12871
rect 12406 12804 14228 12831
rect 17019 12831 17031 12865
rect 17092 12860 17098 12912
rect 19334 12900 19340 12912
rect 18248 12872 19340 12900
rect 17065 12834 17078 12860
rect 17065 12831 17077 12834
rect 17019 12825 17077 12831
rect 7834 12724 7840 12776
rect 7892 12724 7898 12776
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8754 12764 8760 12776
rect 8444 12736 8760 12764
rect 8444 12724 8450 12736
rect 8754 12724 8760 12736
rect 8812 12764 8818 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8812 12736 8953 12764
rect 8812 12724 8818 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12733 10103 12767
rect 11624 12764 11652 12792
rect 10045 12727 10103 12733
rect 10704 12736 11652 12764
rect 11701 12767 11759 12773
rect 7852 12696 7880 12724
rect 8665 12699 8723 12705
rect 8665 12696 8677 12699
rect 7852 12668 8677 12696
rect 8665 12665 8677 12668
rect 8711 12665 8723 12699
rect 8665 12659 8723 12665
rect 6328 12600 7788 12628
rect 6328 12588 6334 12600
rect 8294 12588 8300 12640
rect 8352 12628 8358 12640
rect 8754 12628 8760 12640
rect 8352 12600 8760 12628
rect 8352 12588 8358 12600
rect 8754 12588 8760 12600
rect 8812 12588 8818 12640
rect 9306 12588 9312 12640
rect 9364 12628 9370 12640
rect 10060 12628 10088 12727
rect 10704 12628 10732 12736
rect 11701 12733 11713 12767
rect 11747 12733 11759 12767
rect 11701 12727 11759 12733
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 11716 12696 11744 12727
rect 11296 12668 11744 12696
rect 11296 12656 11302 12668
rect 9364 12600 10732 12628
rect 9364 12588 9370 12600
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 12406 12628 12434 12804
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18248 12841 18276 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 21174 12900 21180 12912
rect 19628 12872 21180 12900
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 18012 12804 18245 12832
rect 18012 12792 18018 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18507 12835 18565 12841
rect 18507 12801 18519 12835
rect 18553 12832 18565 12835
rect 18598 12832 18604 12844
rect 18553 12804 18604 12832
rect 18553 12801 18565 12804
rect 18507 12795 18565 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 19628 12841 19656 12872
rect 21174 12860 21180 12872
rect 21232 12860 21238 12912
rect 22370 12900 22376 12912
rect 21284 12872 22376 12900
rect 21284 12841 21312 12872
rect 22370 12860 22376 12872
rect 22428 12860 22434 12912
rect 22664 12871 22692 12928
rect 22631 12865 22692 12871
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19880 12835 19938 12841
rect 19880 12801 19892 12835
rect 19926 12832 19938 12835
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 19926 12804 21281 12832
rect 19926 12801 19938 12804
rect 19880 12795 19938 12801
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 21545 12835 21603 12841
rect 21545 12801 21557 12835
rect 21591 12801 21603 12835
rect 21545 12795 21603 12801
rect 22097 12835 22155 12841
rect 22097 12801 22109 12835
rect 22143 12801 22155 12835
rect 22097 12795 22155 12801
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 13909 12767 13967 12773
rect 13909 12764 13921 12767
rect 13872 12736 13921 12764
rect 13872 12724 13878 12736
rect 13909 12733 13921 12736
rect 13955 12733 13967 12767
rect 13909 12727 13967 12733
rect 16761 12767 16819 12773
rect 16761 12733 16773 12767
rect 16807 12733 16819 12767
rect 21560 12764 21588 12795
rect 16761 12727 16819 12733
rect 21008 12736 21588 12764
rect 11020 12600 12434 12628
rect 11020 12588 11026 12600
rect 12710 12588 12716 12640
rect 12768 12588 12774 12640
rect 14918 12588 14924 12640
rect 14976 12588 14982 12640
rect 16776 12628 16804 12727
rect 19242 12656 19248 12708
rect 19300 12656 19306 12708
rect 21008 12705 21036 12736
rect 22112 12708 22140 12795
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 22631 12831 22643 12865
rect 22677 12832 22692 12865
rect 23937 12903 23995 12909
rect 23937 12869 23949 12903
rect 23983 12900 23995 12903
rect 24394 12900 24400 12912
rect 23983 12872 24400 12900
rect 23983 12869 23995 12872
rect 23937 12863 23995 12869
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 22677 12831 23060 12832
rect 22631 12825 23060 12831
rect 22664 12804 23060 12825
rect 22204 12764 22232 12792
rect 22373 12767 22431 12773
rect 22373 12764 22385 12767
rect 22204 12736 22385 12764
rect 20993 12699 21051 12705
rect 20993 12665 21005 12699
rect 21039 12665 21051 12699
rect 20993 12659 21051 12665
rect 22094 12656 22100 12708
rect 22152 12656 22158 12708
rect 17126 12628 17132 12640
rect 16776 12600 17132 12628
rect 17126 12588 17132 12600
rect 17184 12588 17190 12640
rect 17770 12588 17776 12640
rect 17828 12588 17834 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 21085 12631 21143 12637
rect 21085 12628 21097 12631
rect 20404 12600 21097 12628
rect 20404 12588 20410 12600
rect 21085 12597 21097 12600
rect 21131 12597 21143 12631
rect 21085 12591 21143 12597
rect 21450 12588 21456 12640
rect 21508 12628 21514 12640
rect 22204 12628 22232 12736
rect 22373 12733 22385 12736
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 21508 12600 22232 12628
rect 21508 12588 21514 12600
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 23032 12628 23060 12804
rect 22704 12600 23060 12628
rect 22704 12588 22710 12600
rect 24210 12588 24216 12640
rect 24268 12588 24274 12640
rect 1104 12538 24840 12560
rect 1104 12486 3917 12538
rect 3969 12486 3981 12538
rect 4033 12486 4045 12538
rect 4097 12486 4109 12538
rect 4161 12486 4173 12538
rect 4225 12486 9851 12538
rect 9903 12486 9915 12538
rect 9967 12486 9979 12538
rect 10031 12486 10043 12538
rect 10095 12486 10107 12538
rect 10159 12486 15785 12538
rect 15837 12486 15849 12538
rect 15901 12486 15913 12538
rect 15965 12486 15977 12538
rect 16029 12486 16041 12538
rect 16093 12486 21719 12538
rect 21771 12486 21783 12538
rect 21835 12486 21847 12538
rect 21899 12486 21911 12538
rect 21963 12486 21975 12538
rect 22027 12486 24840 12538
rect 1104 12464 24840 12486
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3568 12396 3985 12424
rect 3568 12384 3574 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 5994 12424 6000 12436
rect 3973 12387 4031 12393
rect 5552 12396 6000 12424
rect 4982 12316 4988 12368
rect 5040 12356 5046 12368
rect 5552 12365 5580 12396
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 9766 12424 9772 12436
rect 7024 12396 9772 12424
rect 5537 12359 5595 12365
rect 5040 12328 5488 12356
rect 5040 12316 5046 12328
rect 5460 12300 5488 12328
rect 5537 12325 5549 12359
rect 5583 12325 5595 12359
rect 5537 12319 5595 12325
rect 6748 12328 6960 12356
rect 1302 12248 1308 12300
rect 1360 12288 1366 12300
rect 1765 12291 1823 12297
rect 1765 12288 1777 12291
rect 1360 12260 1777 12288
rect 1360 12248 1366 12260
rect 1765 12257 1777 12260
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1949 12291 2007 12297
rect 1949 12257 1961 12291
rect 1995 12288 2007 12291
rect 2130 12288 2136 12300
rect 1995 12260 2136 12288
rect 1995 12257 2007 12260
rect 1949 12251 2007 12257
rect 1964 12084 1992 12251
rect 2130 12248 2136 12260
rect 2188 12248 2194 12300
rect 2406 12248 2412 12300
rect 2464 12248 2470 12300
rect 2498 12248 2504 12300
rect 2556 12288 2562 12300
rect 2866 12297 2872 12300
rect 2685 12291 2743 12297
rect 2685 12288 2697 12291
rect 2556 12260 2697 12288
rect 2556 12248 2562 12260
rect 2685 12257 2697 12260
rect 2731 12257 2743 12291
rect 2685 12251 2743 12257
rect 2823 12291 2872 12297
rect 2823 12257 2835 12291
rect 2869 12257 2872 12291
rect 2823 12251 2872 12257
rect 2866 12248 2872 12251
rect 2924 12248 2930 12300
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3326 12288 3332 12300
rect 3007 12260 3332 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3326 12248 3332 12260
rect 3384 12248 3390 12300
rect 3896 12260 5304 12288
rect 3896 12229 3924 12260
rect 5276 12232 5304 12260
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5500 12260 5825 12288
rect 5500 12248 5506 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6089 12291 6147 12297
rect 5960 12248 5973 12288
rect 6089 12257 6101 12291
rect 6135 12288 6147 12291
rect 6748 12288 6776 12328
rect 6932 12300 6960 12328
rect 6135 12260 6776 12288
rect 6135 12257 6147 12260
rect 6089 12251 6147 12257
rect 6822 12248 6828 12300
rect 6880 12248 6886 12300
rect 6914 12248 6920 12300
rect 6972 12248 6978 12300
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 4433 12223 4491 12229
rect 4433 12220 4445 12223
rect 4396 12192 4445 12220
rect 4396 12180 4402 12192
rect 4433 12189 4445 12192
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 4893 12223 4951 12229
rect 4893 12220 4905 12223
rect 4580 12192 4905 12220
rect 4580 12180 4586 12192
rect 4893 12189 4905 12192
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12189 5135 12223
rect 5077 12183 5135 12189
rect 5092 12152 5120 12183
rect 5258 12180 5264 12232
rect 5316 12180 5322 12232
rect 5945 12229 5973 12248
rect 7024 12229 7052 12396
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 21542 12384 21548 12436
rect 21600 12424 21606 12436
rect 22278 12424 22284 12436
rect 21600 12396 22284 12424
rect 21600 12384 21606 12396
rect 22278 12384 22284 12396
rect 22336 12384 22342 12436
rect 22649 12427 22707 12433
rect 22649 12393 22661 12427
rect 22695 12424 22707 12427
rect 24121 12427 24179 12433
rect 22695 12396 23428 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 7466 12316 7472 12368
rect 7524 12316 7530 12368
rect 15565 12359 15623 12365
rect 15565 12325 15577 12359
rect 15611 12356 15623 12359
rect 16298 12356 16304 12368
rect 15611 12328 16304 12356
rect 15611 12325 15623 12328
rect 15565 12319 15623 12325
rect 16298 12316 16304 12328
rect 16356 12356 16362 12368
rect 23293 12359 23351 12365
rect 16356 12328 17172 12356
rect 16356 12316 16362 12328
rect 12532 12300 12584 12306
rect 7208 12260 7788 12288
rect 7208 12232 7236 12260
rect 5945 12223 6009 12229
rect 5945 12189 5963 12223
rect 5997 12189 6009 12223
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 5945 12183 6009 12189
rect 6654 12192 7021 12220
rect 5945 12182 5994 12183
rect 3436 12124 5120 12152
rect 3436 12084 3464 12124
rect 1964 12056 3464 12084
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 3605 12087 3663 12093
rect 3605 12084 3617 12087
rect 3568 12056 3617 12084
rect 3568 12044 3574 12056
rect 3605 12053 3617 12056
rect 3651 12053 3663 12087
rect 3605 12047 3663 12053
rect 3694 12044 3700 12096
rect 3752 12084 3758 12096
rect 4525 12087 4583 12093
rect 4525 12084 4537 12087
rect 3752 12056 4537 12084
rect 3752 12044 3758 12056
rect 4525 12053 4537 12056
rect 4571 12053 4583 12087
rect 5092 12084 5120 12124
rect 5902 12084 5908 12096
rect 5092 12056 5908 12084
rect 4525 12047 4583 12053
rect 5902 12044 5908 12056
rect 5960 12084 5966 12096
rect 6654 12084 6682 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7190 12180 7196 12232
rect 7248 12180 7254 12232
rect 7760 12229 7788 12260
rect 7834 12248 7840 12300
rect 7892 12297 7898 12300
rect 7892 12291 7920 12297
rect 7908 12257 7920 12291
rect 7892 12251 7920 12257
rect 7892 12248 7898 12251
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 13964 12260 14122 12288
rect 13964 12248 13970 12260
rect 17034 12248 17040 12300
rect 17092 12248 17098 12300
rect 17144 12288 17172 12328
rect 23293 12325 23305 12359
rect 23339 12325 23351 12359
rect 23293 12319 23351 12325
rect 17430 12291 17488 12297
rect 17430 12288 17442 12291
rect 17144 12260 17442 12288
rect 17430 12257 17442 12260
rect 17476 12257 17488 12291
rect 17430 12251 17488 12257
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12288 17647 12291
rect 17770 12288 17776 12300
rect 17635 12260 17776 12288
rect 17635 12257 17647 12260
rect 17589 12251 17647 12257
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 12532 12242 12584 12248
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 11885 12223 11943 12229
rect 11885 12189 11897 12223
rect 11931 12220 11943 12223
rect 12710 12220 12716 12232
rect 11931 12210 12480 12220
rect 12636 12210 12716 12220
rect 11931 12192 12716 12210
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 12452 12182 12664 12192
rect 12710 12180 12716 12192
rect 12768 12180 12774 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 14458 12220 14464 12232
rect 12860 12192 14464 12220
rect 12860 12180 12866 12192
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 14645 12223 14703 12229
rect 14645 12189 14657 12223
rect 14691 12220 14703 12223
rect 14918 12220 14924 12232
rect 14691 12192 14924 12220
rect 14691 12189 14703 12192
rect 14645 12183 14703 12189
rect 14918 12180 14924 12192
rect 14976 12180 14982 12232
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 11793 12155 11851 12161
rect 9088 12124 11744 12152
rect 9088 12112 9094 12124
rect 5960 12056 6682 12084
rect 5960 12044 5966 12056
rect 6730 12044 6736 12096
rect 6788 12044 6794 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8665 12087 8723 12093
rect 8665 12084 8677 12087
rect 8352 12056 8677 12084
rect 8352 12044 8358 12056
rect 8665 12053 8677 12056
rect 8711 12053 8723 12087
rect 8665 12047 8723 12053
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12084 11575 12087
rect 11606 12084 11612 12096
rect 11563 12056 11612 12084
rect 11563 12053 11575 12056
rect 11517 12047 11575 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11716 12084 11744 12124
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 12158 12152 12164 12164
rect 11839 12124 12164 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 12253 12155 12311 12161
rect 12253 12121 12265 12155
rect 12299 12152 12311 12155
rect 12342 12152 12348 12164
rect 12299 12124 12348 12152
rect 12299 12121 12311 12124
rect 12253 12115 12311 12121
rect 12342 12112 12348 12124
rect 12400 12112 12406 12164
rect 12544 12124 12848 12152
rect 12544 12084 12572 12124
rect 11716 12056 12572 12084
rect 12618 12044 12624 12096
rect 12676 12044 12682 12096
rect 12820 12093 12848 12124
rect 13998 12112 14004 12164
rect 14056 12152 14062 12164
rect 14553 12155 14611 12161
rect 14553 12152 14565 12155
rect 14056 12124 14565 12152
rect 14056 12112 14062 12124
rect 14553 12121 14565 12124
rect 14599 12152 14611 12155
rect 14734 12152 14740 12164
rect 14599 12124 14740 12152
rect 14599 12121 14611 12124
rect 14553 12115 14611 12121
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 15013 12155 15071 12161
rect 15013 12121 15025 12155
rect 15059 12121 15071 12155
rect 15013 12115 15071 12121
rect 12805 12087 12863 12093
rect 12805 12053 12817 12087
rect 12851 12053 12863 12087
rect 12805 12047 12863 12053
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 14277 12087 14335 12093
rect 14277 12084 14289 12087
rect 14240 12056 14289 12084
rect 14240 12044 14246 12056
rect 14277 12053 14289 12056
rect 14323 12053 14335 12087
rect 14277 12047 14335 12053
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 15028 12084 15056 12115
rect 16408 12096 16436 12183
rect 16482 12180 16488 12232
rect 16540 12220 16546 12232
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 16540 12192 16589 12220
rect 16540 12180 16546 12192
rect 16577 12189 16589 12192
rect 16623 12220 16635 12223
rect 16758 12220 16764 12232
rect 16623 12192 16764 12220
rect 16623 12189 16635 12192
rect 16577 12183 16635 12189
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 20162 12229 20168 12232
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 20131 12223 20168 12229
rect 20131 12189 20143 12223
rect 20131 12183 20168 12189
rect 19904 12152 19932 12183
rect 20162 12180 20168 12183
rect 20220 12180 20226 12232
rect 21266 12180 21272 12232
rect 21324 12180 21330 12232
rect 22094 12220 22100 12232
rect 21376 12192 22100 12220
rect 20806 12152 20812 12164
rect 19904 12124 20812 12152
rect 20806 12112 20812 12124
rect 20864 12152 20870 12164
rect 21376 12152 21404 12192
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23308 12220 23336 12319
rect 23247 12192 23336 12220
rect 23400 12220 23428 12396
rect 24121 12393 24133 12427
rect 24167 12424 24179 12427
rect 25130 12424 25136 12436
rect 24167 12396 25136 12424
rect 24167 12393 24179 12396
rect 24121 12387 24179 12393
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 23753 12359 23811 12365
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 25222 12356 25228 12368
rect 23799 12328 25228 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 25222 12316 25228 12328
rect 25280 12316 25286 12368
rect 25682 12288 25688 12300
rect 23584 12260 25688 12288
rect 23584 12229 23612 12260
rect 25682 12248 25688 12260
rect 25740 12248 25746 12300
rect 23477 12223 23535 12229
rect 23477 12220 23489 12223
rect 23400 12192 23489 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23477 12189 23489 12192
rect 23523 12189 23535 12223
rect 23477 12183 23535 12189
rect 23569 12223 23627 12229
rect 23569 12189 23581 12223
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 20864 12124 21404 12152
rect 21536 12155 21594 12161
rect 20864 12112 20870 12124
rect 21536 12121 21548 12155
rect 21582 12152 21594 12155
rect 21634 12152 21640 12164
rect 21582 12124 21640 12152
rect 21582 12121 21594 12124
rect 21536 12115 21594 12121
rect 21634 12112 21640 12124
rect 21692 12112 21698 12164
rect 23032 12152 23060 12183
rect 23842 12180 23848 12232
rect 23900 12220 23906 12232
rect 23937 12223 23995 12229
rect 23937 12220 23949 12223
rect 23900 12192 23949 12220
rect 23900 12180 23906 12192
rect 23937 12189 23949 12192
rect 23983 12189 23995 12223
rect 23937 12183 23995 12189
rect 22066 12124 23060 12152
rect 14516 12056 15056 12084
rect 14516 12044 14522 12056
rect 15378 12044 15384 12096
rect 15436 12044 15442 12096
rect 16390 12044 16396 12096
rect 16448 12044 16454 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 16632 12056 18245 12084
rect 16632 12044 16638 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 20901 12087 20959 12093
rect 20901 12053 20913 12087
rect 20947 12084 20959 12087
rect 21818 12084 21824 12096
rect 20947 12056 21824 12084
rect 20947 12053 20959 12056
rect 20901 12047 20959 12053
rect 21818 12044 21824 12056
rect 21876 12084 21882 12096
rect 22066 12084 22094 12124
rect 21876 12056 22094 12084
rect 21876 12044 21882 12056
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 23106 12044 23112 12096
rect 23164 12044 23170 12096
rect 1104 11994 25000 12016
rect 1104 11942 6884 11994
rect 6936 11942 6948 11994
rect 7000 11942 7012 11994
rect 7064 11942 7076 11994
rect 7128 11942 7140 11994
rect 7192 11942 12818 11994
rect 12870 11942 12882 11994
rect 12934 11942 12946 11994
rect 12998 11942 13010 11994
rect 13062 11942 13074 11994
rect 13126 11942 18752 11994
rect 18804 11942 18816 11994
rect 18868 11942 18880 11994
rect 18932 11942 18944 11994
rect 18996 11942 19008 11994
rect 19060 11942 24686 11994
rect 24738 11942 24750 11994
rect 24802 11942 24814 11994
rect 24866 11942 24878 11994
rect 24930 11942 24942 11994
rect 24994 11942 25000 11994
rect 1104 11920 25000 11942
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 2869 11883 2927 11889
rect 2869 11880 2881 11883
rect 2464 11852 2881 11880
rect 2464 11840 2470 11852
rect 2869 11849 2881 11852
rect 2915 11849 2927 11883
rect 2869 11843 2927 11849
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 3694 11880 3700 11892
rect 3568 11852 3700 11880
rect 3568 11840 3574 11852
rect 3694 11840 3700 11852
rect 3752 11840 3758 11892
rect 4525 11883 4583 11889
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 4890 11880 4896 11892
rect 4571 11852 4896 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 5905 11883 5963 11889
rect 5905 11849 5917 11883
rect 5951 11880 5963 11883
rect 5994 11880 6000 11892
rect 5951 11852 6000 11880
rect 5951 11849 5963 11852
rect 5905 11843 5963 11849
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 7834 11880 7840 11892
rect 6932 11852 7840 11880
rect 3421 11771 3479 11777
rect 2131 11747 2189 11753
rect 2131 11713 2143 11747
rect 2177 11744 2189 11747
rect 2177 11716 2774 11744
rect 2177 11713 2189 11716
rect 2131 11707 2189 11713
rect 1857 11679 1915 11685
rect 1857 11645 1869 11679
rect 1903 11645 1915 11679
rect 2746 11676 2774 11716
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3421 11744 3433 11771
rect 3384 11737 3433 11744
rect 3467 11737 3479 11771
rect 3384 11731 3479 11737
rect 3384 11716 3464 11731
rect 3384 11704 3390 11716
rect 3510 11704 3516 11756
rect 3568 11704 3574 11756
rect 3787 11747 3845 11753
rect 3787 11713 3799 11747
rect 3833 11744 3845 11747
rect 3878 11744 3884 11756
rect 3833 11716 3884 11744
rect 3833 11713 3845 11716
rect 3787 11707 3845 11713
rect 3878 11704 3884 11716
rect 3936 11704 3942 11756
rect 5167 11747 5225 11753
rect 5167 11744 5179 11747
rect 4172 11716 5179 11744
rect 2746 11648 3372 11676
rect 1857 11639 1915 11645
rect 1872 11540 1900 11639
rect 2746 11580 3280 11608
rect 2222 11540 2228 11552
rect 1872 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2590 11500 2596 11552
rect 2648 11540 2654 11552
rect 2746 11540 2774 11580
rect 3252 11549 3280 11580
rect 2648 11512 2774 11540
rect 3237 11543 3295 11549
rect 2648 11500 2654 11512
rect 3237 11509 3249 11543
rect 3283 11509 3295 11543
rect 3344 11540 3372 11648
rect 4172 11540 4200 11716
rect 5167 11713 5179 11716
rect 5213 11744 5225 11747
rect 5258 11744 5264 11756
rect 5213 11716 5264 11744
rect 5213 11713 5225 11716
rect 5167 11707 5225 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 6932 11753 6960 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8018 11880 8024 11892
rect 7975 11852 8024 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 12526 11840 12532 11892
rect 12584 11840 12590 11892
rect 13906 11840 13912 11892
rect 13964 11840 13970 11892
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 16408 11852 16988 11880
rect 7282 11812 7288 11824
rect 7206 11784 7288 11812
rect 7206 11783 7234 11784
rect 7175 11777 7234 11783
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6880 11716 6929 11744
rect 6880 11704 6886 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 7175 11743 7187 11777
rect 7221 11746 7234 11777
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 8938 11772 8944 11824
rect 8996 11812 9002 11824
rect 12066 11812 12072 11824
rect 8996 11784 10732 11812
rect 8996 11772 9002 11784
rect 8297 11747 8355 11753
rect 7221 11743 7233 11746
rect 7175 11737 7233 11743
rect 6917 11707 6975 11713
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 4706 11636 4712 11688
rect 4764 11676 4770 11688
rect 4893 11679 4951 11685
rect 4893 11676 4905 11679
rect 4764 11648 4905 11676
rect 4764 11636 4770 11648
rect 4893 11645 4905 11648
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 8312 11608 8340 11707
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8571 11747 8629 11753
rect 8571 11744 8583 11747
rect 8536 11716 8583 11744
rect 8536 11704 8542 11716
rect 8571 11713 8583 11716
rect 8617 11713 8629 11747
rect 8571 11707 8629 11713
rect 8312 11580 8430 11608
rect 3344 11512 4200 11540
rect 3237 11503 3295 11509
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 8294 11540 8300 11552
rect 5408 11512 8300 11540
rect 5408 11500 5414 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8402 11540 8430 11580
rect 9122 11568 9128 11620
rect 9180 11608 9186 11620
rect 10594 11608 10600 11620
rect 9180 11580 10600 11608
rect 9180 11568 9186 11580
rect 10594 11568 10600 11580
rect 10652 11568 10658 11620
rect 8570 11540 8576 11552
rect 8402 11512 8576 11540
rect 8570 11500 8576 11512
rect 8628 11540 8634 11552
rect 8754 11540 8760 11552
rect 8628 11512 8760 11540
rect 8628 11500 8634 11512
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 9309 11543 9367 11549
rect 9309 11509 9321 11543
rect 9355 11540 9367 11543
rect 9674 11540 9680 11552
rect 9355 11512 9680 11540
rect 9355 11509 9367 11512
rect 9309 11503 9367 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 10704 11540 10732 11784
rect 11532 11784 12072 11812
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11532 11753 11560 11784
rect 12066 11772 12072 11784
rect 12124 11812 12130 11824
rect 12124 11784 12940 11812
rect 12124 11772 12130 11784
rect 12912 11753 12940 11784
rect 14550 11772 14556 11824
rect 14608 11812 14614 11824
rect 16408 11812 16436 11852
rect 16960 11812 16988 11852
rect 17402 11852 17693 11880
rect 17126 11812 17132 11824
rect 14608 11784 16436 11812
rect 14608 11772 14614 11784
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11296 11716 11529 11744
rect 11296 11704 11302 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11791 11747 11849 11753
rect 11791 11713 11803 11747
rect 11837 11744 11849 11747
rect 12897 11747 12955 11753
rect 11837 11716 12434 11744
rect 11837 11713 11849 11716
rect 11791 11707 11849 11713
rect 12406 11608 12434 11716
rect 12897 11713 12909 11747
rect 12943 11713 12955 11747
rect 12897 11707 12955 11713
rect 13171 11747 13229 11753
rect 13171 11713 13183 11747
rect 13217 11744 13229 11747
rect 13538 11744 13544 11756
rect 13217 11716 13544 11744
rect 13217 11713 13229 11716
rect 13171 11707 13229 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 14936 11753 14964 11784
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 15194 11744 15200 11756
rect 15155 11716 15200 11744
rect 14921 11707 14979 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 16408 11676 16436 11784
rect 16500 11784 16804 11812
rect 16960 11784 17132 11812
rect 16500 11756 16528 11784
rect 16482 11704 16488 11756
rect 16540 11704 16546 11756
rect 16776 11744 16804 11784
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 16850 11744 16856 11756
rect 16776 11716 16856 11744
rect 16850 11704 16856 11716
rect 16908 11753 16914 11756
rect 16908 11747 16969 11753
rect 16908 11713 16923 11747
rect 16957 11713 16969 11747
rect 16908 11707 16969 11713
rect 16908 11704 16914 11707
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17402 11744 17430 11852
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 17681 11843 17739 11849
rect 21453 11883 21511 11889
rect 21453 11849 21465 11883
rect 21499 11880 21511 11883
rect 22738 11880 22744 11892
rect 21499 11852 22744 11880
rect 21499 11849 21511 11852
rect 21453 11843 21511 11849
rect 22738 11840 22744 11852
rect 22796 11840 22802 11892
rect 22830 11840 22836 11892
rect 22888 11840 22894 11892
rect 23106 11840 23112 11892
rect 23164 11840 23170 11892
rect 23385 11883 23443 11889
rect 23385 11849 23397 11883
rect 23431 11880 23443 11883
rect 23474 11880 23480 11892
rect 23431 11852 23480 11880
rect 23431 11849 23443 11852
rect 23385 11843 23443 11849
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 22848 11812 22876 11840
rect 22388 11784 22876 11812
rect 17092 11716 17430 11744
rect 17092 11704 17098 11716
rect 17862 11704 17868 11756
rect 17920 11704 17926 11756
rect 17954 11704 17960 11756
rect 18012 11744 18018 11756
rect 18291 11747 18349 11753
rect 18291 11744 18303 11747
rect 18012 11716 18303 11744
rect 18012 11704 18018 11716
rect 18291 11713 18303 11716
rect 18337 11713 18349 11747
rect 18291 11707 18349 11713
rect 21634 11704 21640 11756
rect 21692 11704 21698 11756
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 22388 11753 22416 11784
rect 22373 11747 22431 11753
rect 21784 11716 22094 11744
rect 21784 11704 21790 11716
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16408 11648 16681 11676
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 17880 11676 17908 11704
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17880 11648 18061 11676
rect 16669 11639 16727 11645
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 21818 11636 21824 11688
rect 21876 11676 21882 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 21876 11648 21925 11676
rect 21876 11636 21882 11648
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 22066 11676 22094 11716
rect 22373 11713 22385 11747
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11744 22799 11747
rect 23124 11744 23152 11840
rect 23216 11784 23612 11812
rect 23216 11756 23244 11784
rect 22787 11716 23152 11744
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23198 11704 23204 11756
rect 23256 11704 23262 11756
rect 23293 11747 23351 11753
rect 23293 11713 23305 11747
rect 23339 11744 23351 11747
rect 23474 11744 23480 11756
rect 23339 11716 23480 11744
rect 23339 11713 23351 11716
rect 23293 11707 23351 11713
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 23584 11753 23612 11784
rect 23569 11747 23627 11753
rect 23569 11713 23581 11747
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 23661 11747 23719 11753
rect 23661 11713 23673 11747
rect 23707 11713 23719 11747
rect 23661 11707 23719 11713
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11713 24179 11747
rect 24121 11707 24179 11713
rect 23676 11676 23704 11707
rect 22066 11648 23704 11676
rect 21913 11639 21971 11645
rect 12894 11608 12900 11620
rect 12406 11580 12900 11608
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 15856 11580 16804 11608
rect 15856 11540 15884 11580
rect 10704 11512 15884 11540
rect 15933 11543 15991 11549
rect 15933 11509 15945 11543
rect 15979 11540 15991 11543
rect 16298 11540 16304 11552
rect 15979 11512 16304 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16776 11540 16804 11580
rect 19150 11568 19156 11620
rect 19208 11608 19214 11620
rect 22649 11611 22707 11617
rect 22649 11608 22661 11611
rect 19208 11580 22661 11608
rect 19208 11568 19214 11580
rect 22649 11577 22661 11580
rect 22695 11577 22707 11611
rect 22649 11571 22707 11577
rect 23109 11611 23167 11617
rect 23109 11577 23121 11611
rect 23155 11608 23167 11611
rect 24136 11608 24164 11707
rect 23155 11580 24164 11608
rect 23155 11577 23167 11580
rect 23109 11571 23167 11577
rect 18322 11540 18328 11552
rect 16776 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19058 11500 19064 11552
rect 19116 11500 19122 11552
rect 23842 11500 23848 11552
rect 23900 11500 23906 11552
rect 24397 11543 24455 11549
rect 24397 11509 24409 11543
rect 24443 11540 24455 11543
rect 25222 11540 25228 11552
rect 24443 11512 25228 11540
rect 24443 11509 24455 11512
rect 24397 11503 24455 11509
rect 25222 11500 25228 11512
rect 25280 11500 25286 11552
rect 1104 11450 24840 11472
rect 1104 11398 3917 11450
rect 3969 11398 3981 11450
rect 4033 11398 4045 11450
rect 4097 11398 4109 11450
rect 4161 11398 4173 11450
rect 4225 11398 9851 11450
rect 9903 11398 9915 11450
rect 9967 11398 9979 11450
rect 10031 11398 10043 11450
rect 10095 11398 10107 11450
rect 10159 11398 15785 11450
rect 15837 11398 15849 11450
rect 15901 11398 15913 11450
rect 15965 11398 15977 11450
rect 16029 11398 16041 11450
rect 16093 11398 21719 11450
rect 21771 11398 21783 11450
rect 21835 11398 21847 11450
rect 21899 11398 21911 11450
rect 21963 11398 21975 11450
rect 22027 11398 24840 11450
rect 1104 11376 24840 11398
rect 1762 11296 1768 11348
rect 1820 11296 1826 11348
rect 2314 11296 2320 11348
rect 2372 11296 2378 11348
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 3660 11308 4537 11336
rect 3660 11296 3666 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 5077 11339 5135 11345
rect 5077 11305 5089 11339
rect 5123 11305 5135 11339
rect 5077 11299 5135 11305
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 5092 11268 5120 11299
rect 6730 11296 6736 11348
rect 6788 11296 6794 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7524 11308 7665 11336
rect 7524 11296 7530 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 10042 11296 10048 11348
rect 10100 11336 10106 11348
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 10100 11308 17080 11336
rect 10100 11296 10106 11308
rect 3200 11240 5120 11268
rect 5445 11271 5503 11277
rect 3200 11228 3206 11240
rect 5445 11237 5457 11271
rect 5491 11237 5503 11271
rect 6748 11268 6776 11296
rect 9030 11268 9036 11280
rect 5445 11231 5503 11237
rect 5644 11240 6776 11268
rect 7300 11240 9036 11268
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 3605 11135 3663 11141
rect 2004 11104 3372 11132
rect 2004 11092 2010 11104
rect 474 11024 480 11076
rect 532 11064 538 11076
rect 1673 11067 1731 11073
rect 1673 11064 1685 11067
rect 532 11036 1685 11064
rect 532 11024 538 11036
rect 1673 11033 1685 11036
rect 1719 11033 1731 11067
rect 1673 11027 1731 11033
rect 2222 11024 2228 11076
rect 2280 11024 2286 11076
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2832 11036 2973 11064
rect 2832 11024 2838 11036
rect 2961 11033 2973 11036
rect 3007 11033 3019 11067
rect 3344 11064 3372 11104
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 4985 11135 5043 11141
rect 3651 11104 4936 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 3881 11067 3939 11073
rect 3881 11064 3893 11067
rect 3344 11036 3893 11064
rect 2961 11027 3019 11033
rect 3881 11033 3893 11036
rect 3927 11033 3939 11067
rect 3881 11027 3939 11033
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4433 11067 4491 11073
rect 4433 11064 4445 11067
rect 4304 11036 4445 11064
rect 4304 11024 4310 11036
rect 4433 11033 4445 11036
rect 4479 11033 4491 11067
rect 4908 11064 4936 11104
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5460 11132 5488 11231
rect 5644 11141 5672 11240
rect 5031 11104 5488 11132
rect 5629 11135 5687 11141
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 5629 11101 5641 11135
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11132 6699 11135
rect 6822 11132 6828 11144
rect 6687 11104 6828 11132
rect 6687 11101 6699 11104
rect 6641 11095 6699 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 6915 11135 6973 11141
rect 6915 11101 6927 11135
rect 6961 11132 6973 11135
rect 7006 11132 7012 11144
rect 6961 11104 7012 11132
rect 6961 11101 6973 11104
rect 6915 11095 6973 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7300 11064 7328 11240
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 12894 11228 12900 11280
rect 12952 11268 12958 11280
rect 15102 11268 15108 11280
rect 12952 11240 15108 11268
rect 12952 11228 12958 11240
rect 15102 11228 15108 11240
rect 15160 11228 15166 11280
rect 15746 11268 15752 11280
rect 15210 11240 15752 11268
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 9578 11203 9636 11209
rect 8987 11172 9352 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 9324 11144 9352 11172
rect 9578 11169 9590 11203
rect 9624 11200 9636 11203
rect 9674 11200 9680 11212
rect 9624 11172 9680 11200
rect 9624 11169 9636 11172
rect 9578 11163 9636 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 15210 11200 15238 11240
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 15838 11228 15844 11280
rect 15896 11228 15902 11280
rect 17052 11277 17080 11308
rect 17144 11308 18153 11336
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 9916 11172 15238 11200
rect 9916 11160 9922 11172
rect 16114 11160 16120 11212
rect 16172 11160 16178 11212
rect 16206 11160 16212 11212
rect 16264 11209 16270 11212
rect 16264 11203 16292 11209
rect 16280 11169 16292 11203
rect 16264 11163 16292 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11200 16451 11203
rect 17144 11200 17172 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 18380 11308 18736 11336
rect 18380 11296 18386 11308
rect 18708 11277 18736 11308
rect 19058 11296 19064 11348
rect 19116 11296 19122 11348
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 21082 11336 21088 11348
rect 19668 11308 21088 11336
rect 19668 11296 19674 11308
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 23198 11336 23204 11348
rect 22066 11308 23204 11336
rect 18693 11271 18751 11277
rect 18693 11237 18705 11271
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 16439 11172 17172 11200
rect 18877 11203 18935 11209
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 18877 11169 18889 11203
rect 18923 11200 18935 11203
rect 19076 11200 19104 11296
rect 18923 11172 19104 11200
rect 18923 11169 18935 11172
rect 18877 11163 18935 11169
rect 16264 11160 16270 11163
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 9122 11132 9128 11144
rect 7892 11104 9128 11132
rect 7892 11092 7898 11104
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9950 11092 9956 11144
rect 10008 11141 10014 11144
rect 10008 11135 10036 11141
rect 10024 11101 10036 11135
rect 10008 11095 10036 11101
rect 10008 11092 10014 11095
rect 10134 11092 10140 11144
rect 10192 11092 10198 11144
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15381 11135 15439 11141
rect 15381 11101 15393 11135
rect 15427 11101 15439 11135
rect 15381 11095 15439 11101
rect 4908 11036 7328 11064
rect 4433 11027 4491 11033
rect 8018 11024 8024 11076
rect 8076 11064 8082 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 8076 11036 9168 11064
rect 8076 11024 8082 11036
rect 1486 10956 1492 11008
rect 1544 10996 1550 11008
rect 2682 10996 2688 11008
rect 1544 10968 2688 10996
rect 1544 10956 1550 10968
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 3050 10956 3056 11008
rect 3108 10956 3114 11008
rect 3418 10956 3424 11008
rect 3476 10956 3482 11008
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 5350 10996 5356 11008
rect 4580 10968 5356 10996
rect 4580 10956 4586 10968
rect 5350 10956 5356 10968
rect 5408 10956 5414 11008
rect 7282 10956 7288 11008
rect 7340 10996 7346 11008
rect 8110 10996 8116 11008
rect 7340 10968 8116 10996
rect 7340 10956 7346 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 9140 10996 9168 11036
rect 10612 11036 10793 11064
rect 10612 10996 10640 11036
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 14918 11064 14924 11076
rect 12584 11036 14924 11064
rect 12584 11024 12590 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 9140 10968 10640 10996
rect 15396 10996 15424 11095
rect 17126 11092 17132 11144
rect 17184 11092 17190 11144
rect 17402 11132 17408 11144
rect 17363 11104 17408 11132
rect 17402 11092 17408 11104
rect 17460 11132 17466 11144
rect 17770 11132 17776 11144
rect 17460 11104 17776 11132
rect 17460 11092 17466 11104
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 18693 11135 18751 11141
rect 18693 11132 18705 11135
rect 18656 11104 18705 11132
rect 18656 11092 18662 11104
rect 18693 11101 18705 11104
rect 18739 11101 18751 11135
rect 19076 11132 19104 11172
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19076 11104 19257 11132
rect 18693 11095 18751 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19886 11132 19892 11144
rect 19475 11104 19892 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 20254 11092 20260 11144
rect 20312 11092 20318 11144
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 19061 11067 19119 11073
rect 17092 11036 19012 11064
rect 17092 11024 17098 11036
rect 16850 10996 16856 11008
rect 15396 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 18984 10996 19012 11036
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 19337 11067 19395 11073
rect 19337 11064 19349 11067
rect 19107 11036 19349 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19337 11033 19349 11036
rect 19383 11033 19395 11067
rect 20993 11067 21051 11073
rect 20993 11064 21005 11067
rect 19337 11027 19395 11033
rect 19444 11036 21005 11064
rect 19444 10996 19472 11036
rect 20993 11033 21005 11036
rect 21039 11033 21051 11067
rect 20993 11027 21051 11033
rect 21358 11024 21364 11076
rect 21416 11064 21422 11076
rect 22066 11064 22094 11308
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 23474 11296 23480 11348
rect 23532 11336 23538 11348
rect 23753 11339 23811 11345
rect 23753 11336 23765 11339
rect 23532 11308 23765 11336
rect 23532 11296 23538 11308
rect 23753 11305 23765 11308
rect 23799 11305 23811 11339
rect 23753 11299 23811 11305
rect 22462 11092 22468 11144
rect 22520 11132 22526 11144
rect 22646 11132 22652 11144
rect 22520 11104 22652 11132
rect 22520 11092 22526 11104
rect 22646 11092 22652 11104
rect 22704 11092 22710 11144
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 21416 11036 22094 11064
rect 21416 11024 21422 11036
rect 22756 11008 22784 11095
rect 22922 11092 22928 11144
rect 22980 11132 22986 11144
rect 23015 11135 23073 11141
rect 23015 11132 23027 11135
rect 22980 11104 23027 11132
rect 22980 11092 22986 11104
rect 23015 11101 23027 11104
rect 23061 11101 23073 11135
rect 23015 11095 23073 11101
rect 18984 10968 19472 10996
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 22738 10996 22744 11008
rect 22336 10968 22744 10996
rect 22336 10956 22342 10968
rect 22738 10956 22744 10968
rect 22796 10956 22802 11008
rect 1104 10906 25000 10928
rect 1104 10854 6884 10906
rect 6936 10854 6948 10906
rect 7000 10854 7012 10906
rect 7064 10854 7076 10906
rect 7128 10854 7140 10906
rect 7192 10854 12818 10906
rect 12870 10854 12882 10906
rect 12934 10854 12946 10906
rect 12998 10854 13010 10906
rect 13062 10854 13074 10906
rect 13126 10854 18752 10906
rect 18804 10854 18816 10906
rect 18868 10854 18880 10906
rect 18932 10854 18944 10906
rect 18996 10854 19008 10906
rect 19060 10854 24686 10906
rect 24738 10854 24750 10906
rect 24802 10854 24814 10906
rect 24866 10854 24878 10906
rect 24930 10854 24942 10906
rect 24994 10854 25000 10906
rect 1104 10832 25000 10854
rect 1578 10752 1584 10804
rect 1636 10752 1642 10804
rect 2222 10752 2228 10804
rect 2280 10792 2286 10804
rect 3789 10795 3847 10801
rect 3789 10792 3801 10795
rect 2280 10764 3801 10792
rect 2280 10752 2286 10764
rect 3789 10761 3801 10764
rect 3835 10761 3847 10795
rect 3789 10755 3847 10761
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5810 10792 5816 10804
rect 4764 10764 5816 10792
rect 4764 10752 4770 10764
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6178 10752 6184 10804
rect 6236 10792 6242 10804
rect 6546 10792 6552 10804
rect 6236 10764 6552 10792
rect 6236 10752 6242 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7374 10752 7380 10804
rect 7432 10752 7438 10804
rect 9490 10752 9496 10804
rect 9548 10752 9554 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10192 10764 10241 10792
rect 10192 10752 10198 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10965 10795 11023 10801
rect 10965 10761 10977 10795
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 16206 10792 16212 10804
rect 14967 10764 16212 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 1486 10684 1492 10736
rect 1544 10684 1550 10736
rect 7392 10724 7420 10752
rect 9508 10724 9536 10752
rect 3896 10696 4090 10724
rect 2499 10669 2557 10675
rect 2130 10616 2136 10668
rect 2188 10616 2194 10668
rect 2499 10635 2511 10669
rect 2545 10656 2557 10669
rect 3896 10656 3924 10696
rect 2545 10635 3924 10656
rect 2499 10629 3924 10635
rect 2514 10628 3924 10629
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 4062 10656 4090 10696
rect 4862 10696 7420 10724
rect 9324 10696 9536 10724
rect 4339 10659 4397 10665
rect 4339 10656 4351 10659
rect 4062 10628 4351 10656
rect 3973 10619 4031 10625
rect 4339 10625 4351 10628
rect 4385 10656 4397 10659
rect 4862 10656 4890 10696
rect 4385 10628 4890 10656
rect 4385 10625 4397 10628
rect 4339 10619 4397 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2240 10520 2268 10551
rect 3237 10523 3295 10529
rect 2240 10492 2360 10520
rect 2332 10464 2360 10492
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3510 10520 3516 10532
rect 3283 10492 3516 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3510 10480 3516 10492
rect 3568 10480 3574 10532
rect 1946 10412 1952 10464
rect 2004 10412 2010 10464
rect 2314 10412 2320 10464
rect 2372 10412 2378 10464
rect 3988 10452 4016 10619
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5868 10628 6377 10656
rect 5868 10616 5874 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6639 10659 6697 10665
rect 6639 10656 6651 10659
rect 6604 10628 6651 10656
rect 6604 10616 6610 10628
rect 6639 10625 6651 10628
rect 6685 10625 6697 10659
rect 6639 10619 6697 10625
rect 8570 10616 8576 10668
rect 8628 10656 8634 10668
rect 9217 10659 9275 10665
rect 9217 10656 9229 10659
rect 8628 10628 9229 10656
rect 8628 10616 8634 10628
rect 9217 10625 9229 10628
rect 9263 10656 9275 10659
rect 9324 10656 9352 10696
rect 9582 10684 9588 10736
rect 9640 10724 9646 10736
rect 10980 10724 11008 10755
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 19058 10792 19064 10804
rect 16298 10764 19064 10792
rect 9640 10696 11008 10724
rect 9640 10684 9646 10696
rect 13630 10684 13636 10736
rect 13688 10724 13694 10736
rect 14182 10724 14188 10736
rect 13688 10696 14188 10724
rect 13688 10684 13694 10696
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 14737 10727 14795 10733
rect 14737 10693 14749 10727
rect 14783 10693 14795 10727
rect 14737 10687 14795 10693
rect 9263 10628 9352 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9491 10659 9549 10665
rect 9491 10656 9503 10659
rect 9456 10628 9503 10656
rect 9456 10616 9462 10628
rect 9491 10625 9503 10628
rect 9537 10625 9549 10659
rect 9491 10619 9549 10625
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 11238 10656 11244 10668
rect 10827 10628 11244 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11882 10656 11888 10668
rect 11440 10628 11888 10656
rect 4062 10548 4068 10600
rect 4120 10548 4126 10600
rect 7558 10520 7564 10532
rect 4908 10492 6500 10520
rect 4908 10452 4936 10492
rect 3988 10424 4936 10452
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 5077 10455 5135 10461
rect 5077 10452 5089 10455
rect 5040 10424 5089 10452
rect 5040 10412 5046 10424
rect 5077 10421 5089 10424
rect 5123 10421 5135 10455
rect 6472 10452 6500 10492
rect 7300 10492 7564 10520
rect 7300 10452 7328 10492
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 6472 10424 7328 10452
rect 5077 10415 5135 10421
rect 7374 10412 7380 10464
rect 7432 10412 7438 10464
rect 7466 10412 7472 10464
rect 7524 10452 7530 10464
rect 11440 10452 11468 10628
rect 11882 10616 11888 10628
rect 11940 10656 11946 10668
rect 12311 10659 12369 10665
rect 12311 10656 12323 10659
rect 11940 10628 12323 10656
rect 11940 10616 11946 10628
rect 12311 10625 12323 10628
rect 12357 10625 12369 10659
rect 12311 10619 12369 10625
rect 13906 10616 13912 10668
rect 13964 10616 13970 10668
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 14369 10659 14427 10665
rect 14369 10656 14381 10659
rect 14332 10628 14381 10656
rect 14332 10616 14338 10628
rect 14369 10625 14381 10628
rect 14415 10656 14427 10659
rect 14458 10656 14464 10668
rect 14415 10628 14464 10656
rect 14415 10625 14427 10628
rect 14369 10619 14427 10625
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 14752 10656 14780 10687
rect 15746 10684 15752 10736
rect 15804 10724 15810 10736
rect 16298 10724 16326 10764
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19426 10792 19432 10804
rect 19168 10764 19432 10792
rect 19168 10724 19196 10764
rect 19426 10752 19432 10764
rect 19484 10752 19490 10804
rect 20070 10752 20076 10804
rect 20128 10792 20134 10804
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 20128 10764 20269 10792
rect 20128 10752 20134 10764
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 15804 10696 16326 10724
rect 17788 10696 19196 10724
rect 15804 10684 15810 10696
rect 14918 10656 14924 10668
rect 14752 10628 14924 10656
rect 14918 10616 14924 10628
rect 14976 10656 14982 10668
rect 15378 10656 15384 10668
rect 14976 10628 15384 10656
rect 14976 10616 14982 10628
rect 15378 10616 15384 10628
rect 15436 10616 15442 10668
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16298 10656 16304 10668
rect 15896 10628 16304 10656
rect 15896 10616 15902 10628
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 17788 10665 17816 10696
rect 19334 10686 19340 10698
rect 19260 10665 19340 10686
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10625 17739 10659
rect 17681 10619 17739 10625
rect 17773 10659 17831 10665
rect 17773 10625 17785 10659
rect 17819 10625 17831 10659
rect 18040 10659 18098 10665
rect 18040 10656 18052 10659
rect 17773 10619 17831 10625
rect 17880 10628 18052 10656
rect 11514 10548 11520 10600
rect 11572 10588 11578 10600
rect 12066 10588 12072 10600
rect 11572 10560 12072 10588
rect 11572 10548 11578 10560
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 13081 10523 13139 10529
rect 13081 10489 13093 10523
rect 13127 10520 13139 10523
rect 13464 10520 13492 10574
rect 15194 10548 15200 10600
rect 15252 10588 15258 10600
rect 16390 10588 16396 10600
rect 15252 10560 16396 10588
rect 15252 10548 15258 10560
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 17696 10588 17724 10619
rect 17880 10588 17908 10628
rect 18040 10625 18052 10628
rect 18086 10656 18098 10659
rect 19245 10659 19340 10665
rect 19245 10656 19257 10659
rect 18086 10628 19012 10656
rect 18086 10625 18098 10628
rect 18040 10619 18098 10625
rect 17696 10560 17908 10588
rect 13127 10492 13492 10520
rect 18984 10520 19012 10628
rect 19076 10628 19257 10656
rect 19076 10600 19104 10628
rect 19245 10625 19257 10628
rect 19291 10658 19340 10659
rect 19291 10625 19303 10658
rect 19334 10646 19340 10658
rect 19392 10646 19398 10698
rect 19509 10656 19515 10668
rect 19567 10665 19573 10668
rect 19477 10628 19515 10656
rect 19245 10619 19303 10625
rect 19509 10616 19515 10628
rect 19567 10619 19577 10665
rect 20272 10656 20300 10755
rect 20714 10752 20720 10804
rect 20772 10752 20778 10804
rect 20901 10795 20959 10801
rect 20901 10761 20913 10795
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 20625 10659 20683 10665
rect 20625 10656 20637 10659
rect 20272 10628 20637 10656
rect 20625 10625 20637 10628
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 19567 10616 19573 10619
rect 20714 10616 20720 10668
rect 20772 10616 20778 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 20916 10656 20944 10755
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 22646 10792 22652 10804
rect 22428 10764 22652 10792
rect 22428 10752 22434 10764
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 21192 10696 23026 10724
rect 20855 10628 20944 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 19058 10548 19064 10600
rect 19116 10548 19122 10600
rect 20732 10588 20760 10616
rect 21192 10588 21220 10696
rect 22998 10665 23026 10696
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10625 22707 10659
rect 22649 10619 22707 10625
rect 22983 10659 23041 10665
rect 22983 10625 22995 10659
rect 23029 10625 23041 10659
rect 22983 10619 23041 10625
rect 20732 10560 21220 10588
rect 18984 10492 19288 10520
rect 13127 10489 13139 10492
rect 13081 10483 13139 10489
rect 7524 10424 11468 10452
rect 7524 10412 7530 10424
rect 17494 10412 17500 10464
rect 17552 10412 17558 10464
rect 19150 10412 19156 10464
rect 19208 10412 19214 10464
rect 19260 10452 19288 10492
rect 19334 10452 19340 10464
rect 19260 10424 19340 10452
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22428 10424 22477 10452
rect 22428 10412 22434 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 22664 10452 22692 10619
rect 22738 10548 22744 10600
rect 22796 10548 22802 10600
rect 23753 10455 23811 10461
rect 23753 10452 23765 10455
rect 22664 10424 23765 10452
rect 22465 10415 22523 10421
rect 23753 10421 23765 10424
rect 23799 10421 23811 10455
rect 23753 10415 23811 10421
rect 1104 10362 24840 10384
rect 1104 10310 3917 10362
rect 3969 10310 3981 10362
rect 4033 10310 4045 10362
rect 4097 10310 4109 10362
rect 4161 10310 4173 10362
rect 4225 10310 9851 10362
rect 9903 10310 9915 10362
rect 9967 10310 9979 10362
rect 10031 10310 10043 10362
rect 10095 10310 10107 10362
rect 10159 10310 15785 10362
rect 15837 10310 15849 10362
rect 15901 10310 15913 10362
rect 15965 10310 15977 10362
rect 16029 10310 16041 10362
rect 16093 10310 21719 10362
rect 21771 10310 21783 10362
rect 21835 10310 21847 10362
rect 21899 10310 21911 10362
rect 21963 10310 21975 10362
rect 22027 10310 24840 10362
rect 1104 10288 24840 10310
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2556 10220 4568 10248
rect 2556 10208 2562 10220
rect 382 10072 388 10124
rect 440 10112 446 10124
rect 1765 10115 1823 10121
rect 1765 10112 1777 10115
rect 440 10084 1777 10112
rect 440 10072 446 10084
rect 1765 10081 1777 10084
rect 1811 10081 1823 10115
rect 1765 10075 1823 10081
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2038 10112 2044 10124
rect 1995 10084 2044 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2038 10072 2044 10084
rect 2096 10072 2102 10124
rect 2406 10072 2412 10124
rect 2464 10072 2470 10124
rect 2516 10112 2544 10208
rect 3804 10152 4384 10180
rect 2685 10115 2743 10121
rect 2685 10112 2697 10115
rect 2516 10084 2697 10112
rect 2685 10081 2697 10084
rect 2731 10081 2743 10115
rect 2685 10075 2743 10081
rect 2961 10115 3019 10121
rect 2961 10081 2973 10115
rect 3007 10112 3019 10115
rect 3510 10112 3516 10124
rect 3007 10084 3516 10112
rect 3007 10081 3019 10084
rect 2961 10075 3019 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 2866 10053 2872 10056
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 2823 10047 2872 10053
rect 2823 10013 2835 10047
rect 2869 10013 2872 10047
rect 2823 10007 2872 10013
rect 1486 9868 1492 9920
rect 1544 9868 1550 9920
rect 1688 9908 1716 10007
rect 2866 10004 2872 10007
rect 2924 10004 2930 10056
rect 3804 10053 3832 10152
rect 4356 10124 4384 10152
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 4430 10072 4436 10124
rect 4488 10072 4494 10124
rect 4540 10112 4568 10220
rect 7374 10208 7380 10260
rect 7432 10208 7438 10260
rect 7558 10208 7564 10260
rect 7616 10208 7622 10260
rect 11514 10248 11520 10260
rect 9968 10220 11520 10248
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 5592 10152 6500 10180
rect 5592 10140 5598 10152
rect 4890 10121 4896 10124
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 4540 10084 4721 10112
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 4847 10115 4896 10121
rect 4847 10081 4859 10115
rect 4893 10081 4896 10115
rect 4847 10075 4896 10081
rect 4890 10072 4896 10075
rect 4948 10072 4954 10124
rect 4982 10072 4988 10124
rect 5040 10072 5046 10124
rect 5350 10072 5356 10124
rect 5408 10112 5414 10124
rect 5408 10084 5580 10112
rect 5408 10072 5414 10084
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 5552 10044 5580 10084
rect 5902 10072 5908 10124
rect 5960 10072 5966 10124
rect 6362 10072 6368 10124
rect 6420 10072 6426 10124
rect 6472 10112 6500 10152
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6472 10084 6653 10112
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6730 10072 6736 10124
rect 6788 10121 6794 10124
rect 6788 10115 6816 10121
rect 6804 10081 6816 10115
rect 6788 10075 6816 10081
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7392 10112 7420 10208
rect 9968 10121 9996 10220
rect 11514 10208 11520 10220
rect 11572 10208 11578 10260
rect 13998 10208 14004 10260
rect 14056 10248 14062 10260
rect 15105 10251 15163 10257
rect 15105 10248 15117 10251
rect 14056 10220 15117 10248
rect 14056 10208 14062 10220
rect 15105 10217 15117 10220
rect 15151 10217 15163 10251
rect 15105 10211 15163 10217
rect 17494 10208 17500 10260
rect 17552 10208 17558 10260
rect 18322 10208 18328 10260
rect 18380 10208 18386 10260
rect 18417 10251 18475 10257
rect 18417 10217 18429 10251
rect 18463 10248 18475 10251
rect 18598 10248 18604 10260
rect 18463 10220 18604 10248
rect 18463 10217 18475 10220
rect 18417 10211 18475 10217
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 19150 10208 19156 10260
rect 19208 10208 19214 10260
rect 19334 10208 19340 10260
rect 19392 10248 19398 10260
rect 19610 10248 19616 10260
rect 19392 10220 19616 10248
rect 19392 10208 19398 10220
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 20165 10251 20223 10257
rect 20165 10217 20177 10251
rect 20211 10248 20223 10251
rect 20254 10248 20260 10260
rect 20211 10220 20260 10248
rect 20211 10217 20223 10220
rect 20165 10211 20223 10217
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 10965 10183 11023 10189
rect 10965 10149 10977 10183
rect 11011 10149 11023 10183
rect 10965 10143 11023 10149
rect 6963 10084 7420 10112
rect 9953 10115 10011 10121
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 9953 10081 9965 10115
rect 9999 10081 10011 10115
rect 10980 10112 11008 10143
rect 10980 10084 11362 10112
rect 9953 10075 10011 10081
rect 6788 10072 6794 10075
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5552 10016 5733 10044
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 11698 10044 11704 10056
rect 5721 10007 5779 10013
rect 10210 10017 11704 10044
rect 10210 9983 10223 10017
rect 10257 10016 11704 10017
rect 10257 9983 10269 10016
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12618 10044 12624 10056
rect 11931 10016 12624 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 14056 10016 14105 10044
rect 14056 10004 14062 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14367 10047 14425 10053
rect 14367 10044 14379 10047
rect 14093 10007 14151 10013
rect 14182 10016 14379 10044
rect 10210 9977 10269 9983
rect 10210 9976 10238 9977
rect 9600 9948 10238 9976
rect 9600 9920 9628 9948
rect 10410 9936 10416 9988
rect 10468 9976 10474 9988
rect 10962 9976 10968 9988
rect 10468 9948 10968 9976
rect 10468 9936 10474 9948
rect 10962 9936 10968 9948
rect 11020 9976 11026 9988
rect 11793 9979 11851 9985
rect 11020 9948 11744 9976
rect 11020 9936 11026 9948
rect 3605 9911 3663 9917
rect 3605 9908 3617 9911
rect 1688 9880 3617 9908
rect 3605 9877 3617 9880
rect 3651 9877 3663 9911
rect 3605 9871 3663 9877
rect 5626 9868 5632 9920
rect 5684 9868 5690 9920
rect 5810 9868 5816 9920
rect 5868 9908 5874 9920
rect 8478 9908 8484 9920
rect 5868 9880 8484 9908
rect 5868 9868 5874 9880
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11606 9908 11612 9920
rect 11563 9880 11612 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 11716 9908 11744 9948
rect 11793 9945 11805 9979
rect 11839 9976 11851 9979
rect 11974 9976 11980 9988
rect 11839 9948 11980 9976
rect 11839 9945 11851 9948
rect 11793 9939 11851 9945
rect 11974 9936 11980 9948
rect 12032 9976 12038 9988
rect 12158 9976 12164 9988
rect 12032 9948 12164 9976
rect 12032 9936 12038 9948
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 12253 9979 12311 9985
rect 12253 9945 12265 9979
rect 12299 9976 12311 9979
rect 12342 9976 12348 9988
rect 12299 9948 12348 9976
rect 12299 9945 12311 9948
rect 12253 9939 12311 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 12452 9948 12848 9976
rect 12452 9908 12480 9948
rect 11716 9880 12480 9908
rect 12621 9911 12679 9917
rect 12621 9877 12633 9911
rect 12667 9908 12679 9911
rect 12710 9908 12716 9920
rect 12667 9880 12716 9908
rect 12667 9877 12679 9880
rect 12621 9871 12679 9877
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 12820 9917 12848 9948
rect 13722 9936 13728 9988
rect 13780 9976 13786 9988
rect 14182 9976 14210 10016
rect 14367 10013 14379 10016
rect 14413 10044 14425 10047
rect 17512 10044 17540 10208
rect 18340 10180 18368 10208
rect 19058 10180 19064 10192
rect 18340 10152 19064 10180
rect 19058 10140 19064 10152
rect 19116 10140 19122 10192
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 14413 10016 15792 10044
rect 17512 10016 18337 10044
rect 14413 10013 14425 10016
rect 14367 10007 14425 10013
rect 15764 9988 15792 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10044 19119 10047
rect 19168 10044 19196 10208
rect 20349 10183 20407 10189
rect 20349 10149 20361 10183
rect 20395 10149 20407 10183
rect 20349 10143 20407 10149
rect 19107 10016 19196 10044
rect 20073 10047 20131 10053
rect 19107 10013 19119 10016
rect 19061 10007 19119 10013
rect 20073 10013 20085 10047
rect 20119 10044 20131 10047
rect 20364 10044 20392 10143
rect 20806 10072 20812 10124
rect 20864 10072 20870 10124
rect 20119 10016 20392 10044
rect 20533 10047 20591 10053
rect 20119 10013 20131 10016
rect 20073 10007 20131 10013
rect 20533 10013 20545 10047
rect 20579 10044 20591 10047
rect 20579 10016 20668 10044
rect 20579 10013 20591 10016
rect 20533 10007 20591 10013
rect 13780 9948 14210 9976
rect 13780 9936 13786 9948
rect 15746 9936 15752 9988
rect 15804 9936 15810 9988
rect 20640 9920 20668 10016
rect 20824 9976 20852 10072
rect 21083 10047 21141 10053
rect 21083 10013 21095 10047
rect 21129 10044 21141 10047
rect 21174 10044 21180 10056
rect 21129 10016 21180 10044
rect 21129 10013 21141 10016
rect 21083 10007 21141 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 22738 10004 22744 10056
rect 22796 10004 22802 10056
rect 23014 10053 23020 10056
rect 22983 10047 23020 10053
rect 22983 10013 22995 10047
rect 22983 10007 23020 10013
rect 23014 10004 23020 10007
rect 23072 10004 23078 10056
rect 21450 9976 21456 9988
rect 20824 9948 21456 9976
rect 21450 9936 21456 9948
rect 21508 9936 21514 9988
rect 12805 9911 12863 9917
rect 12805 9877 12817 9911
rect 12851 9877 12863 9911
rect 12805 9871 12863 9877
rect 18877 9911 18935 9917
rect 18877 9877 18889 9911
rect 18923 9908 18935 9911
rect 19886 9908 19892 9920
rect 18923 9880 19892 9908
rect 18923 9877 18935 9880
rect 18877 9871 18935 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20622 9868 20628 9920
rect 20680 9868 20686 9920
rect 21174 9868 21180 9920
rect 21232 9908 21238 9920
rect 21542 9908 21548 9920
rect 21232 9880 21548 9908
rect 21232 9868 21238 9880
rect 21542 9868 21548 9880
rect 21600 9868 21606 9920
rect 21818 9868 21824 9920
rect 21876 9868 21882 9920
rect 22278 9868 22284 9920
rect 22336 9868 22342 9920
rect 23750 9868 23756 9920
rect 23808 9868 23814 9920
rect 1104 9818 25000 9840
rect 1104 9766 6884 9818
rect 6936 9766 6948 9818
rect 7000 9766 7012 9818
rect 7064 9766 7076 9818
rect 7128 9766 7140 9818
rect 7192 9766 12818 9818
rect 12870 9766 12882 9818
rect 12934 9766 12946 9818
rect 12998 9766 13010 9818
rect 13062 9766 13074 9818
rect 13126 9766 18752 9818
rect 18804 9766 18816 9818
rect 18868 9766 18880 9818
rect 18932 9766 18944 9818
rect 18996 9766 19008 9818
rect 19060 9766 24686 9818
rect 24738 9766 24750 9818
rect 24802 9766 24814 9818
rect 24866 9766 24878 9818
rect 24930 9766 24942 9818
rect 24994 9766 25000 9818
rect 1104 9744 25000 9766
rect 1578 9664 1584 9716
rect 1636 9664 1642 9716
rect 1780 9676 2360 9704
rect 1596 9601 1624 9664
rect 1581 9595 1639 9601
rect 1581 9561 1593 9595
rect 1627 9561 1639 9595
rect 1780 9578 1808 9676
rect 2332 9648 2360 9676
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 2685 9707 2743 9713
rect 2685 9704 2697 9707
rect 2464 9676 2697 9704
rect 2464 9664 2470 9676
rect 2685 9673 2697 9676
rect 2731 9673 2743 9707
rect 2685 9667 2743 9673
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3326 9704 3332 9716
rect 2924 9676 3332 9704
rect 2924 9664 2930 9676
rect 3326 9664 3332 9676
rect 3384 9664 3390 9716
rect 4430 9664 4436 9716
rect 4488 9704 4494 9716
rect 4525 9707 4583 9713
rect 4525 9704 4537 9707
rect 4488 9676 4537 9704
rect 4488 9664 4494 9676
rect 4525 9673 4537 9676
rect 4571 9673 4583 9707
rect 4525 9667 4583 9673
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6362 9704 6368 9716
rect 5951 9676 6368 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 10502 9704 10508 9716
rect 7668 9676 9168 9704
rect 2314 9596 2320 9648
rect 2372 9596 2378 9648
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 3418 9636 3424 9648
rect 2556 9608 3424 9636
rect 2556 9596 2562 9608
rect 3418 9596 3424 9608
rect 3476 9596 3482 9648
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 3878 9636 3884 9648
rect 3568 9608 3884 9636
rect 3568 9596 3574 9608
rect 3878 9596 3884 9608
rect 3936 9596 3942 9648
rect 1688 9577 1808 9578
rect 1581 9555 1639 9561
rect 1673 9571 1808 9577
rect 1673 9537 1685 9571
rect 1719 9550 1808 9571
rect 1947 9571 2005 9577
rect 1719 9537 1731 9550
rect 1673 9531 1731 9537
rect 1947 9537 1959 9571
rect 1993 9568 2005 9571
rect 2038 9568 2044 9580
rect 1993 9540 2044 9568
rect 1993 9537 2005 9540
rect 1947 9531 2005 9537
rect 2038 9528 2044 9540
rect 2096 9568 2102 9580
rect 2096 9540 2360 9568
rect 2096 9528 2102 9540
rect 2332 9500 2360 9540
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 3755 9571 3813 9577
rect 3755 9568 3767 9571
rect 3344 9540 3767 9568
rect 3344 9500 3372 9540
rect 3755 9537 3767 9540
rect 3801 9537 3813 9571
rect 3755 9531 3813 9537
rect 4338 9528 4344 9580
rect 4396 9568 4402 9580
rect 5074 9568 5080 9580
rect 4396 9540 5080 9568
rect 4396 9528 4402 9540
rect 5074 9528 5080 9540
rect 5132 9577 5138 9580
rect 5132 9571 5193 9577
rect 5132 9537 5147 9571
rect 5181 9537 5193 9571
rect 5132 9531 5193 9537
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7558 9568 7564 9580
rect 7515 9540 7564 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 5132 9528 5138 9531
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 2332 9472 3372 9500
rect 3510 9460 3516 9512
rect 3568 9460 3574 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 4893 9503 4951 9509
rect 4893 9500 4905 9503
rect 4764 9472 4905 9500
rect 4764 9460 4770 9472
rect 4893 9469 4905 9472
rect 4939 9469 4951 9503
rect 4893 9463 4951 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 7668 9509 7696 9676
rect 9140 9636 9168 9676
rect 9600 9676 10508 9704
rect 9600 9636 9628 9676
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 10744 9676 11100 9704
rect 10744 9664 10750 9676
rect 9140 9608 9628 9636
rect 11072 9636 11100 9676
rect 11238 9664 11244 9716
rect 11296 9664 11302 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12805 9707 12863 9713
rect 12805 9704 12817 9707
rect 12676 9676 12817 9704
rect 12676 9664 12682 9676
rect 12805 9673 12817 9676
rect 12851 9673 12863 9707
rect 12805 9667 12863 9673
rect 14366 9664 14372 9716
rect 14424 9704 14430 9716
rect 15194 9704 15200 9716
rect 14424 9676 15200 9704
rect 14424 9664 14430 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 20990 9704 20996 9716
rect 15804 9676 20996 9704
rect 15804 9664 15810 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 21082 9664 21088 9716
rect 21140 9664 21146 9716
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 21818 9704 21824 9716
rect 21600 9676 21824 9704
rect 21600 9664 21606 9676
rect 21818 9664 21824 9676
rect 21876 9704 21882 9716
rect 21876 9676 22140 9704
rect 21876 9664 21882 9676
rect 11514 9636 11520 9648
rect 11072 9608 11520 9636
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 7653 9503 7711 9509
rect 7653 9500 7665 9503
rect 6604 9472 7665 9500
rect 6604 9460 6610 9472
rect 7653 9469 7665 9472
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 8110 9460 8116 9512
rect 8168 9460 8174 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 8404 9500 8432 9531
rect 8662 9528 8668 9580
rect 8720 9528 8726 9580
rect 9600 9577 9628 9608
rect 11514 9596 11520 9608
rect 11572 9636 11578 9648
rect 17310 9636 17316 9648
rect 11572 9608 17316 9636
rect 11572 9596 11578 9608
rect 17310 9596 17316 9608
rect 17368 9596 17374 9648
rect 18138 9596 18144 9648
rect 18196 9636 18202 9648
rect 19972 9639 20030 9645
rect 18196 9608 18451 9636
rect 18196 9596 18202 9608
rect 9585 9571 9643 9577
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 10410 9528 10416 9580
rect 10468 9577 10474 9580
rect 10468 9571 10496 9577
rect 10484 9537 10496 9571
rect 10468 9531 10496 9537
rect 10468 9528 10474 9531
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 12067 9571 12125 9577
rect 12067 9568 12079 9571
rect 11164 9540 12079 9568
rect 8260 9472 8432 9500
rect 8527 9503 8585 9509
rect 8260 9460 8266 9472
rect 8527 9469 8539 9503
rect 8573 9500 8585 9503
rect 9030 9500 9036 9512
rect 8573 9472 9036 9500
rect 8573 9469 8585 9472
rect 8527 9463 8585 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9140 9472 9413 9500
rect 9140 9444 9168 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 10134 9500 10140 9512
rect 9732 9472 10140 9500
rect 9732 9460 9738 9472
rect 10134 9460 10140 9472
rect 10192 9460 10198 9512
rect 10321 9503 10379 9509
rect 10321 9469 10333 9503
rect 10367 9500 10379 9503
rect 10778 9500 10784 9512
rect 10367 9472 10784 9500
rect 10367 9469 10379 9472
rect 10321 9463 10379 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11164 9500 11192 9540
rect 12067 9537 12079 9540
rect 12113 9568 12125 9571
rect 16942 9568 16948 9580
rect 12113 9540 16948 9568
rect 12113 9537 12125 9540
rect 12067 9531 12125 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 18322 9528 18328 9580
rect 18380 9528 18386 9580
rect 18423 9568 18451 9608
rect 18583 9601 18641 9607
rect 18583 9568 18595 9601
rect 18423 9567 18595 9568
rect 18629 9567 18641 9601
rect 19972 9605 19984 9639
rect 20018 9636 20030 9639
rect 20622 9636 20628 9648
rect 20018 9608 20628 9636
rect 20018 9605 20030 9608
rect 19972 9599 20030 9605
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 22112 9577 22140 9676
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 22296 9577 22324 9664
rect 22830 9636 22836 9648
rect 22572 9608 22836 9636
rect 22572 9577 22600 9608
rect 22830 9596 22836 9608
rect 22888 9596 22894 9648
rect 18423 9561 18641 9567
rect 21821 9571 21879 9577
rect 18423 9540 18626 9561
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 21821 9531 21879 9537
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9537 22615 9571
rect 22983 9571 23041 9577
rect 22983 9568 22995 9571
rect 22557 9531 22615 9537
rect 22664 9540 22995 9568
rect 11020 9472 11192 9500
rect 11793 9503 11851 9509
rect 11020 9460 11026 9472
rect 11793 9469 11805 9503
rect 11839 9469 11851 9503
rect 11793 9463 11851 9469
rect 2746 9404 3188 9432
rect 1397 9367 1455 9373
rect 1397 9333 1409 9367
rect 1443 9364 1455 9367
rect 2746 9364 2774 9404
rect 1443 9336 2774 9364
rect 1443 9333 1455 9336
rect 1397 9327 1455 9333
rect 3050 9324 3056 9376
rect 3108 9324 3114 9376
rect 3160 9364 3188 9404
rect 9122 9392 9128 9444
rect 9180 9392 9186 9444
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9401 9367 9435
rect 9309 9395 9367 9401
rect 10045 9435 10103 9441
rect 10045 9401 10057 9435
rect 10091 9401 10103 9435
rect 10045 9395 10103 9401
rect 4246 9364 4252 9376
rect 3160 9336 4252 9364
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 5994 9324 6000 9376
rect 6052 9364 6058 9376
rect 9324 9364 9352 9395
rect 6052 9336 9352 9364
rect 10060 9364 10088 9395
rect 10318 9364 10324 9376
rect 10060 9336 10324 9364
rect 6052 9324 6058 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 11808 9364 11836 9463
rect 19702 9460 19708 9512
rect 19760 9460 19766 9512
rect 21836 9500 21864 9531
rect 21836 9472 22416 9500
rect 13998 9392 14004 9444
rect 14056 9432 14062 9444
rect 18138 9432 18144 9444
rect 14056 9404 18144 9432
rect 14056 9392 14062 9404
rect 18138 9392 18144 9404
rect 18196 9392 18202 9444
rect 22388 9441 22416 9472
rect 22373 9435 22431 9441
rect 18984 9404 19656 9432
rect 12158 9364 12164 9376
rect 11808 9336 12164 9364
rect 12158 9324 12164 9336
rect 12216 9364 12222 9376
rect 14016 9364 14044 9392
rect 12216 9336 14044 9364
rect 12216 9324 12222 9336
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 17126 9364 17132 9376
rect 15528 9336 17132 9364
rect 15528 9324 15534 9336
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17494 9324 17500 9376
rect 17552 9364 17558 9376
rect 18984 9364 19012 9404
rect 17552 9336 19012 9364
rect 19337 9367 19395 9373
rect 17552 9324 17558 9336
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19518 9364 19524 9376
rect 19383 9336 19524 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19628 9364 19656 9404
rect 20640 9404 22324 9432
rect 20640 9364 20668 9404
rect 19628 9336 20668 9364
rect 21913 9367 21971 9373
rect 21913 9333 21925 9367
rect 21959 9364 21971 9367
rect 22094 9364 22100 9376
rect 21959 9336 22100 9364
rect 21959 9333 21971 9336
rect 21913 9327 21971 9333
rect 22094 9324 22100 9336
rect 22152 9324 22158 9376
rect 22186 9324 22192 9376
rect 22244 9324 22250 9376
rect 22296 9364 22324 9404
rect 22373 9401 22385 9435
rect 22419 9401 22431 9435
rect 22373 9395 22431 9401
rect 22664 9364 22692 9540
rect 22983 9537 22995 9540
rect 23029 9537 23041 9571
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 22983 9531 23041 9537
rect 23768 9540 24317 9568
rect 22738 9460 22744 9512
rect 22796 9460 22802 9512
rect 22296 9336 22692 9364
rect 22756 9364 22784 9460
rect 23768 9441 23796 9540
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 24210 9460 24216 9512
rect 24268 9460 24274 9512
rect 23753 9435 23811 9441
rect 23753 9401 23765 9435
rect 23799 9401 23811 9435
rect 24228 9432 24256 9460
rect 23753 9395 23811 9401
rect 23860 9404 24256 9432
rect 23860 9364 23888 9404
rect 22756 9336 23888 9364
rect 24118 9324 24124 9376
rect 24176 9324 24182 9376
rect 1104 9274 24840 9296
rect 1104 9222 3917 9274
rect 3969 9222 3981 9274
rect 4033 9222 4045 9274
rect 4097 9222 4109 9274
rect 4161 9222 4173 9274
rect 4225 9222 9851 9274
rect 9903 9222 9915 9274
rect 9967 9222 9979 9274
rect 10031 9222 10043 9274
rect 10095 9222 10107 9274
rect 10159 9222 15785 9274
rect 15837 9222 15849 9274
rect 15901 9222 15913 9274
rect 15965 9222 15977 9274
rect 16029 9222 16041 9274
rect 16093 9222 21719 9274
rect 21771 9222 21783 9274
rect 21835 9222 21847 9274
rect 21899 9222 21911 9274
rect 21963 9222 21975 9274
rect 22027 9222 24840 9274
rect 1104 9200 24840 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 1360 9132 2697 9160
rect 1360 9120 1366 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 2685 9123 2743 9129
rect 3050 9120 3056 9172
rect 3108 9160 3114 9172
rect 3108 9132 3188 9160
rect 3108 9120 3114 9132
rect 1670 9052 1676 9104
rect 1728 9092 1734 9104
rect 2225 9095 2283 9101
rect 2225 9092 2237 9095
rect 1728 9064 2237 9092
rect 1728 9052 1734 9064
rect 2225 9061 2237 9064
rect 2271 9061 2283 9095
rect 2225 9055 2283 9061
rect 2590 9024 2596 9036
rect 1596 8996 2596 9024
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8956 1547 8959
rect 1596 8956 1624 8996
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 1535 8928 1624 8956
rect 1535 8925 1547 8928
rect 1489 8919 1547 8925
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2041 8959 2099 8965
rect 2041 8956 2053 8959
rect 1728 8928 2053 8956
rect 1728 8916 1734 8928
rect 2041 8925 2053 8928
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 3160 8965 3188 9132
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4065 9163 4123 9169
rect 4065 9160 4077 9163
rect 3844 9132 4077 9160
rect 3844 9120 3850 9132
rect 4065 9129 4077 9132
rect 4111 9129 4123 9163
rect 4065 9123 4123 9129
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 8481 9163 8539 9169
rect 7616 9132 8156 9160
rect 7616 9120 7622 9132
rect 3145 8959 3203 8965
rect 2280 8928 2774 8956
rect 2280 8916 2286 8928
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 1268 8860 2268 8888
rect 1268 8848 1274 8860
rect 658 8780 664 8832
rect 716 8820 722 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 716 8792 1593 8820
rect 716 8780 722 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 2240 8820 2268 8860
rect 2590 8848 2596 8900
rect 2648 8848 2654 8900
rect 2746 8888 2774 8928
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3602 8916 3608 8968
rect 3660 8956 3666 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 3660 8928 3985 8956
rect 3660 8916 3666 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 4249 8919 4307 8925
rect 7392 8928 7481 8956
rect 2746 8860 3832 8888
rect 3804 8829 3832 8860
rect 3237 8823 3295 8829
rect 3237 8820 3249 8823
rect 2240 8792 3249 8820
rect 1581 8783 1639 8789
rect 3237 8789 3249 8792
rect 3283 8789 3295 8823
rect 3237 8783 3295 8789
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8789 3847 8823
rect 4264 8820 4292 8919
rect 7392 8900 7420 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7743 8959 7801 8965
rect 7743 8956 7755 8959
rect 7469 8919 7527 8925
rect 7668 8928 7755 8956
rect 7668 8900 7696 8928
rect 7743 8925 7755 8928
rect 7789 8925 7801 8959
rect 7743 8919 7801 8925
rect 6362 8848 6368 8900
rect 6420 8888 6426 8900
rect 7282 8888 7288 8900
rect 6420 8860 7288 8888
rect 6420 8848 6426 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 7374 8848 7380 8900
rect 7432 8848 7438 8900
rect 7650 8848 7656 8900
rect 7708 8848 7714 8900
rect 8128 8888 8156 9132
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 8662 9160 8668 9172
rect 8527 9132 8668 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9088 9132 10548 9160
rect 9088 9120 9094 9132
rect 10520 9092 10548 9132
rect 10594 9120 10600 9172
rect 10652 9160 10658 9172
rect 10781 9163 10839 9169
rect 10781 9160 10793 9163
rect 10652 9132 10793 9160
rect 10652 9120 10658 9132
rect 10781 9129 10793 9132
rect 10827 9129 10839 9163
rect 10781 9123 10839 9129
rect 13464 9132 22416 9160
rect 13354 9092 13360 9104
rect 10520 9064 13360 9092
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 9769 9027 9827 9033
rect 9769 9024 9781 9027
rect 8956 8996 9781 9024
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8956 8956 8984 8996
rect 9769 8993 9781 8996
rect 9815 8993 9827 9027
rect 9769 8987 9827 8993
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 13464 9024 13492 9132
rect 13998 9052 14004 9104
rect 14056 9092 14062 9104
rect 22388 9092 22416 9132
rect 22462 9120 22468 9172
rect 22520 9160 22526 9172
rect 22649 9163 22707 9169
rect 22649 9160 22661 9163
rect 22520 9132 22661 9160
rect 22520 9120 22526 9132
rect 22649 9129 22661 9132
rect 22695 9129 22707 9163
rect 22649 9123 22707 9129
rect 23382 9120 23388 9172
rect 23440 9120 23446 9172
rect 23937 9163 23995 9169
rect 23937 9129 23949 9163
rect 23983 9160 23995 9163
rect 24026 9160 24032 9172
rect 23983 9132 24032 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 24026 9120 24032 9132
rect 24084 9120 24090 9172
rect 24118 9120 24124 9172
rect 24176 9120 24182 9172
rect 22738 9092 22744 9104
rect 14056 9064 14136 9092
rect 22388 9064 22744 9092
rect 14056 9052 14062 9064
rect 14108 9033 14136 9064
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 10560 8996 13492 9024
rect 14093 9027 14151 9033
rect 10560 8984 10566 8996
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14093 8987 14151 8993
rect 15470 8984 15476 9036
rect 15528 8984 15534 9036
rect 16298 9024 16304 9036
rect 16132 8996 16304 9024
rect 8536 8928 8984 8956
rect 8536 8916 8542 8928
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 10042 8956 10048 8968
rect 10003 8928 10048 8956
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 14335 8959 14393 8965
rect 14335 8956 14347 8959
rect 10152 8928 11652 8956
rect 9140 8888 9168 8916
rect 8128 8860 9168 8888
rect 9324 8888 9352 8916
rect 10152 8888 10180 8928
rect 9324 8860 10180 8888
rect 10226 8848 10232 8900
rect 10284 8888 10290 8900
rect 11514 8888 11520 8900
rect 10284 8860 11520 8888
rect 10284 8848 10290 8860
rect 11514 8848 11520 8860
rect 11572 8848 11578 8900
rect 11624 8888 11652 8928
rect 14108 8928 14347 8956
rect 14108 8888 14136 8928
rect 14335 8925 14347 8928
rect 14381 8925 14393 8959
rect 14335 8919 14393 8925
rect 15747 8959 15805 8965
rect 15747 8925 15759 8959
rect 15793 8956 15805 8959
rect 16132 8956 16160 8996
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16850 8984 16856 9036
rect 16908 8984 16914 9036
rect 15793 8928 16160 8956
rect 17095 8959 17153 8965
rect 15793 8925 15805 8928
rect 15747 8919 15805 8925
rect 17095 8925 17107 8959
rect 17141 8925 17153 8959
rect 17095 8919 17153 8925
rect 11624 8860 14136 8888
rect 14734 8820 14740 8832
rect 4264 8792 14740 8820
rect 3789 8783 3847 8789
rect 14734 8780 14740 8792
rect 14792 8780 14798 8832
rect 15102 8780 15108 8832
rect 15160 8780 15166 8832
rect 15470 8780 15476 8832
rect 15528 8820 15534 8832
rect 15762 8820 15790 8919
rect 17110 8888 17138 8919
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 17644 8928 18644 8956
rect 17644 8916 17650 8928
rect 18616 8900 18644 8928
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 22278 8956 22284 8968
rect 21324 8928 22284 8956
rect 21324 8916 21330 8928
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22370 8916 22376 8968
rect 22428 8916 22434 8968
rect 22925 8959 22983 8965
rect 22925 8925 22937 8959
rect 22971 8956 22983 8959
rect 23566 8956 23572 8968
rect 22971 8928 23572 8956
rect 22971 8925 22983 8928
rect 22925 8919 22983 8925
rect 23566 8916 23572 8928
rect 23624 8916 23630 8968
rect 23661 8959 23719 8965
rect 23661 8925 23673 8959
rect 23707 8956 23719 8959
rect 24136 8956 24164 9120
rect 23707 8928 24164 8956
rect 23707 8925 23719 8928
rect 23661 8919 23719 8925
rect 16132 8860 17138 8888
rect 16132 8832 16160 8860
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 21174 8888 21180 8900
rect 18656 8860 21180 8888
rect 18656 8848 18662 8860
rect 21174 8848 21180 8860
rect 21232 8848 21238 8900
rect 21536 8891 21594 8897
rect 21536 8857 21548 8891
rect 21582 8888 21594 8891
rect 22388 8888 22416 8916
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 21582 8860 22324 8888
rect 22388 8860 23121 8888
rect 21582 8857 21594 8860
rect 21536 8851 21594 8857
rect 15528 8792 15790 8820
rect 15528 8780 15534 8792
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 16482 8780 16488 8832
rect 16540 8780 16546 8832
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17184 8792 17877 8820
rect 17184 8780 17190 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 17865 8783 17923 8789
rect 18138 8780 18144 8832
rect 18196 8820 18202 8832
rect 20254 8820 20260 8832
rect 18196 8792 20260 8820
rect 18196 8780 18202 8792
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 22296 8820 22324 8860
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23109 8851 23167 8857
rect 22741 8823 22799 8829
rect 22741 8820 22753 8823
rect 22296 8792 22753 8820
rect 22741 8789 22753 8792
rect 22787 8820 22799 8823
rect 22830 8820 22836 8832
rect 22787 8792 22836 8820
rect 22787 8789 22799 8792
rect 22741 8783 22799 8789
rect 22830 8780 22836 8792
rect 22888 8780 22894 8832
rect 1104 8730 25000 8752
rect 1104 8678 6884 8730
rect 6936 8678 6948 8730
rect 7000 8678 7012 8730
rect 7064 8678 7076 8730
rect 7128 8678 7140 8730
rect 7192 8678 12818 8730
rect 12870 8678 12882 8730
rect 12934 8678 12946 8730
rect 12998 8678 13010 8730
rect 13062 8678 13074 8730
rect 13126 8678 18752 8730
rect 18804 8678 18816 8730
rect 18868 8678 18880 8730
rect 18932 8678 18944 8730
rect 18996 8678 19008 8730
rect 19060 8678 24686 8730
rect 24738 8678 24750 8730
rect 24802 8678 24814 8730
rect 24866 8678 24878 8730
rect 24930 8678 24942 8730
rect 24994 8678 25000 8730
rect 1104 8656 25000 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1452 8588 1593 8616
rect 1452 8576 1458 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 1581 8579 1639 8585
rect 2746 8588 7113 8616
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 1946 8548 1952 8560
rect 1535 8520 1952 8548
rect 1535 8517 1547 8520
rect 1489 8511 1547 8517
rect 1946 8508 1952 8520
rect 2004 8508 2010 8560
rect 2593 8551 2651 8557
rect 2593 8517 2605 8551
rect 2639 8548 2651 8551
rect 2746 8548 2774 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8389 8619 8447 8625
rect 8389 8616 8401 8619
rect 8168 8588 8401 8616
rect 8168 8576 8174 8588
rect 8389 8585 8401 8588
rect 8435 8585 8447 8619
rect 8389 8579 8447 8585
rect 10137 8619 10195 8625
rect 10137 8585 10149 8619
rect 10183 8616 10195 8619
rect 10318 8616 10324 8628
rect 10183 8588 10324 8616
rect 10183 8585 10195 8588
rect 10137 8579 10195 8585
rect 10318 8576 10324 8588
rect 10376 8576 10382 8628
rect 12989 8619 13047 8625
rect 10428 8588 12940 8616
rect 2639 8520 2774 8548
rect 2639 8517 2651 8520
rect 2593 8511 2651 8517
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 7742 8548 7748 8560
rect 6052 8520 7748 8548
rect 6052 8508 6058 8520
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 2038 8440 2044 8492
rect 2096 8440 2102 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8480 2467 8483
rect 2866 8480 2872 8492
rect 2455 8452 2872 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 7651 8483 7709 8489
rect 7651 8480 7663 8483
rect 7616 8452 7663 8480
rect 7616 8440 7622 8452
rect 7651 8449 7663 8452
rect 7697 8449 7709 8483
rect 9367 8483 9425 8489
rect 9367 8480 9379 8483
rect 7651 8443 7709 8449
rect 8496 8452 9379 8480
rect 842 8372 848 8424
rect 900 8412 906 8424
rect 900 8384 3924 8412
rect 900 8372 906 8384
rect 1026 8304 1032 8356
rect 1084 8344 1090 8356
rect 2777 8347 2835 8353
rect 2777 8344 2789 8347
rect 1084 8316 2789 8344
rect 1084 8304 1090 8316
rect 2777 8313 2789 8316
rect 2823 8313 2835 8347
rect 2777 8307 2835 8313
rect 3326 8304 3332 8356
rect 3384 8304 3390 8356
rect 3896 8353 3924 8384
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7374 8412 7380 8424
rect 6788 8384 7380 8412
rect 6788 8372 6794 8384
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 8496 8356 8524 8452
rect 9367 8449 9379 8452
rect 9413 8480 9425 8483
rect 10428 8480 10456 8588
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11701 8551 11759 8557
rect 11701 8548 11713 8551
rect 11664 8520 11713 8548
rect 11664 8508 11670 8520
rect 11701 8517 11713 8520
rect 11747 8517 11759 8551
rect 11701 8511 11759 8517
rect 11974 8508 11980 8560
rect 12032 8508 12038 8560
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 12308 8520 12449 8548
rect 12308 8508 12314 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 12805 8551 12863 8557
rect 12805 8517 12817 8551
rect 12851 8517 12863 8551
rect 12805 8511 12863 8517
rect 9413 8452 10456 8480
rect 9413 8449 9425 8452
rect 9367 8443 9425 8449
rect 12066 8440 12072 8492
rect 12124 8440 12130 8492
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12820 8480 12848 8511
rect 12676 8452 12848 8480
rect 12912 8480 12940 8588
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13354 8616 13360 8628
rect 13035 8588 13360 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 16666 8576 16672 8628
rect 16724 8616 16730 8628
rect 17129 8619 17187 8625
rect 17129 8616 17141 8619
rect 16724 8588 17141 8616
rect 16724 8576 16730 8588
rect 17129 8585 17141 8588
rect 17175 8585 17187 8619
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 17129 8579 17187 8585
rect 17512 8588 19625 8616
rect 13170 8508 13176 8560
rect 13228 8548 13234 8560
rect 13630 8548 13636 8560
rect 13228 8520 13636 8548
rect 13228 8508 13234 8520
rect 13630 8508 13636 8520
rect 13688 8548 13694 8560
rect 13817 8551 13875 8557
rect 13817 8548 13829 8551
rect 13688 8520 13829 8548
rect 13688 8508 13694 8520
rect 13817 8517 13829 8520
rect 13863 8517 13875 8551
rect 13817 8511 13875 8517
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8548 14243 8551
rect 14231 8520 14688 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 13538 8480 13544 8492
rect 12912 8452 13544 8480
rect 12676 8440 12682 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 14056 8452 14105 8480
rect 14056 8440 14062 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14274 8440 14280 8492
rect 14332 8480 14338 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14332 8452 14565 8480
rect 14332 8440 14338 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14660 8480 14688 8520
rect 14918 8508 14924 8560
rect 14976 8508 14982 8560
rect 15102 8508 15108 8560
rect 15160 8508 15166 8560
rect 17310 8508 17316 8560
rect 17368 8548 17374 8560
rect 17512 8557 17540 8588
rect 19613 8585 19625 8588
rect 19659 8585 19671 8619
rect 19613 8579 19671 8585
rect 22186 8576 22192 8628
rect 22244 8576 22250 8628
rect 23290 8616 23296 8628
rect 22480 8588 23296 8616
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 17368 8520 17417 8548
rect 17368 8508 17374 8520
rect 17405 8517 17417 8520
rect 17451 8517 17463 8551
rect 17405 8511 17463 8517
rect 17497 8551 17555 8557
rect 17497 8517 17509 8551
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 22204 8548 22232 8576
rect 22480 8560 22508 8588
rect 23290 8576 23296 8588
rect 23348 8576 23354 8628
rect 23750 8576 23756 8628
rect 23808 8576 23814 8628
rect 18196 8520 19472 8548
rect 22204 8520 22324 8548
rect 18196 8508 18202 8520
rect 15120 8480 15148 8508
rect 14660 8452 15148 8480
rect 14553 8443 14611 8449
rect 17862 8440 17868 8492
rect 17920 8440 17926 8492
rect 18247 8483 18305 8489
rect 18247 8449 18259 8483
rect 18293 8480 18305 8483
rect 18293 8452 18368 8480
rect 18293 8449 18305 8452
rect 18247 8443 18305 8449
rect 11520 8424 11572 8430
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 9125 8415 9183 8421
rect 9125 8412 9137 8415
rect 8628 8384 9137 8412
rect 8628 8372 8634 8384
rect 9125 8381 9137 8384
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 11520 8366 11572 8372
rect 13820 8424 13872 8430
rect 15562 8412 15568 8424
rect 13820 8366 13872 8372
rect 15120 8384 15568 8412
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8313 3939 8347
rect 3881 8307 3939 8313
rect 8478 8304 8484 8356
rect 8536 8304 8542 8356
rect 10042 8304 10048 8356
rect 10100 8344 10106 8356
rect 10502 8344 10508 8356
rect 10100 8316 10508 8344
rect 10100 8304 10106 8316
rect 10502 8304 10508 8316
rect 10560 8344 10566 8356
rect 10870 8344 10876 8356
rect 10560 8316 10876 8344
rect 10560 8304 10566 8316
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 15120 8353 15148 8384
rect 15562 8372 15568 8384
rect 15620 8372 15626 8424
rect 17678 8372 17684 8424
rect 17736 8372 17742 8424
rect 15105 8347 15163 8353
rect 15105 8313 15117 8347
rect 15151 8313 15163 8347
rect 18340 8344 18368 8452
rect 18598 8440 18604 8492
rect 18656 8440 18662 8492
rect 18782 8440 18788 8492
rect 18840 8480 18846 8492
rect 18875 8483 18933 8489
rect 18875 8480 18887 8483
rect 18840 8452 18887 8480
rect 18840 8440 18846 8452
rect 18875 8449 18887 8452
rect 18921 8480 18933 8483
rect 19334 8480 19340 8492
rect 18921 8452 19340 8480
rect 18921 8449 18933 8452
rect 18875 8443 18933 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19444 8344 19472 8520
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19576 8452 19993 8480
rect 19576 8440 19582 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20162 8440 20168 8492
rect 20220 8440 20226 8492
rect 21542 8440 21548 8492
rect 21600 8480 21606 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21600 8452 21833 8480
rect 21600 8440 21606 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22189 8483 22247 8489
rect 22189 8480 22201 8483
rect 22152 8452 22201 8480
rect 22152 8440 22158 8452
rect 22189 8449 22201 8452
rect 22235 8449 22247 8483
rect 22296 8480 22324 8520
rect 22462 8508 22468 8560
rect 22520 8508 22526 8560
rect 22738 8508 22744 8560
rect 22796 8548 22802 8560
rect 22925 8551 22983 8557
rect 22925 8548 22937 8551
rect 22796 8520 22937 8548
rect 22796 8508 22802 8520
rect 22925 8517 22937 8520
rect 22971 8517 22983 8551
rect 23768 8548 23796 8576
rect 23768 8520 24532 8548
rect 22925 8511 22983 8517
rect 22649 8483 22707 8489
rect 22649 8480 22661 8483
rect 22296 8452 22661 8480
rect 22189 8443 22247 8449
rect 22649 8449 22661 8452
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 23014 8440 23020 8492
rect 23072 8480 23078 8492
rect 23477 8483 23535 8489
rect 23477 8480 23489 8483
rect 23072 8452 23489 8480
rect 23072 8440 23078 8452
rect 23477 8449 23489 8452
rect 23523 8449 23535 8483
rect 23477 8443 23535 8449
rect 24026 8440 24032 8492
rect 24084 8440 24090 8492
rect 24504 8489 24532 8520
rect 24489 8483 24547 8489
rect 24489 8449 24501 8483
rect 24535 8449 24547 8483
rect 24489 8443 24547 8449
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 22462 8412 22468 8424
rect 20680 8384 22468 8412
rect 20680 8372 20686 8384
rect 22462 8372 22468 8384
rect 22520 8372 22526 8424
rect 23293 8415 23351 8421
rect 22572 8384 22784 8412
rect 22572 8344 22600 8384
rect 18340 8316 18736 8344
rect 19444 8316 22600 8344
rect 22756 8344 22784 8384
rect 23293 8381 23305 8415
rect 23339 8412 23351 8415
rect 23566 8412 23572 8424
rect 23339 8384 23572 8412
rect 23339 8381 23351 8384
rect 23293 8375 23351 8381
rect 23566 8372 23572 8384
rect 23624 8372 23630 8424
rect 23937 8347 23995 8353
rect 23937 8344 23949 8347
rect 22756 8316 23949 8344
rect 15105 8307 15163 8313
rect 18708 8288 18736 8316
rect 23937 8313 23949 8316
rect 23983 8313 23995 8347
rect 23937 8307 23995 8313
rect 24228 8316 24440 8344
rect 474 8236 480 8288
rect 532 8276 538 8288
rect 2406 8276 2412 8288
rect 532 8248 2412 8276
rect 532 8236 538 8248
rect 2406 8236 2412 8248
rect 2464 8236 2470 8288
rect 2682 8236 2688 8288
rect 2740 8276 2746 8288
rect 11698 8276 11704 8288
rect 2740 8248 11704 8276
rect 2740 8236 2746 8248
rect 11698 8236 11704 8248
rect 11756 8236 11762 8288
rect 18417 8279 18475 8285
rect 18417 8245 18429 8279
rect 18463 8276 18475 8279
rect 18598 8276 18604 8288
rect 18463 8248 18604 8276
rect 18463 8245 18475 8248
rect 18417 8239 18475 8245
rect 18598 8236 18604 8248
rect 18656 8236 18662 8288
rect 18690 8236 18696 8288
rect 18748 8236 18754 8288
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20073 8279 20131 8285
rect 20073 8276 20085 8279
rect 20036 8248 20085 8276
rect 20036 8236 20042 8248
rect 20073 8245 20085 8248
rect 20119 8245 20131 8279
rect 20073 8239 20131 8245
rect 22738 8236 22744 8288
rect 22796 8276 22802 8288
rect 24228 8276 24256 8316
rect 22796 8248 24256 8276
rect 22796 8236 22802 8248
rect 24302 8236 24308 8288
rect 24360 8236 24366 8288
rect 24412 8276 24440 8316
rect 24670 8276 24676 8288
rect 24412 8248 24676 8276
rect 24670 8236 24676 8248
rect 24728 8236 24734 8288
rect 1104 8186 24840 8208
rect 1104 8134 3917 8186
rect 3969 8134 3981 8186
rect 4033 8134 4045 8186
rect 4097 8134 4109 8186
rect 4161 8134 4173 8186
rect 4225 8134 9851 8186
rect 9903 8134 9915 8186
rect 9967 8134 9979 8186
rect 10031 8134 10043 8186
rect 10095 8134 10107 8186
rect 10159 8134 15785 8186
rect 15837 8134 15849 8186
rect 15901 8134 15913 8186
rect 15965 8134 15977 8186
rect 16029 8134 16041 8186
rect 16093 8134 21719 8186
rect 21771 8134 21783 8186
rect 21835 8134 21847 8186
rect 21899 8134 21911 8186
rect 21963 8134 21975 8186
rect 22027 8134 24840 8186
rect 1104 8112 24840 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 1854 8072 1860 8084
rect 1811 8044 1860 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 2096 8044 3341 8072
rect 2096 8032 2102 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 5350 8072 5356 8084
rect 3329 8035 3387 8041
rect 4908 8044 5356 8072
rect 4706 8004 4712 8016
rect 2746 7976 4712 8004
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 1504 7732 1532 7831
rect 1964 7800 1992 7831
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2223 7871 2281 7877
rect 2223 7868 2235 7871
rect 2188 7840 2235 7868
rect 2188 7828 2194 7840
rect 2223 7837 2235 7840
rect 2269 7837 2281 7871
rect 2746 7868 2774 7976
rect 4706 7964 4712 7976
rect 4764 7964 4770 8016
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 3844 7908 4292 7936
rect 3844 7896 3850 7908
rect 2223 7831 2281 7837
rect 2332 7840 2774 7868
rect 3513 7871 3571 7877
rect 2038 7800 2044 7812
rect 1964 7772 2044 7800
rect 2038 7760 2044 7772
rect 2096 7800 2102 7812
rect 2332 7800 2360 7840
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 3973 7871 4031 7877
rect 3559 7840 3924 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 2096 7772 2360 7800
rect 2096 7760 2102 7772
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 3896 7800 3924 7840
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4154 7868 4160 7880
rect 4019 7840 4160 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 4264 7877 4292 7908
rect 4430 7896 4436 7948
rect 4488 7936 4494 7948
rect 4908 7936 4936 8044
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 7190 8072 7196 8084
rect 7024 8044 7196 8072
rect 5905 8007 5963 8013
rect 5905 7973 5917 8007
rect 5951 8004 5963 8007
rect 6917 8007 6975 8013
rect 6917 8004 6929 8007
rect 5951 7976 6929 8004
rect 5951 7973 5963 7976
rect 5905 7967 5963 7973
rect 6917 7973 6929 7976
rect 6963 7973 6975 8007
rect 6917 7967 6975 7973
rect 4488 7908 4936 7936
rect 4488 7896 4494 7908
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 6457 7939 6515 7945
rect 6457 7905 6469 7939
rect 6503 7936 6515 7939
rect 6546 7936 6552 7948
rect 6503 7908 6552 7936
rect 6503 7905 6515 7908
rect 6457 7899 6515 7905
rect 6546 7896 6552 7908
rect 6604 7896 6610 7948
rect 7024 7936 7052 8044
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7340 8044 8125 8072
rect 7340 8032 7346 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 10873 8075 10931 8081
rect 8113 8035 8171 8041
rect 9876 8044 10824 8072
rect 7374 7945 7380 7948
rect 7193 7939 7251 7945
rect 7193 7936 7205 7939
rect 7024 7908 7205 7936
rect 7193 7905 7205 7908
rect 7239 7905 7251 7939
rect 7193 7899 7251 7905
rect 7331 7939 7380 7945
rect 7331 7905 7343 7939
rect 7377 7905 7380 7939
rect 7331 7899 7380 7905
rect 7374 7896 7380 7899
rect 7432 7936 7438 7948
rect 9876 7945 9904 8044
rect 10796 7948 10824 8044
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11514 8072 11520 8084
rect 10919 8044 11520 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 12124 8044 12265 8072
rect 12124 8032 12130 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12618 8072 12624 8084
rect 12492 8044 12624 8072
rect 12492 8032 12498 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13814 8072 13820 8084
rect 13679 8044 13820 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 16482 8072 16488 8084
rect 15948 8044 16488 8072
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 15838 8004 15844 8016
rect 15436 7976 15844 8004
rect 15436 7964 15442 7976
rect 9861 7939 9919 7945
rect 7432 7908 9101 7936
rect 7432 7896 7438 7908
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 5167 7871 5225 7877
rect 5167 7837 5179 7871
rect 5213 7868 5225 7871
rect 6362 7868 6368 7880
rect 5213 7840 6368 7868
rect 5213 7837 5225 7840
rect 5167 7831 5225 7837
rect 6362 7828 6368 7840
rect 6420 7828 6426 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 5902 7800 5908 7812
rect 2464 7772 2636 7800
rect 2464 7760 2470 7772
rect 2498 7732 2504 7744
rect 1504 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2608 7732 2636 7772
rect 2746 7772 3832 7800
rect 3896 7772 5908 7800
rect 2746 7732 2774 7772
rect 2608 7704 2774 7732
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 3804 7741 3832 7772
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 3789 7735 3847 7741
rect 3789 7701 3801 7735
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3936 7704 4077 7732
rect 3936 7692 3942 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 6380 7732 6408 7828
rect 9073 7800 9101 7908
rect 9861 7905 9873 7939
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10778 7896 10784 7948
rect 10836 7936 10842 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 10836 7908 11253 7936
rect 10836 7896 10842 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 11241 7899 11299 7905
rect 12158 7896 12164 7948
rect 12216 7936 12222 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12216 7908 12633 7936
rect 12216 7896 12222 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 13354 7896 13360 7948
rect 13412 7936 13418 7948
rect 15488 7945 15516 7976
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 15948 8013 15976 8044
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16908 8044 17908 8072
rect 16908 8032 16914 8044
rect 15933 8007 15991 8013
rect 15933 7973 15945 8007
rect 15979 7973 15991 8007
rect 15933 7967 15991 7973
rect 15473 7939 15531 7945
rect 15473 7936 15485 7939
rect 13412 7908 15485 7936
rect 13412 7896 13418 7908
rect 15473 7905 15485 7908
rect 15519 7905 15531 7939
rect 15473 7899 15531 7905
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 16326 7939 16384 7945
rect 16326 7936 16338 7939
rect 15620 7908 16338 7936
rect 15620 7896 15626 7908
rect 16326 7905 16338 7908
rect 16372 7905 16384 7939
rect 16326 7899 16384 7905
rect 16485 7939 16543 7945
rect 16485 7905 16497 7939
rect 16531 7936 16543 7939
rect 17126 7936 17132 7948
rect 16531 7908 17132 7936
rect 16531 7905 16543 7908
rect 16485 7899 16543 7905
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 17880 7936 17908 8044
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18690 8072 18696 8084
rect 18472 8044 18696 8072
rect 18472 8032 18478 8044
rect 18690 8032 18696 8044
rect 18748 8072 18754 8084
rect 19889 8075 19947 8081
rect 18748 8044 19564 8072
rect 18748 8032 18754 8044
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 18598 8004 18604 8016
rect 18012 7976 18604 8004
rect 18012 7964 18018 7976
rect 18598 7964 18604 7976
rect 18656 7964 18662 8016
rect 19429 8007 19487 8013
rect 19429 8004 19441 8007
rect 18708 7976 19441 8004
rect 18708 7936 18736 7976
rect 19429 7973 19441 7976
rect 19475 7973 19487 8007
rect 19429 7967 19487 7973
rect 17880 7908 18736 7936
rect 18877 7939 18935 7945
rect 18877 7905 18889 7939
rect 18923 7936 18935 7939
rect 19536 7936 19564 8044
rect 19889 8041 19901 8075
rect 19935 8072 19947 8075
rect 20162 8072 20168 8084
rect 19935 8044 20168 8072
rect 19935 8041 19947 8044
rect 19889 8035 19947 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 22462 8072 22468 8084
rect 21048 8044 22468 8072
rect 21048 8032 21054 8044
rect 22462 8032 22468 8044
rect 22520 8032 22526 8084
rect 22649 8075 22707 8081
rect 22649 8041 22661 8075
rect 22695 8072 22707 8075
rect 23014 8072 23020 8084
rect 22695 8044 23020 8072
rect 22695 8041 22707 8044
rect 22649 8035 22707 8041
rect 23014 8032 23020 8044
rect 23072 8032 23078 8084
rect 20070 7964 20076 8016
rect 20128 8004 20134 8016
rect 22738 8004 22744 8016
rect 20128 7976 22744 8004
rect 20128 7964 20134 7976
rect 22738 7964 22744 7976
rect 22796 7964 22802 8016
rect 21177 7939 21235 7945
rect 21177 7936 21189 7939
rect 18923 7908 19472 7936
rect 19536 7908 21189 7936
rect 18923 7905 18935 7908
rect 18877 7899 18935 7905
rect 10135 7871 10193 7877
rect 10135 7837 10147 7871
rect 10181 7868 10193 7871
rect 11515 7871 11573 7877
rect 10181 7840 11192 7868
rect 10181 7837 10193 7840
rect 10135 7831 10193 7837
rect 10962 7800 10968 7812
rect 9073 7772 10968 7800
rect 10962 7760 10968 7772
rect 11020 7760 11026 7812
rect 11164 7800 11192 7840
rect 11515 7837 11527 7871
rect 11561 7868 11573 7871
rect 11882 7868 11888 7880
rect 11561 7840 11888 7868
rect 11561 7837 11573 7840
rect 11515 7831 11573 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 12879 7841 12937 7847
rect 11422 7800 11428 7812
rect 11164 7772 11428 7800
rect 11422 7760 11428 7772
rect 11480 7760 11486 7812
rect 12879 7807 12891 7841
rect 12925 7838 12937 7841
rect 12925 7807 12940 7838
rect 14734 7828 14740 7880
rect 14792 7828 14798 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15378 7868 15384 7880
rect 15335 7840 15384 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15378 7828 15384 7840
rect 15436 7828 15442 7880
rect 16206 7828 16212 7880
rect 16264 7828 16270 7880
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7837 17279 7871
rect 17221 7831 17279 7837
rect 12879 7801 12940 7807
rect 12912 7732 12940 7801
rect 6380 7704 12940 7732
rect 14752 7732 14780 7828
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 14752 7704 17141 7732
rect 4065 7695 4123 7701
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 17236 7732 17264 7831
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17495 7871 17553 7877
rect 17495 7868 17507 7871
rect 17460 7840 17507 7868
rect 17460 7828 17466 7840
rect 17495 7837 17507 7840
rect 17541 7868 17553 7871
rect 17541 7840 18552 7868
rect 17541 7837 17553 7840
rect 17495 7831 17553 7837
rect 17310 7760 17316 7812
rect 17368 7800 17374 7812
rect 18524 7800 18552 7840
rect 18598 7828 18604 7880
rect 18656 7868 18662 7880
rect 19444 7877 19472 7908
rect 21177 7905 21189 7908
rect 21223 7905 21235 7939
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 21177 7899 21235 7905
rect 22388 7908 22845 7936
rect 22388 7880 22416 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 22833 7899 22891 7905
rect 18785 7871 18843 7877
rect 18785 7868 18797 7871
rect 18656 7840 18797 7868
rect 18656 7828 18662 7840
rect 18785 7837 18797 7840
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19576 7840 19625 7868
rect 19576 7828 19582 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19944 7840 20085 7868
rect 19944 7828 19950 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20346 7828 20352 7880
rect 20404 7828 20410 7880
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 21082 7828 21088 7880
rect 21140 7828 21146 7880
rect 22370 7828 22376 7880
rect 22428 7828 22434 7880
rect 22465 7871 22523 7877
rect 22465 7837 22477 7871
rect 22511 7837 22523 7871
rect 22465 7831 22523 7837
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7868 22615 7871
rect 23658 7868 23664 7880
rect 22603 7840 23664 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 19334 7800 19340 7812
rect 17368 7772 18368 7800
rect 18524 7772 19340 7800
rect 17368 7760 17374 7772
rect 17586 7732 17592 7744
rect 17236 7704 17592 7732
rect 17129 7695 17187 7701
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 17678 7692 17684 7744
rect 17736 7732 17742 7744
rect 18233 7735 18291 7741
rect 18233 7732 18245 7735
rect 17736 7704 18245 7732
rect 17736 7692 17742 7704
rect 18233 7701 18245 7704
rect 18279 7701 18291 7735
rect 18340 7732 18368 7772
rect 19334 7760 19340 7772
rect 19392 7760 19398 7812
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 19978 7800 19984 7812
rect 19843 7772 19984 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 22480 7800 22508 7831
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 23100 7803 23158 7809
rect 22480 7772 22784 7800
rect 20806 7732 20812 7744
rect 18340 7704 20812 7732
rect 18233 7695 18291 7701
rect 20806 7692 20812 7704
rect 20864 7692 20870 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 22756 7732 22784 7772
rect 23100 7769 23112 7803
rect 23146 7800 23158 7803
rect 23934 7800 23940 7812
rect 23146 7772 23940 7800
rect 23146 7769 23158 7772
rect 23100 7763 23158 7769
rect 23934 7760 23940 7772
rect 23992 7760 23998 7812
rect 24213 7735 24271 7741
rect 24213 7732 24225 7735
rect 22756 7704 24225 7732
rect 24213 7701 24225 7704
rect 24259 7701 24271 7735
rect 24213 7695 24271 7701
rect 1104 7642 25000 7664
rect 1104 7590 6884 7642
rect 6936 7590 6948 7642
rect 7000 7590 7012 7642
rect 7064 7590 7076 7642
rect 7128 7590 7140 7642
rect 7192 7590 12818 7642
rect 12870 7590 12882 7642
rect 12934 7590 12946 7642
rect 12998 7590 13010 7642
rect 13062 7590 13074 7642
rect 13126 7590 18752 7642
rect 18804 7590 18816 7642
rect 18868 7590 18880 7642
rect 18932 7590 18944 7642
rect 18996 7590 19008 7642
rect 19060 7590 24686 7642
rect 24738 7590 24750 7642
rect 24802 7590 24814 7642
rect 24866 7590 24878 7642
rect 24930 7590 24942 7642
rect 24994 7590 25000 7642
rect 1104 7568 25000 7590
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2590 7528 2596 7540
rect 2179 7500 2596 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4249 7531 4307 7537
rect 4249 7528 4261 7531
rect 4212 7500 4261 7528
rect 4212 7488 4218 7500
rect 4249 7497 4261 7500
rect 4295 7497 4307 7531
rect 4249 7491 4307 7497
rect 4890 7488 4896 7540
rect 4948 7528 4954 7540
rect 5810 7528 5816 7540
rect 4948 7500 5816 7528
rect 4948 7488 4954 7500
rect 5810 7488 5816 7500
rect 5868 7528 5874 7540
rect 6730 7528 6736 7540
rect 5868 7500 6736 7528
rect 5868 7488 5874 7500
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2363 7364 2820 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 382 7284 388 7336
rect 440 7324 446 7336
rect 1854 7324 1860 7336
rect 440 7296 1860 7324
rect 440 7284 446 7296
rect 1854 7284 1860 7296
rect 1912 7324 1918 7336
rect 2409 7327 2467 7333
rect 2409 7324 2421 7327
rect 1912 7296 2421 7324
rect 1912 7284 1918 7296
rect 2409 7293 2421 7296
rect 2455 7293 2467 7327
rect 2409 7287 2467 7293
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 2682 7324 2688 7336
rect 2639 7296 2688 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 2792 7188 2820 7364
rect 3418 7352 3424 7404
rect 3476 7401 3482 7404
rect 3476 7395 3504 7401
rect 3492 7361 3504 7395
rect 3476 7355 3504 7361
rect 3476 7352 3482 7355
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 6472 7401 6500 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7466 7488 7472 7540
rect 7524 7488 7530 7540
rect 9306 7528 9312 7540
rect 8220 7500 9312 7528
rect 8220 7460 8248 7500
rect 9306 7488 9312 7500
rect 9364 7488 9370 7540
rect 9674 7488 9680 7540
rect 9732 7488 9738 7540
rect 9766 7488 9772 7540
rect 9824 7528 9830 7540
rect 13354 7528 13360 7540
rect 9824 7500 13360 7528
rect 9824 7488 9830 7500
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 13998 7528 14004 7540
rect 13556 7500 14004 7528
rect 9490 7460 9496 7472
rect 6748 7432 8248 7460
rect 9416 7432 9496 7460
rect 6748 7431 6776 7432
rect 6715 7425 6776 7431
rect 6457 7395 6515 7401
rect 6457 7361 6469 7395
rect 6503 7361 6515 7395
rect 6715 7391 6727 7425
rect 6761 7394 6776 7425
rect 8279 7425 8337 7431
rect 6761 7391 6773 7394
rect 6715 7385 6773 7391
rect 8279 7391 8291 7425
rect 8325 7422 8337 7425
rect 8325 7392 8340 7422
rect 8662 7392 8668 7404
rect 8325 7391 8668 7392
rect 8279 7385 8668 7391
rect 8312 7364 8668 7385
rect 6457 7355 6515 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3053 7327 3111 7333
rect 3053 7324 3065 7327
rect 3016 7296 3065 7324
rect 3016 7284 3022 7296
rect 3053 7293 3065 7296
rect 3099 7293 3111 7327
rect 3053 7287 3111 7293
rect 3329 7327 3387 7333
rect 3329 7293 3341 7327
rect 3375 7324 3387 7327
rect 4341 7327 4399 7333
rect 3375 7296 4200 7324
rect 3375 7293 3387 7296
rect 3329 7287 3387 7293
rect 4172 7256 4200 7296
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4430 7324 4436 7336
rect 4387 7296 4436 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 4522 7284 4528 7336
rect 4580 7284 4586 7336
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5074 7324 5080 7336
rect 4672 7296 5080 7324
rect 4672 7284 4678 7296
rect 5074 7284 5080 7296
rect 5132 7324 5138 7336
rect 5378 7327 5436 7333
rect 5378 7324 5390 7327
rect 5132 7296 5390 7324
rect 5132 7284 5138 7296
rect 5378 7293 5390 7296
rect 5424 7293 5436 7327
rect 5378 7287 5436 7293
rect 5534 7284 5540 7336
rect 5592 7284 5598 7336
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7293 8079 7327
rect 9214 7324 9220 7336
rect 8021 7287 8079 7293
rect 8680 7296 9220 7324
rect 4632 7256 4660 7284
rect 4172 7228 4660 7256
rect 4982 7216 4988 7268
rect 5040 7216 5046 7268
rect 6181 7259 6239 7265
rect 6181 7225 6193 7259
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 6196 7188 6224 7219
rect 2792 7160 6224 7188
rect 6362 7148 6368 7200
rect 6420 7188 6426 7200
rect 8036 7188 8064 7287
rect 8680 7188 8708 7296
rect 9214 7284 9220 7296
rect 9272 7324 9278 7336
rect 9416 7333 9444 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 9692 7411 9720 7488
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 13556 7469 13584 7500
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7497 14427 7531
rect 14369 7491 14427 7497
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 16666 7528 16672 7540
rect 14599 7500 16672 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 13265 7463 13323 7469
rect 13265 7460 13277 7463
rect 13228 7432 13277 7460
rect 13228 7420 13234 7432
rect 13265 7429 13277 7432
rect 13311 7429 13323 7463
rect 13265 7423 13323 7429
rect 13541 7463 13599 7469
rect 13541 7429 13553 7463
rect 13587 7429 13599 7463
rect 13541 7423 13599 7429
rect 14384 7460 14412 7491
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 18414 7528 18420 7540
rect 16776 7500 18420 7528
rect 14918 7460 14924 7472
rect 14384 7432 14924 7460
rect 9675 7405 9733 7411
rect 9675 7371 9687 7405
rect 9721 7371 9733 7405
rect 14384 7404 14412 7432
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 15838 7420 15844 7472
rect 15896 7460 15902 7472
rect 16776 7460 16804 7500
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 19521 7531 19579 7537
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 19886 7528 19892 7540
rect 19567 7500 19892 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 19981 7531 20039 7537
rect 19981 7497 19993 7531
rect 20027 7528 20039 7531
rect 20622 7528 20628 7540
rect 20027 7500 20628 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 21545 7531 21603 7537
rect 21545 7497 21557 7531
rect 21591 7497 21603 7531
rect 21545 7491 21603 7497
rect 23293 7531 23351 7537
rect 23293 7497 23305 7531
rect 23339 7528 23351 7531
rect 23566 7528 23572 7540
rect 23339 7500 23572 7528
rect 23339 7497 23351 7500
rect 23293 7491 23351 7497
rect 15896 7432 16804 7460
rect 15896 7420 15902 7432
rect 16942 7420 16948 7472
rect 17000 7460 17006 7472
rect 17310 7460 17316 7472
rect 17000 7432 17316 7460
rect 17000 7420 17006 7432
rect 17310 7420 17316 7432
rect 17368 7420 17374 7472
rect 19702 7460 19708 7472
rect 18156 7432 19708 7460
rect 9675 7365 9733 7371
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13906 7392 13912 7404
rect 13679 7364 13912 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13906 7352 13912 7364
rect 13964 7352 13970 7404
rect 14001 7395 14059 7401
rect 14001 7361 14013 7395
rect 14047 7392 14059 7395
rect 14182 7392 14188 7404
rect 14047 7364 14188 7392
rect 14047 7361 14059 7364
rect 14001 7355 14059 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 18156 7401 18184 7432
rect 19702 7420 19708 7432
rect 19760 7460 19766 7472
rect 19760 7432 20208 7460
rect 19760 7420 19766 7432
rect 18141 7395 18199 7401
rect 18141 7361 18153 7395
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18408 7395 18466 7401
rect 18408 7361 18420 7395
rect 18454 7392 18466 7395
rect 18782 7392 18788 7404
rect 18454 7364 18788 7392
rect 18454 7361 18466 7364
rect 18408 7355 18466 7361
rect 18782 7352 18788 7364
rect 18840 7352 18846 7404
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 9401 7327 9459 7333
rect 9401 7324 9413 7327
rect 9272 7296 9413 7324
rect 9272 7284 9278 7296
rect 9401 7293 9413 7296
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 13446 7284 13452 7336
rect 13504 7284 13510 7336
rect 6420 7160 8708 7188
rect 6420 7148 6426 7160
rect 9030 7148 9036 7200
rect 9088 7148 9094 7200
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9766 7188 9772 7200
rect 9548 7160 9772 7188
rect 9548 7148 9554 7160
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 10376 7160 10425 7188
rect 10376 7148 10382 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 19904 7188 19932 7355
rect 20180 7336 20208 7432
rect 20432 7395 20490 7401
rect 20432 7361 20444 7395
rect 20478 7392 20490 7395
rect 20898 7392 20904 7404
rect 20478 7364 20904 7392
rect 20478 7361 20490 7364
rect 20432 7355 20490 7361
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 21560 7392 21588 7491
rect 23566 7488 23572 7500
rect 23624 7488 23630 7540
rect 23658 7488 23664 7540
rect 23716 7488 23722 7540
rect 23934 7488 23940 7540
rect 23992 7528 23998 7540
rect 23992 7500 24532 7528
rect 23992 7488 23998 7500
rect 22554 7431 22560 7472
rect 22539 7425 22560 7431
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21560 7364 22017 7392
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22539 7391 22551 7425
rect 22612 7420 22618 7472
rect 22585 7394 22600 7420
rect 22585 7391 22597 7394
rect 22539 7385 22597 7391
rect 22005 7355 22063 7361
rect 20162 7284 20168 7336
rect 20220 7284 20226 7336
rect 21542 7284 21548 7336
rect 21600 7324 21606 7336
rect 22094 7324 22100 7336
rect 21600 7296 22100 7324
rect 21600 7284 21606 7296
rect 22094 7284 22100 7296
rect 22152 7324 22158 7336
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22152 7296 22293 7324
rect 22152 7284 22158 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22281 7287 22339 7293
rect 23676 7256 23704 7488
rect 23845 7463 23903 7469
rect 23845 7429 23857 7463
rect 23891 7460 23903 7463
rect 24302 7460 24308 7472
rect 23891 7432 24308 7460
rect 23891 7429 23903 7432
rect 23845 7423 23903 7429
rect 24302 7420 24308 7432
rect 24360 7420 24366 7472
rect 24394 7352 24400 7404
rect 24452 7392 24458 7404
rect 24504 7401 24532 7500
rect 24489 7395 24547 7401
rect 24489 7392 24501 7395
rect 24452 7364 24501 7392
rect 24452 7352 24458 7364
rect 24489 7361 24501 7364
rect 24535 7361 24547 7395
rect 24489 7355 24547 7361
rect 24121 7327 24179 7333
rect 24121 7293 24133 7327
rect 24167 7324 24179 7327
rect 25314 7324 25320 7336
rect 24167 7296 25320 7324
rect 24167 7293 24179 7296
rect 24121 7287 24179 7293
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 24305 7259 24363 7265
rect 24305 7256 24317 7259
rect 23676 7228 24317 7256
rect 24305 7225 24317 7228
rect 24351 7225 24363 7259
rect 24305 7219 24363 7225
rect 20806 7188 20812 7200
rect 19904 7160 20812 7188
rect 10413 7151 10471 7157
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 21358 7148 21364 7200
rect 21416 7188 21422 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21416 7160 21833 7188
rect 21416 7148 21422 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21821 7151 21879 7157
rect 1104 7098 24840 7120
rect 1104 7046 3917 7098
rect 3969 7046 3981 7098
rect 4033 7046 4045 7098
rect 4097 7046 4109 7098
rect 4161 7046 4173 7098
rect 4225 7046 9851 7098
rect 9903 7046 9915 7098
rect 9967 7046 9979 7098
rect 10031 7046 10043 7098
rect 10095 7046 10107 7098
rect 10159 7046 15785 7098
rect 15837 7046 15849 7098
rect 15901 7046 15913 7098
rect 15965 7046 15977 7098
rect 16029 7046 16041 7098
rect 16093 7046 21719 7098
rect 21771 7046 21783 7098
rect 21835 7046 21847 7098
rect 21899 7046 21911 7098
rect 21963 7046 21975 7098
rect 22027 7046 24840 7098
rect 1104 7024 24840 7046
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3602 6984 3608 6996
rect 3375 6956 3608 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3602 6944 3608 6956
rect 3660 6944 3666 6996
rect 4890 6984 4896 6996
rect 4540 6956 4896 6984
rect 4154 6916 4160 6928
rect 2976 6888 4160 6916
rect 1578 6808 1584 6860
rect 1636 6848 1642 6860
rect 1949 6851 2007 6857
rect 1949 6848 1961 6851
rect 1636 6820 1961 6848
rect 1636 6808 1642 6820
rect 1949 6817 1961 6820
rect 1995 6817 2007 6851
rect 1949 6811 2007 6817
rect 2038 6808 2044 6860
rect 2096 6848 2102 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2096 6820 2329 6848
rect 2096 6808 2102 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2976 6792 3004 6888
rect 4154 6876 4160 6888
rect 4212 6916 4218 6928
rect 4540 6916 4568 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5534 6944 5540 6996
rect 5592 6944 5598 6996
rect 5902 6944 5908 6996
rect 5960 6984 5966 6996
rect 5960 6956 13400 6984
rect 5960 6944 5966 6956
rect 4212 6888 4568 6916
rect 4212 6876 4218 6888
rect 4540 6857 4568 6888
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 9088 6888 9597 6916
rect 9088 6876 9094 6888
rect 9585 6885 9597 6888
rect 9631 6885 9643 6919
rect 9585 6879 9643 6885
rect 10778 6876 10784 6928
rect 10836 6916 10842 6928
rect 13372 6916 13400 6956
rect 13446 6944 13452 6996
rect 13504 6984 13510 6996
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 13504 6956 13553 6984
rect 13504 6944 13510 6956
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13541 6947 13599 6953
rect 17954 6944 17960 6996
rect 18012 6944 18018 6996
rect 18598 6944 18604 6996
rect 18656 6944 18662 6996
rect 20346 6944 20352 6996
rect 20404 6944 20410 6996
rect 20717 6987 20775 6993
rect 20717 6953 20729 6987
rect 20763 6984 20775 6987
rect 20806 6984 20812 6996
rect 20763 6956 20812 6984
rect 20763 6953 20775 6956
rect 20717 6947 20775 6953
rect 20806 6944 20812 6956
rect 20864 6944 20870 6996
rect 21082 6944 21088 6996
rect 21140 6944 21146 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 22186 6984 22192 6996
rect 21324 6956 22192 6984
rect 21324 6944 21330 6956
rect 22186 6944 22192 6956
rect 22244 6944 22250 6996
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22336 6956 24164 6984
rect 22336 6944 22342 6956
rect 17972 6916 18000 6944
rect 10836 6888 12434 6916
rect 13372 6888 18000 6916
rect 10836 6876 10842 6888
rect 4525 6851 4583 6857
rect 3988 6820 4476 6848
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2222 6780 2228 6792
rect 1719 6752 2228 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2575 6753 2633 6759
rect 2575 6719 2587 6753
rect 2621 6750 2633 6753
rect 2621 6724 2636 6750
rect 2958 6740 2964 6792
rect 3016 6740 3022 6792
rect 3988 6789 4016 6820
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 2575 6713 2596 6719
rect 2590 6672 2596 6713
rect 2648 6672 2654 6724
rect 3418 6672 3424 6724
rect 3476 6712 3482 6724
rect 3476 6684 4108 6712
rect 3476 6672 3482 6684
rect 2038 6604 2044 6656
rect 2096 6644 2102 6656
rect 2608 6644 2636 6672
rect 2096 6616 2636 6644
rect 2096 6604 2102 6616
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 4080 6653 4108 6684
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3752 6616 3801 6644
rect 3752 6604 3758 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4065 6647 4123 6653
rect 4065 6613 4077 6647
rect 4111 6613 4123 6647
rect 4264 6644 4292 6743
rect 4448 6712 4476 6820
rect 4525 6817 4537 6851
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 7558 6848 7564 6860
rect 6788 6820 7564 6848
rect 6788 6808 6794 6820
rect 7558 6808 7564 6820
rect 7616 6808 7622 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6848 9183 6851
rect 9490 6848 9496 6860
rect 9171 6820 9496 6848
rect 9171 6817 9183 6820
rect 9125 6811 9183 6817
rect 4799 6783 4857 6789
rect 4799 6749 4811 6783
rect 4845 6780 4857 6783
rect 6178 6780 6184 6792
rect 4845 6752 6184 6780
rect 4845 6749 4857 6752
rect 4799 6743 4857 6749
rect 6178 6740 6184 6752
rect 6236 6740 6242 6792
rect 8956 6724 8984 6811
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9858 6808 9864 6860
rect 9916 6808 9922 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 12406 6848 12434 6888
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12406 6820 12541 6848
rect 10042 6789 10048 6792
rect 9999 6783 10048 6789
rect 9999 6749 10011 6783
rect 10045 6749 10048 6783
rect 9999 6743 10048 6749
rect 10042 6740 10048 6743
rect 10100 6740 10106 6792
rect 8386 6712 8392 6724
rect 4448 6684 8392 6712
rect 8386 6672 8392 6684
rect 8444 6672 8450 6724
rect 8938 6672 8944 6724
rect 8996 6672 9002 6724
rect 12406 6712 12434 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 17862 6848 17868 6860
rect 15436 6820 17868 6848
rect 15436 6808 15442 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 20364 6848 20392 6944
rect 20622 6876 20628 6928
rect 20680 6916 20686 6928
rect 22649 6919 22707 6925
rect 22649 6916 22661 6919
rect 20680 6888 22661 6916
rect 20680 6876 20686 6888
rect 22649 6885 22661 6888
rect 22695 6885 22707 6919
rect 22649 6879 22707 6885
rect 22738 6876 22744 6928
rect 22796 6876 22802 6928
rect 22005 6851 22063 6857
rect 20364 6820 21036 6848
rect 12802 6780 12808 6792
rect 12763 6752 12808 6780
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18840 6752 19196 6780
rect 18840 6740 18846 6752
rect 13262 6712 13268 6724
rect 12406 6684 13268 6712
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 19168 6656 19196 6752
rect 19334 6740 19340 6792
rect 19392 6740 19398 6792
rect 19518 6740 19524 6792
rect 19576 6780 19582 6792
rect 19611 6783 19669 6789
rect 19611 6780 19623 6783
rect 19576 6752 19623 6780
rect 19576 6740 19582 6752
rect 19611 6749 19623 6752
rect 19657 6749 19669 6783
rect 20530 6780 20536 6792
rect 19611 6743 19669 6749
rect 19720 6752 20536 6780
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 4264 6616 10793 6644
rect 4065 6607 4123 6613
rect 10781 6613 10793 6616
rect 10827 6613 10839 6647
rect 10781 6607 10839 6613
rect 17678 6604 17684 6656
rect 17736 6644 17742 6656
rect 18046 6644 18052 6656
rect 17736 6616 18052 6644
rect 17736 6604 17742 6616
rect 18046 6604 18052 6616
rect 18104 6604 18110 6656
rect 19150 6604 19156 6656
rect 19208 6604 19214 6656
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 19720 6644 19748 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 21008 6789 21036 6820
rect 22005 6817 22017 6851
rect 22051 6817 22063 6851
rect 22005 6811 22063 6817
rect 20993 6783 21051 6789
rect 20993 6749 21005 6783
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6780 21235 6783
rect 21358 6780 21364 6792
rect 21223 6752 21364 6780
rect 21223 6749 21235 6752
rect 21177 6743 21235 6749
rect 21358 6740 21364 6752
rect 21416 6740 21422 6792
rect 21450 6740 21456 6792
rect 21508 6740 21514 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21910 6780 21916 6792
rect 21591 6752 21916 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 20916 6712 20944 6740
rect 21082 6712 21088 6724
rect 20916 6684 21088 6712
rect 21082 6672 21088 6684
rect 21140 6672 21146 6724
rect 19484 6616 19748 6644
rect 19484 6604 19490 6616
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21266 6644 21272 6656
rect 20588 6616 21272 6644
rect 20588 6604 20594 6616
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 21634 6604 21640 6656
rect 21692 6644 21698 6656
rect 21729 6647 21787 6653
rect 21729 6644 21741 6647
rect 21692 6616 21741 6644
rect 21692 6604 21698 6616
rect 21729 6613 21741 6616
rect 21775 6613 21787 6647
rect 22020 6644 22048 6811
rect 22186 6740 22192 6792
rect 22244 6740 22250 6792
rect 22756 6789 22784 6876
rect 24026 6808 24032 6860
rect 24084 6808 24090 6860
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 23198 6740 23204 6792
rect 23256 6740 23262 6792
rect 23382 6740 23388 6792
rect 23440 6740 23446 6792
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 22278 6672 22284 6724
rect 22336 6712 22342 6724
rect 23216 6712 23244 6740
rect 23492 6712 23520 6743
rect 23566 6740 23572 6792
rect 23624 6780 23630 6792
rect 24136 6789 24164 6956
rect 23937 6783 23995 6789
rect 23937 6780 23949 6783
rect 23624 6752 23949 6780
rect 23624 6740 23630 6752
rect 23937 6749 23949 6752
rect 23983 6749 23995 6783
rect 23937 6743 23995 6749
rect 24121 6783 24179 6789
rect 24121 6749 24133 6783
rect 24167 6749 24179 6783
rect 24121 6743 24179 6749
rect 22336 6684 22968 6712
rect 23216 6684 23520 6712
rect 22336 6672 22342 6684
rect 22940 6656 22968 6684
rect 22830 6644 22836 6656
rect 22020 6616 22836 6644
rect 21729 6607 21787 6613
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 22922 6604 22928 6656
rect 22980 6604 22986 6656
rect 23198 6604 23204 6656
rect 23256 6604 23262 6656
rect 23569 6647 23627 6653
rect 23569 6613 23581 6647
rect 23615 6644 23627 6647
rect 24026 6644 24032 6656
rect 23615 6616 24032 6644
rect 23615 6613 23627 6616
rect 23569 6607 23627 6613
rect 24026 6604 24032 6616
rect 24084 6604 24090 6656
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 3421 6443 3479 6449
rect 3421 6440 3433 6443
rect 1360 6412 3433 6440
rect 1360 6400 1366 6412
rect 3421 6409 3433 6412
rect 3467 6409 3479 6443
rect 3421 6403 3479 6409
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 4706 6440 4712 6452
rect 3660 6412 4712 6440
rect 3660 6400 3666 6412
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 5626 6400 5632 6452
rect 5684 6400 5690 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 5736 6412 8309 6440
rect 1210 6332 1216 6384
rect 1268 6372 1274 6384
rect 2593 6375 2651 6381
rect 2593 6372 2605 6375
rect 1268 6344 2605 6372
rect 1268 6332 1274 6344
rect 2593 6341 2605 6344
rect 2639 6341 2651 6375
rect 2593 6335 2651 6341
rect 2682 6332 2688 6384
rect 2740 6372 2746 6384
rect 3234 6372 3240 6384
rect 2740 6344 3240 6372
rect 2740 6332 2746 6344
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 3375 6344 4660 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 2130 6304 2136 6316
rect 1535 6276 2136 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 3786 6304 3792 6316
rect 2823 6276 3792 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 2240 6236 2268 6267
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4154 6304 4160 6316
rect 4019 6276 4160 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4247 6307 4305 6313
rect 4247 6273 4259 6307
rect 4293 6304 4305 6307
rect 4338 6304 4344 6316
rect 4293 6276 4344 6304
rect 4293 6273 4305 6276
rect 4247 6267 4305 6273
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4632 6236 4660 6344
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5644 6304 5672 6400
rect 5583 6276 5672 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 2240 6208 3924 6236
rect 4632 6208 5672 6236
rect 1302 6128 1308 6180
rect 1360 6168 1366 6180
rect 1360 6140 2774 6168
rect 1360 6128 1366 6140
rect 1394 6060 1400 6112
rect 1452 6100 1458 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1452 6072 1593 6100
rect 1452 6060 1458 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 2746 6100 2774 6140
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2746 6072 2881 6100
rect 1581 6063 1639 6069
rect 2869 6069 2881 6072
rect 2915 6069 2927 6103
rect 3896 6100 3924 6208
rect 5644 6177 5672 6208
rect 5629 6171 5687 6177
rect 4632 6140 5488 6168
rect 4632 6100 4660 6140
rect 3896 6072 4660 6100
rect 2869 6063 2927 6069
rect 5350 6060 5356 6112
rect 5408 6060 5414 6112
rect 5460 6100 5488 6140
rect 5629 6137 5641 6171
rect 5675 6137 5687 6171
rect 5629 6131 5687 6137
rect 5736 6100 5764 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 9490 6440 9496 6452
rect 8297 6403 8355 6409
rect 9048 6412 9496 6440
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 6086 6264 6092 6316
rect 6144 6264 6150 6316
rect 6270 6264 6276 6316
rect 6328 6304 6334 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6328 6276 6377 6304
rect 6328 6264 6334 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7374 6264 7380 6316
rect 7432 6313 7438 6316
rect 7432 6307 7460 6313
rect 7448 6273 7460 6307
rect 7432 6267 7460 6273
rect 7432 6264 7438 6267
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 9048 6313 9076 6412
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10042 6440 10048 6452
rect 9916 6412 10048 6440
rect 9916 6400 9922 6412
rect 10042 6400 10048 6412
rect 10100 6440 10106 6452
rect 10686 6440 10692 6452
rect 10100 6412 10692 6440
rect 10100 6400 10106 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 12434 6440 12440 6452
rect 11716 6412 12440 6440
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8251 6276 8493 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 9033 6307 9091 6313
rect 9033 6273 9045 6307
rect 9079 6273 9091 6307
rect 9033 6267 9091 6273
rect 9766 6264 9772 6316
rect 9824 6264 9830 6316
rect 9858 6264 9864 6316
rect 9916 6313 9922 6316
rect 9916 6307 9944 6313
rect 9932 6273 9944 6307
rect 9916 6267 9944 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6304 11575 6307
rect 11606 6304 11612 6316
rect 11563 6276 11612 6304
rect 11563 6273 11575 6276
rect 11517 6267 11575 6273
rect 9916 6264 9922 6267
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 5902 6196 5908 6248
rect 5960 6236 5966 6248
rect 6178 6236 6184 6248
rect 5960 6208 6184 6236
rect 5960 6196 5966 6208
rect 6178 6196 6184 6208
rect 6236 6236 6242 6248
rect 8849 6239 8907 6245
rect 6236 6208 6868 6236
rect 6236 6196 6242 6208
rect 6840 6180 6868 6208
rect 6932 6208 7972 6236
rect 6822 6128 6828 6180
rect 6880 6128 6886 6180
rect 6932 6112 6960 6208
rect 7006 6128 7012 6180
rect 7064 6128 7070 6180
rect 5460 6072 5764 6100
rect 5902 6060 5908 6112
rect 5960 6060 5966 6112
rect 6914 6060 6920 6112
rect 6972 6060 6978 6112
rect 7944 6100 7972 6208
rect 8849 6205 8861 6239
rect 8895 6236 8907 6239
rect 8938 6236 8944 6248
rect 8895 6208 8944 6236
rect 8895 6205 8907 6208
rect 8849 6199 8907 6205
rect 8864 6168 8892 6199
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 10045 6239 10103 6245
rect 10045 6205 10057 6239
rect 10091 6236 10103 6239
rect 10226 6236 10232 6248
rect 10091 6208 10232 6236
rect 10091 6205 10103 6208
rect 10045 6199 10103 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 10594 6196 10600 6248
rect 10652 6236 10658 6248
rect 11716 6245 11744 6412
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13964 6412 14473 6440
rect 13964 6400 13970 6412
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 16758 6440 16764 6452
rect 15620 6412 16764 6440
rect 15620 6400 15626 6412
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 17920 6412 17969 6440
rect 17920 6400 17926 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 20625 6443 20683 6449
rect 20625 6409 20637 6443
rect 20671 6440 20683 6443
rect 21450 6440 21456 6452
rect 20671 6412 21456 6440
rect 20671 6409 20683 6412
rect 20625 6403 20683 6409
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 22186 6440 22192 6452
rect 21744 6412 22192 6440
rect 21269 6375 21327 6381
rect 13280 6344 20668 6372
rect 12526 6264 12532 6316
rect 12584 6313 12590 6316
rect 12584 6307 12633 6313
rect 12584 6273 12587 6307
rect 12621 6273 12633 6307
rect 12584 6267 12633 6273
rect 12584 6264 12590 6267
rect 12710 6264 12716 6316
rect 12768 6264 12774 6316
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 10652 6208 11713 6236
rect 10652 6196 10658 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11940 6208 12449 6236
rect 11940 6196 11946 6208
rect 12437 6205 12449 6208
rect 12483 6236 12495 6239
rect 13280 6236 13308 6344
rect 20640 6316 20668 6344
rect 21269 6341 21281 6375
rect 21315 6372 21327 6375
rect 21744 6372 21772 6412
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 22738 6400 22744 6452
rect 22796 6440 22802 6452
rect 23293 6443 23351 6449
rect 23293 6440 23305 6443
rect 22796 6412 23305 6440
rect 22796 6400 22802 6412
rect 23293 6409 23305 6412
rect 23339 6409 23351 6443
rect 23293 6403 23351 6409
rect 23382 6400 23388 6452
rect 23440 6440 23446 6452
rect 23937 6443 23995 6449
rect 23937 6440 23949 6443
rect 23440 6412 23949 6440
rect 23440 6400 23446 6412
rect 23937 6409 23949 6412
rect 23983 6409 23995 6443
rect 23937 6403 23995 6409
rect 24305 6443 24363 6449
rect 24305 6409 24317 6443
rect 24351 6440 24363 6443
rect 24394 6440 24400 6452
rect 24351 6412 24400 6440
rect 24351 6409 24363 6412
rect 24305 6403 24363 6409
rect 24394 6400 24400 6412
rect 24452 6400 24458 6452
rect 25222 6372 25228 6384
rect 21315 6344 21772 6372
rect 22020 6344 23520 6372
rect 21315 6341 21327 6344
rect 21269 6335 21327 6341
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13691 6307 13749 6313
rect 13691 6304 13703 6307
rect 13412 6276 13703 6304
rect 13412 6264 13418 6276
rect 13691 6273 13703 6276
rect 13737 6273 13749 6307
rect 13691 6267 13749 6273
rect 15195 6307 15253 6313
rect 15195 6273 15207 6307
rect 15241 6304 15253 6307
rect 15286 6304 15292 6316
rect 15241 6276 15292 6304
rect 15241 6273 15253 6276
rect 15195 6267 15253 6273
rect 15286 6264 15292 6276
rect 15344 6304 15350 6316
rect 17681 6307 17739 6313
rect 15344 6276 16528 6304
rect 15344 6264 15350 6276
rect 12483 6208 13308 6236
rect 13449 6239 13507 6245
rect 12483 6205 12495 6208
rect 12437 6199 12495 6205
rect 13449 6205 13461 6239
rect 13495 6205 13507 6239
rect 13449 6199 13507 6205
rect 9398 6168 9404 6180
rect 8864 6140 9404 6168
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 9490 6128 9496 6180
rect 9548 6128 9554 6180
rect 12158 6128 12164 6180
rect 12216 6128 12222 6180
rect 13262 6128 13268 6180
rect 13320 6168 13326 6180
rect 13464 6168 13492 6199
rect 14734 6196 14740 6248
rect 14792 6236 14798 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14792 6208 14933 6236
rect 14792 6196 14798 6208
rect 14921 6205 14933 6208
rect 14967 6205 14979 6239
rect 14921 6199 14979 6205
rect 13320 6140 13492 6168
rect 13320 6128 13326 6140
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 7944 6072 10701 6100
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10778 6060 10784 6112
rect 10836 6100 10842 6112
rect 12434 6100 12440 6112
rect 10836 6072 12440 6100
rect 10836 6060 10842 6072
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 12676 6072 13369 6100
rect 12676 6060 12682 6072
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 15933 6103 15991 6109
rect 15933 6069 15945 6103
rect 15979 6100 15991 6103
rect 16206 6100 16212 6112
rect 15979 6072 16212 6100
rect 15979 6069 15991 6072
rect 15933 6063 15991 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16500 6100 16528 6276
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 18230 6304 18236 6316
rect 17727 6276 18236 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20622 6264 20628 6316
rect 20680 6264 20686 6316
rect 20809 6307 20867 6313
rect 20809 6273 20821 6307
rect 20855 6304 20867 6307
rect 20898 6304 20904 6316
rect 20855 6276 20904 6304
rect 20855 6273 20867 6276
rect 20809 6267 20867 6273
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 21082 6264 21088 6316
rect 21140 6264 21146 6316
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21223 6302 21312 6304
rect 21358 6302 21364 6316
rect 21223 6276 21364 6302
rect 21223 6273 21235 6276
rect 21284 6274 21364 6276
rect 21177 6267 21235 6273
rect 21358 6264 21364 6274
rect 21416 6264 21422 6316
rect 21450 6264 21456 6316
rect 21508 6304 21514 6316
rect 21637 6307 21695 6313
rect 21637 6304 21649 6307
rect 21508 6276 21649 6304
rect 21508 6264 21514 6276
rect 21637 6273 21649 6276
rect 21683 6273 21695 6307
rect 22020 6304 22048 6344
rect 21637 6267 21695 6273
rect 21744 6276 22048 6304
rect 22095 6307 22153 6313
rect 17957 6239 18015 6245
rect 17957 6205 17969 6239
rect 18003 6236 18015 6239
rect 18414 6236 18420 6248
rect 18003 6208 18420 6236
rect 18003 6205 18015 6208
rect 17957 6199 18015 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 21744 6236 21772 6276
rect 22095 6273 22107 6307
rect 22141 6304 22153 6307
rect 22462 6304 22468 6316
rect 22141 6276 22468 6304
rect 22141 6273 22153 6276
rect 22095 6267 22153 6273
rect 22462 6264 22468 6276
rect 22520 6264 22526 6316
rect 22830 6264 22836 6316
rect 22888 6304 22894 6316
rect 23492 6313 23520 6344
rect 24044 6344 25228 6372
rect 23201 6307 23259 6313
rect 23201 6304 23213 6307
rect 22888 6276 23213 6304
rect 22888 6264 22894 6276
rect 23201 6273 23213 6276
rect 23247 6273 23259 6307
rect 23201 6267 23259 6273
rect 23385 6307 23443 6313
rect 23385 6273 23397 6307
rect 23431 6273 23443 6307
rect 23385 6267 23443 6273
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 21284 6228 21772 6236
rect 21100 6208 21772 6228
rect 21100 6200 21312 6208
rect 17773 6171 17831 6177
rect 17773 6137 17785 6171
rect 17819 6168 17831 6171
rect 18138 6168 18144 6180
rect 17819 6140 18144 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 20349 6171 20407 6177
rect 20349 6137 20361 6171
rect 20395 6168 20407 6171
rect 21100 6168 21128 6200
rect 21818 6196 21824 6248
rect 21876 6196 21882 6248
rect 22848 6177 22876 6264
rect 23400 6236 23428 6267
rect 23750 6264 23756 6316
rect 23808 6264 23814 6316
rect 24044 6313 24072 6344
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 24029 6307 24087 6313
rect 24029 6273 24041 6307
rect 24075 6273 24087 6307
rect 24029 6267 24087 6273
rect 24486 6264 24492 6316
rect 24544 6264 24550 6316
rect 23216 6208 23428 6236
rect 20395 6140 21128 6168
rect 21453 6171 21511 6177
rect 20395 6137 20407 6140
rect 20349 6131 20407 6137
rect 21453 6137 21465 6171
rect 21499 6137 21511 6171
rect 21453 6131 21511 6137
rect 22833 6171 22891 6177
rect 22833 6137 22845 6171
rect 22879 6137 22891 6171
rect 22833 6131 22891 6137
rect 17862 6100 17868 6112
rect 16500 6072 17868 6100
rect 17862 6060 17868 6072
rect 17920 6060 17926 6112
rect 20898 6060 20904 6112
rect 20956 6060 20962 6112
rect 21266 6060 21272 6112
rect 21324 6100 21330 6112
rect 21468 6100 21496 6131
rect 21324 6072 21496 6100
rect 21324 6060 21330 6072
rect 21634 6060 21640 6112
rect 21692 6100 21698 6112
rect 23216 6100 23244 6208
rect 24213 6171 24271 6177
rect 24213 6168 24225 6171
rect 23492 6140 24225 6168
rect 21692 6072 23244 6100
rect 21692 6060 21698 6072
rect 23290 6060 23296 6112
rect 23348 6100 23354 6112
rect 23492 6100 23520 6140
rect 24213 6137 24225 6140
rect 24259 6137 24271 6171
rect 24213 6131 24271 6137
rect 23348 6072 23520 6100
rect 23348 6060 23354 6072
rect 23566 6060 23572 6112
rect 23624 6060 23630 6112
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 1762 5856 1768 5908
rect 1820 5856 1826 5908
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 3237 5899 3295 5905
rect 3237 5896 3249 5899
rect 2746 5868 3249 5896
rect 1026 5788 1032 5840
rect 1084 5828 1090 5840
rect 2746 5828 2774 5868
rect 3237 5865 3249 5868
rect 3283 5865 3295 5899
rect 3237 5859 3295 5865
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 5350 5896 5356 5908
rect 3936 5868 5356 5896
rect 3936 5856 3942 5868
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 5537 5899 5595 5905
rect 5537 5865 5549 5899
rect 5583 5865 5595 5899
rect 5537 5859 5595 5865
rect 1084 5800 2774 5828
rect 1084 5788 1090 5800
rect 3326 5788 3332 5840
rect 3384 5828 3390 5840
rect 3384 5800 4016 5828
rect 3384 5788 3390 5800
rect 3694 5760 3700 5772
rect 1688 5732 3700 5760
rect 1688 5701 1716 5732
rect 3694 5720 3700 5732
rect 3752 5720 3758 5772
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 2314 5652 2320 5704
rect 2372 5652 2378 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3878 5692 3884 5704
rect 3191 5664 3884 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 3988 5701 4016 5800
rect 4706 5788 4712 5840
rect 4764 5828 4770 5840
rect 5552 5828 5580 5859
rect 5902 5856 5908 5908
rect 5960 5856 5966 5908
rect 6362 5896 6368 5908
rect 6104 5868 6368 5896
rect 4764 5800 5580 5828
rect 4764 5788 4770 5800
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4154 5692 4160 5704
rect 4019 5664 4160 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 4246 5652 4252 5704
rect 4304 5652 4310 5704
rect 5920 5692 5948 5856
rect 6104 5769 6132 5868
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 7101 5899 7159 5905
rect 6604 5868 7052 5896
rect 6604 5856 6610 5868
rect 7024 5828 7052 5868
rect 7101 5865 7113 5899
rect 7147 5896 7159 5899
rect 7466 5896 7472 5908
rect 7147 5868 7472 5896
rect 7147 5865 7159 5868
rect 7101 5859 7159 5865
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 8481 5899 8539 5905
rect 7576 5868 8432 5896
rect 7576 5828 7604 5868
rect 7024 5800 7604 5828
rect 8404 5828 8432 5868
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 9490 5896 9496 5908
rect 8527 5868 9496 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 10594 5896 10600 5908
rect 9968 5868 10600 5896
rect 9968 5828 9996 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 12158 5896 12164 5908
rect 10919 5868 12164 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12710 5896 12716 5908
rect 12299 5868 12716 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 16206 5896 16212 5908
rect 16040 5868 16212 5896
rect 8404 5800 9996 5828
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 15470 5828 15476 5840
rect 12492 5800 15476 5828
rect 12492 5788 12498 5800
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 15562 5788 15568 5840
rect 15620 5828 15626 5840
rect 15933 5831 15991 5837
rect 15620 5800 15698 5828
rect 15620 5788 15626 5800
rect 6089 5763 6147 5769
rect 6089 5729 6101 5763
rect 6135 5729 6147 5763
rect 6089 5723 6147 5729
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 7469 5763 7527 5769
rect 7469 5760 7481 5763
rect 6880 5732 7481 5760
rect 6880 5720 6886 5732
rect 7469 5729 7481 5732
rect 7515 5729 7527 5763
rect 7469 5723 7527 5729
rect 9214 5720 9220 5772
rect 9272 5760 9278 5772
rect 9272 5732 9904 5760
rect 9272 5720 9278 5732
rect 9876 5704 9904 5732
rect 4356 5664 5948 5692
rect 7743 5695 7801 5701
rect 6347 5665 6405 5671
rect 2593 5627 2651 5633
rect 2593 5593 2605 5627
rect 2639 5624 2651 5627
rect 4356 5624 4384 5664
rect 2639 5596 4384 5624
rect 2639 5593 2651 5596
rect 2593 5587 2651 5593
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 5445 5627 5503 5633
rect 5445 5624 5457 5627
rect 5408 5596 5457 5624
rect 5408 5584 5414 5596
rect 5445 5593 5457 5596
rect 5491 5593 5503 5627
rect 6347 5631 6359 5665
rect 6393 5662 6405 5665
rect 6393 5631 6406 5662
rect 7743 5661 7755 5695
rect 7789 5692 7801 5695
rect 9582 5692 9588 5704
rect 7789 5664 9588 5692
rect 7789 5661 7801 5664
rect 7743 5655 7801 5661
rect 8588 5636 8616 5664
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10135 5695 10193 5701
rect 10135 5692 10147 5695
rect 10100 5664 10147 5692
rect 10100 5652 10106 5664
rect 10135 5661 10147 5664
rect 10181 5692 10193 5695
rect 10778 5692 10784 5704
rect 10181 5664 10784 5692
rect 10181 5661 10193 5664
rect 10135 5655 10193 5661
rect 10778 5652 10784 5664
rect 10836 5652 10842 5704
rect 10962 5652 10968 5704
rect 11020 5692 11026 5704
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11020 5664 11253 5692
rect 11020 5652 11026 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 6347 5625 6406 5631
rect 6378 5624 6406 5625
rect 6378 5596 6960 5624
rect 5445 5587 5503 5593
rect 2866 5516 2872 5568
rect 2924 5516 2930 5568
rect 4982 5516 4988 5568
rect 5040 5516 5046 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 6546 5556 6552 5568
rect 5776 5528 6552 5556
rect 5776 5516 5782 5528
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 6932 5556 6960 5596
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 7374 5624 7380 5636
rect 7064 5596 7380 5624
rect 7064 5584 7070 5596
rect 7374 5584 7380 5596
rect 7432 5584 7438 5636
rect 8386 5584 8392 5636
rect 8444 5584 8450 5636
rect 8570 5584 8576 5636
rect 8628 5584 8634 5636
rect 9398 5584 9404 5636
rect 9456 5624 9462 5636
rect 11054 5624 11060 5636
rect 9456 5596 11060 5624
rect 9456 5584 9462 5596
rect 11054 5584 11060 5596
rect 11112 5584 11118 5636
rect 11256 5624 11284 5655
rect 11514 5652 11520 5704
rect 11572 5692 11578 5704
rect 12526 5692 12532 5704
rect 11572 5664 11615 5692
rect 11716 5664 12532 5692
rect 11572 5652 11578 5664
rect 11716 5624 11744 5664
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5692 15347 5695
rect 15378 5692 15384 5704
rect 15335 5664 15384 5692
rect 15335 5661 15347 5664
rect 15289 5655 15347 5661
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5692 15531 5695
rect 15670 5692 15698 5800
rect 15933 5797 15945 5831
rect 15979 5828 15991 5831
rect 16040 5828 16068 5868
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 18230 5856 18236 5908
rect 18288 5856 18294 5908
rect 19518 5896 19524 5908
rect 19260 5868 19524 5896
rect 15979 5800 16068 5828
rect 15979 5797 15991 5800
rect 15933 5791 15991 5797
rect 16298 5720 16304 5772
rect 16356 5769 16362 5772
rect 16356 5763 16384 5769
rect 16372 5729 16384 5763
rect 16356 5723 16384 5729
rect 16485 5763 16543 5769
rect 16485 5729 16497 5763
rect 16531 5760 16543 5763
rect 17126 5760 17132 5772
rect 16531 5732 17132 5760
rect 16531 5729 16543 5732
rect 16485 5723 16543 5729
rect 16356 5720 16362 5723
rect 17126 5720 17132 5732
rect 17184 5720 17190 5772
rect 19260 5769 19288 5868
rect 19518 5856 19524 5868
rect 19576 5856 19582 5908
rect 21082 5856 21088 5908
rect 21140 5856 21146 5908
rect 21174 5856 21180 5908
rect 21232 5856 21238 5908
rect 21358 5856 21364 5908
rect 21416 5896 21422 5908
rect 21453 5899 21511 5905
rect 21453 5896 21465 5899
rect 21416 5868 21465 5896
rect 21416 5856 21422 5868
rect 21453 5865 21465 5868
rect 21499 5865 21511 5899
rect 22925 5899 22983 5905
rect 22925 5896 22937 5899
rect 21453 5859 21511 5865
rect 21560 5868 22937 5896
rect 21100 5828 21128 5856
rect 21560 5828 21588 5868
rect 22925 5865 22937 5868
rect 22971 5865 22983 5899
rect 22925 5859 22983 5865
rect 23566 5856 23572 5908
rect 23624 5856 23630 5908
rect 21100 5800 21588 5828
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 15519 5664 15698 5692
rect 15519 5661 15531 5664
rect 15473 5655 15531 5661
rect 13906 5624 13912 5636
rect 11256 5596 11744 5624
rect 12452 5596 13912 5624
rect 7650 5556 7656 5568
rect 6932 5528 7656 5556
rect 7650 5516 7656 5528
rect 7708 5516 7714 5568
rect 8404 5556 8432 5584
rect 12452 5556 12480 5596
rect 13906 5584 13912 5596
rect 13964 5584 13970 5636
rect 14918 5584 14924 5636
rect 14976 5624 14982 5636
rect 15488 5624 15516 5655
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 17221 5695 17279 5701
rect 17221 5661 17233 5695
rect 17267 5661 17279 5695
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17221 5655 17279 5661
rect 14976 5596 15516 5624
rect 17236 5624 17264 5655
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 19260 5692 19288 5723
rect 20162 5720 20168 5772
rect 20220 5760 20226 5772
rect 20220 5732 21588 5760
rect 20220 5720 20226 5732
rect 19487 5695 19545 5701
rect 19487 5692 19499 5695
rect 17696 5664 19288 5692
rect 19352 5664 19499 5692
rect 17696 5636 17724 5664
rect 17678 5624 17684 5636
rect 17236 5596 17684 5624
rect 14976 5584 14982 5596
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 19352 5624 19380 5664
rect 19487 5661 19499 5664
rect 19533 5661 19545 5695
rect 19487 5655 19545 5661
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20404 5664 20913 5692
rect 20404 5652 20410 5664
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 20990 5652 20996 5704
rect 21048 5652 21054 5704
rect 21560 5701 21588 5732
rect 21269 5695 21327 5701
rect 21269 5661 21281 5695
rect 21315 5661 21327 5695
rect 21269 5655 21327 5661
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 22370 5692 22376 5704
rect 21591 5664 22376 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 17920 5596 19380 5624
rect 21284 5624 21312 5655
rect 22370 5652 22376 5664
rect 22428 5692 22434 5704
rect 22554 5692 22560 5704
rect 22428 5664 22560 5692
rect 22428 5652 22434 5664
rect 22554 5652 22560 5664
rect 22612 5652 22618 5704
rect 23290 5652 23296 5704
rect 23348 5652 23354 5704
rect 23584 5701 23612 5856
rect 23569 5695 23627 5701
rect 23569 5661 23581 5695
rect 23615 5661 23627 5695
rect 23569 5655 23627 5661
rect 23750 5652 23756 5704
rect 23808 5692 23814 5704
rect 23937 5695 23995 5701
rect 23937 5692 23949 5695
rect 23808 5664 23949 5692
rect 23808 5652 23814 5664
rect 23937 5661 23949 5664
rect 23983 5661 23995 5695
rect 23937 5655 23995 5661
rect 21818 5633 21824 5636
rect 21284 5596 21772 5624
rect 17920 5584 17926 5596
rect 8404 5528 12480 5556
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 17129 5559 17187 5565
rect 17129 5556 17141 5559
rect 16632 5528 17141 5556
rect 16632 5516 16638 5528
rect 17129 5525 17141 5528
rect 17175 5525 17187 5559
rect 17129 5519 17187 5525
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 19392 5528 20269 5556
rect 19392 5516 19398 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 20898 5556 20904 5568
rect 20763 5528 20904 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 21744 5556 21772 5596
rect 21812 5587 21824 5633
rect 21876 5624 21882 5636
rect 21876 5596 21912 5624
rect 21818 5584 21824 5587
rect 21876 5584 21882 5596
rect 22094 5584 22100 5636
rect 22152 5624 22158 5636
rect 22646 5624 22652 5636
rect 22152 5596 22652 5624
rect 22152 5584 22158 5596
rect 22646 5584 22652 5596
rect 22704 5584 22710 5636
rect 23382 5584 23388 5636
rect 23440 5624 23446 5636
rect 24213 5627 24271 5633
rect 24213 5624 24225 5627
rect 23440 5596 24225 5624
rect 23440 5584 23446 5596
rect 24213 5593 24225 5596
rect 24259 5593 24271 5627
rect 24213 5587 24271 5593
rect 22186 5556 22192 5568
rect 21744 5528 22192 5556
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 2130 5312 2136 5364
rect 2188 5352 2194 5364
rect 2590 5352 2596 5364
rect 2188 5324 2596 5352
rect 2188 5312 2194 5324
rect 2590 5312 2596 5324
rect 2648 5312 2654 5364
rect 2682 5312 2688 5364
rect 2740 5352 2746 5364
rect 3326 5352 3332 5364
rect 2740 5324 3332 5352
rect 2740 5312 2746 5324
rect 3326 5312 3332 5324
rect 3384 5352 3390 5364
rect 5258 5352 5264 5364
rect 3384 5324 5264 5352
rect 3384 5312 3390 5324
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5868 5324 6193 5352
rect 5868 5312 5874 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 6181 5315 6239 5321
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 10226 5312 10232 5364
rect 10284 5312 10290 5364
rect 10870 5312 10876 5364
rect 10928 5312 10934 5364
rect 12342 5352 12348 5364
rect 11990 5324 12348 5352
rect 10594 5284 10600 5296
rect 1412 5256 2820 5284
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1412 5225 1440 5256
rect 2792 5225 2820 5256
rect 9508 5256 10600 5284
rect 9508 5255 9536 5256
rect 9475 5249 9536 5255
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 1671 5219 1729 5225
rect 1671 5185 1683 5219
rect 1717 5216 1729 5219
rect 2777 5219 2835 5225
rect 1717 5188 2268 5216
rect 1717 5185 1729 5188
rect 1671 5179 1729 5185
rect 2240 5080 2268 5188
rect 2777 5185 2789 5219
rect 2823 5216 2835 5219
rect 2958 5216 2964 5228
rect 2823 5188 2964 5216
rect 2823 5185 2835 5188
rect 2777 5179 2835 5185
rect 2958 5176 2964 5188
rect 3016 5176 3022 5228
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4430 5216 4436 5228
rect 4387 5188 4436 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4430 5176 4436 5188
rect 4488 5216 4494 5228
rect 4488 5188 4752 5216
rect 4488 5176 4494 5188
rect 4522 5108 4528 5160
rect 4580 5108 4586 5160
rect 4724 5148 4752 5188
rect 5258 5176 5264 5228
rect 5316 5176 5322 5228
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6639 5219 6697 5225
rect 6639 5185 6651 5219
rect 6685 5216 6697 5219
rect 6730 5216 6736 5228
rect 6685 5188 6736 5216
rect 6685 5185 6697 5188
rect 6639 5179 6697 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 9475 5215 9487 5249
rect 9521 5218 9536 5249
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 10888 5284 10916 5312
rect 10652 5256 10916 5284
rect 10652 5244 10658 5256
rect 9521 5215 9533 5218
rect 9475 5209 9533 5215
rect 9858 5176 9864 5228
rect 9916 5176 9922 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10870 5216 10876 5228
rect 10560 5188 10876 5216
rect 10560 5176 10566 5188
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 4890 5148 4896 5160
rect 4724 5120 4896 5148
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 4982 5108 4988 5160
rect 5040 5108 5046 5160
rect 5074 5108 5080 5160
rect 5132 5148 5138 5160
rect 5378 5151 5436 5157
rect 5378 5148 5390 5151
rect 5132 5120 5390 5148
rect 5132 5108 5138 5120
rect 5378 5117 5390 5120
rect 5424 5117 5436 5151
rect 5378 5111 5436 5117
rect 8938 5108 8944 5160
rect 8996 5148 9002 5160
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 8996 5120 9229 5148
rect 8996 5108 9002 5120
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9876 5148 9904 5176
rect 10962 5148 10968 5160
rect 9876 5120 10968 5148
rect 9217 5111 9275 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 4062 5080 4068 5092
rect 2240 5052 2774 5080
rect 2409 5015 2467 5021
rect 2409 4981 2421 5015
rect 2455 5012 2467 5015
rect 2498 5012 2504 5024
rect 2455 4984 2504 5012
rect 2455 4981 2467 4984
rect 2409 4975 2467 4981
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 2746 5012 2774 5052
rect 3436 5052 4068 5080
rect 3436 5012 3464 5052
rect 4062 5040 4068 5052
rect 4120 5040 4126 5092
rect 4338 5040 4344 5092
rect 4396 5080 4402 5092
rect 5092 5080 5120 5108
rect 4396 5052 5120 5080
rect 4396 5040 4402 5052
rect 2746 4984 3464 5012
rect 3602 4972 3608 5024
rect 3660 5012 3666 5024
rect 3789 5015 3847 5021
rect 3789 5012 3801 5015
rect 3660 4984 3801 5012
rect 3660 4972 3666 4984
rect 3789 4981 3801 4984
rect 3835 4981 3847 5015
rect 3789 4975 3847 4981
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 11990 5012 12018 5324
rect 12342 5312 12348 5324
rect 12400 5352 12406 5364
rect 13814 5352 13820 5364
rect 12400 5324 13820 5352
rect 12400 5312 12406 5324
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 13964 5324 16497 5352
rect 13964 5312 13970 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17681 5355 17739 5361
rect 17681 5352 17693 5355
rect 17184 5324 17693 5352
rect 17184 5312 17190 5324
rect 17681 5321 17693 5324
rect 17727 5321 17739 5355
rect 17681 5315 17739 5321
rect 18138 5312 18144 5364
rect 18196 5312 18202 5364
rect 18230 5312 18236 5364
rect 18288 5312 18294 5364
rect 18414 5312 18420 5364
rect 18472 5312 18478 5364
rect 19150 5312 19156 5364
rect 19208 5352 19214 5364
rect 21910 5352 21916 5364
rect 19208 5324 21916 5352
rect 19208 5312 19214 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 22005 5355 22063 5361
rect 22005 5321 22017 5355
rect 22051 5321 22063 5355
rect 22005 5315 22063 5321
rect 24489 5355 24547 5361
rect 24489 5321 24501 5355
rect 24535 5321 24547 5355
rect 24489 5315 24547 5321
rect 16684 5256 17632 5284
rect 16684 5228 16712 5256
rect 17604 5228 17632 5256
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 13078 5216 13084 5228
rect 12759 5188 13084 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5216 14703 5219
rect 14691 5188 15056 5216
rect 14691 5185 14703 5188
rect 14645 5179 14703 5185
rect 13814 5157 13820 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 13633 5151 13691 5157
rect 13633 5148 13645 5151
rect 12897 5111 12955 5117
rect 13464 5120 13645 5148
rect 12912 5080 12940 5111
rect 12406 5052 12940 5080
rect 12406 5024 12434 5052
rect 13354 5040 13360 5092
rect 13412 5040 13418 5092
rect 6052 4984 12018 5012
rect 6052 4972 6058 4984
rect 12342 4972 12348 5024
rect 12400 4984 12434 5024
rect 13464 5012 13492 5120
rect 13633 5117 13645 5120
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 13771 5151 13820 5157
rect 13771 5117 13783 5151
rect 13817 5117 13820 5151
rect 13771 5111 13820 5117
rect 13814 5108 13820 5111
rect 13872 5108 13878 5160
rect 13906 5108 13912 5160
rect 13964 5108 13970 5160
rect 14829 5151 14887 5157
rect 14829 5117 14841 5151
rect 14875 5148 14887 5151
rect 14918 5148 14924 5160
rect 14875 5120 14924 5148
rect 14875 5117 14887 5120
rect 14829 5111 14887 5117
rect 14844 5080 14872 5111
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15028 5148 15056 5188
rect 16666 5176 16672 5228
rect 16724 5176 16730 5228
rect 16943 5219 17001 5225
rect 16943 5185 16955 5219
rect 16989 5216 17001 5219
rect 16989 5188 17356 5216
rect 16989 5185 17001 5188
rect 16943 5179 17001 5185
rect 15378 5148 15384 5160
rect 15028 5120 15384 5148
rect 15378 5108 15384 5120
rect 15436 5108 15442 5160
rect 15562 5108 15568 5160
rect 15620 5108 15626 5160
rect 15746 5157 15752 5160
rect 15703 5151 15752 5157
rect 15703 5117 15715 5151
rect 15749 5117 15752 5151
rect 15703 5111 15752 5117
rect 15746 5108 15752 5111
rect 15804 5108 15810 5160
rect 15841 5151 15899 5157
rect 15841 5117 15853 5151
rect 15887 5148 15899 5151
rect 16390 5148 16396 5160
rect 15887 5120 16396 5148
rect 15887 5117 15899 5120
rect 15841 5111 15899 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 17328 5148 17356 5188
rect 17586 5176 17592 5228
rect 17644 5176 17650 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18049 5219 18107 5225
rect 18049 5216 18061 5219
rect 17736 5188 18061 5216
rect 17736 5176 17742 5188
rect 18049 5185 18061 5188
rect 18095 5185 18107 5219
rect 18248 5216 18276 5312
rect 18432 5256 19656 5284
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 18248 5188 18337 5216
rect 18049 5179 18107 5185
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 17770 5148 17776 5160
rect 17328 5120 17776 5148
rect 17770 5108 17776 5120
rect 17828 5148 17834 5160
rect 18432 5148 18460 5256
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 18555 5188 18644 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 17828 5120 18460 5148
rect 17828 5108 17834 5120
rect 14292 5052 14872 5080
rect 14292 5012 14320 5052
rect 15286 5040 15292 5092
rect 15344 5040 15350 5092
rect 16298 5040 16304 5092
rect 16356 5040 16362 5092
rect 17954 5040 17960 5092
rect 18012 5040 18018 5092
rect 18616 5089 18644 5188
rect 18782 5176 18788 5228
rect 18840 5176 18846 5228
rect 19150 5176 19156 5228
rect 19208 5176 19214 5228
rect 19334 5176 19340 5228
rect 19392 5176 19398 5228
rect 19503 5219 19561 5225
rect 19503 5216 19515 5219
rect 19444 5188 19515 5216
rect 18601 5083 18659 5089
rect 18601 5049 18613 5083
rect 18647 5049 18659 5083
rect 18601 5043 18659 5049
rect 19153 5083 19211 5089
rect 19153 5049 19165 5083
rect 19199 5049 19211 5083
rect 19444 5080 19472 5188
rect 19503 5185 19515 5188
rect 19549 5185 19561 5219
rect 19628 5216 19656 5256
rect 19702 5244 19708 5296
rect 19760 5284 19766 5296
rect 22020 5284 22048 5315
rect 24504 5284 24532 5315
rect 19760 5256 22048 5284
rect 22572 5256 24532 5284
rect 19760 5244 19766 5256
rect 19855 5219 19913 5225
rect 19855 5216 19867 5219
rect 19628 5188 19867 5216
rect 19503 5179 19561 5185
rect 19855 5185 19867 5188
rect 19901 5185 19913 5219
rect 19855 5179 19913 5185
rect 21174 5176 21180 5228
rect 21232 5176 21238 5228
rect 21542 5176 21548 5228
rect 21600 5176 21606 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21652 5188 21833 5216
rect 19610 5108 19616 5160
rect 19668 5108 19674 5160
rect 20990 5148 20996 5160
rect 20640 5120 20996 5148
rect 20640 5089 20668 5120
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21450 5108 21456 5160
rect 21508 5148 21514 5160
rect 21652 5148 21680 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 21910 5176 21916 5228
rect 21968 5176 21974 5228
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 22572 5225 22600 5256
rect 22097 5219 22155 5225
rect 22097 5216 22109 5219
rect 22060 5188 22109 5216
rect 22060 5176 22066 5188
rect 22097 5185 22109 5188
rect 22143 5185 22155 5219
rect 22097 5179 22155 5185
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 22646 5176 22652 5228
rect 22704 5176 22710 5228
rect 22922 5176 22928 5228
rect 22980 5216 22986 5228
rect 23365 5219 23423 5225
rect 23365 5216 23377 5219
rect 22980 5188 23377 5216
rect 22980 5176 22986 5188
rect 23365 5185 23377 5188
rect 23411 5185 23423 5219
rect 23365 5179 23423 5185
rect 21508 5120 21680 5148
rect 21508 5108 21514 5120
rect 20625 5083 20683 5089
rect 19444 5052 19656 5080
rect 19153 5043 19211 5049
rect 13464 4984 14320 5012
rect 12400 4972 12406 4984
rect 14550 4972 14556 5024
rect 14608 4972 14614 5024
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 16316 5012 16344 5040
rect 15804 4984 16344 5012
rect 17972 5012 18000 5040
rect 19168 5012 19196 5043
rect 19628 5024 19656 5052
rect 20625 5049 20637 5083
rect 20671 5049 20683 5083
rect 20625 5043 20683 5049
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 21177 5083 21235 5089
rect 21177 5080 21189 5083
rect 20772 5052 21189 5080
rect 20772 5040 20778 5052
rect 21177 5049 21189 5052
rect 21223 5049 21235 5083
rect 21928 5080 21956 5176
rect 23109 5151 23167 5157
rect 23109 5148 23121 5151
rect 22572 5120 23121 5148
rect 22572 5092 22600 5120
rect 23109 5117 23121 5120
rect 23155 5117 23167 5151
rect 23109 5111 23167 5117
rect 22281 5083 22339 5089
rect 22281 5080 22293 5083
rect 21928 5052 22293 5080
rect 21177 5043 21235 5049
rect 22281 5049 22293 5052
rect 22327 5049 22339 5083
rect 22281 5043 22339 5049
rect 22554 5040 22560 5092
rect 22612 5040 22618 5092
rect 17972 4984 19196 5012
rect 15804 4972 15810 4984
rect 19610 4972 19616 5024
rect 19668 4972 19674 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 21358 5012 21364 5024
rect 20128 4984 21364 5012
rect 20128 4972 20134 4984
rect 21358 4972 21364 4984
rect 21416 4972 21422 5024
rect 22370 4972 22376 5024
rect 22428 4972 22434 5024
rect 22462 4972 22468 5024
rect 22520 5012 22526 5024
rect 22741 5015 22799 5021
rect 22741 5012 22753 5015
rect 22520 4984 22753 5012
rect 22520 4972 22526 4984
rect 22741 4981 22753 4984
rect 22787 4981 22799 5015
rect 22741 4975 22799 4981
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 1486 4768 1492 4820
rect 1544 4768 1550 4820
rect 2314 4768 2320 4820
rect 2372 4808 2378 4820
rect 2372 4780 5488 4808
rect 2372 4768 2378 4780
rect 3786 4700 3792 4752
rect 3844 4700 3850 4752
rect 5460 4740 5488 4780
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12400 4780 13308 4808
rect 12400 4768 12434 4780
rect 12406 4740 12434 4768
rect 5460 4712 12434 4740
rect 13280 4740 13308 4780
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13412 4780 13645 4808
rect 13412 4768 13418 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 14550 4768 14556 4820
rect 14608 4768 14614 4820
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 18782 4768 18788 4820
rect 18840 4768 18846 4820
rect 19150 4768 19156 4820
rect 19208 4808 19214 4820
rect 19337 4811 19395 4817
rect 19337 4808 19349 4811
rect 19208 4780 19349 4808
rect 19208 4768 19214 4780
rect 19337 4777 19349 4780
rect 19383 4777 19395 4811
rect 19337 4771 19395 4777
rect 19610 4768 19616 4820
rect 19668 4768 19674 4820
rect 20346 4768 20352 4820
rect 20404 4768 20410 4820
rect 20714 4808 20720 4820
rect 20447 4780 20720 4808
rect 14366 4740 14372 4752
rect 13280 4712 14372 4740
rect 14366 4700 14372 4712
rect 14424 4700 14430 4752
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4672 2007 4675
rect 2130 4672 2136 4684
rect 1995 4644 2136 4672
rect 1995 4641 2007 4644
rect 1949 4635 2007 4641
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 2406 4632 2412 4684
rect 2464 4632 2470 4684
rect 2682 4632 2688 4684
rect 2740 4632 2746 4684
rect 2823 4675 2881 4681
rect 2823 4641 2835 4675
rect 2869 4672 2881 4675
rect 3510 4672 3516 4684
rect 2869 4644 3516 4672
rect 2869 4641 2881 4644
rect 2823 4635 2881 4641
rect 3510 4632 3516 4644
rect 3568 4672 3574 4684
rect 4338 4672 4344 4684
rect 3568 4644 4344 4672
rect 3568 4632 3574 4644
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 6362 4632 6368 4684
rect 6420 4632 6426 4684
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 1811 4576 1900 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 1688 4468 1716 4567
rect 1872 4548 1900 4576
rect 2958 4564 2964 4616
rect 3016 4564 3022 4616
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4262 4566 4292 4567
rect 1854 4496 1860 4548
rect 1912 4496 1918 4548
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 1688 4440 3617 4468
rect 3605 4437 3617 4440
rect 3651 4437 3663 4471
rect 3605 4431 3663 4437
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 3752 4440 4077 4468
rect 3752 4428 3758 4440
rect 4065 4437 4077 4440
rect 4111 4437 4123 4471
rect 4262 4468 4290 4566
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 4540 4536 4568 4567
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 6380 4536 6408 4632
rect 12618 4564 12624 4616
rect 12676 4564 12682 4616
rect 12802 4564 12808 4616
rect 12860 4604 12866 4616
rect 12895 4607 12953 4613
rect 12895 4604 12907 4607
rect 12860 4576 12907 4604
rect 12860 4564 12866 4576
rect 12895 4573 12907 4576
rect 12941 4604 12953 4607
rect 13538 4604 13544 4616
rect 12941 4576 13544 4604
rect 12941 4573 12953 4576
rect 12895 4567 12953 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 4396 4508 6408 4536
rect 4396 4496 4402 4508
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 14568 4536 14596 4768
rect 18877 4743 18935 4749
rect 18877 4709 18889 4743
rect 18923 4740 18935 4743
rect 20447 4740 20475 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 20993 4811 21051 4817
rect 20993 4777 21005 4811
rect 21039 4808 21051 4811
rect 21174 4808 21180 4820
rect 21039 4780 21180 4808
rect 21039 4777 21051 4780
rect 20993 4771 21051 4777
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21269 4811 21327 4817
rect 21269 4777 21281 4811
rect 21315 4808 21327 4811
rect 21542 4808 21548 4820
rect 21315 4780 21548 4808
rect 21315 4777 21327 4780
rect 21269 4771 21327 4777
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 22094 4768 22100 4820
rect 22152 4808 22158 4820
rect 22189 4811 22247 4817
rect 22189 4808 22201 4811
rect 22152 4780 22201 4808
rect 22152 4768 22158 4780
rect 22189 4777 22201 4780
rect 22235 4777 22247 4811
rect 23198 4808 23204 4820
rect 22189 4771 22247 4777
rect 22296 4780 23204 4808
rect 22296 4740 22324 4780
rect 23198 4768 23204 4780
rect 23256 4768 23262 4820
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 25406 4808 25412 4820
rect 24075 4780 25412 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 25406 4768 25412 4780
rect 25464 4768 25470 4820
rect 18923 4712 20475 4740
rect 20548 4712 22324 4740
rect 18923 4709 18935 4712
rect 18877 4703 18935 4709
rect 19334 4632 19340 4684
rect 19392 4632 19398 4684
rect 20548 4672 20576 4712
rect 20272 4644 20576 4672
rect 14734 4564 14740 4616
rect 14792 4604 14798 4616
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 14792 4576 15393 4604
rect 14792 4564 14798 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 6880 4508 14596 4536
rect 15396 4536 15424 4567
rect 15562 4564 15568 4616
rect 15620 4604 15626 4616
rect 15655 4607 15713 4613
rect 15655 4604 15667 4607
rect 15620 4576 15667 4604
rect 15620 4564 15626 4576
rect 15655 4573 15667 4576
rect 15701 4604 15713 4607
rect 16114 4604 16120 4616
rect 15701 4576 16120 4604
rect 15701 4573 15713 4576
rect 15655 4567 15713 4573
rect 16114 4564 16120 4576
rect 16172 4564 16178 4616
rect 16666 4564 16672 4616
rect 16724 4564 16730 4616
rect 17405 4607 17463 4613
rect 17405 4573 17417 4607
rect 17451 4604 17463 4607
rect 18598 4604 18604 4616
rect 17451 4576 18604 4604
rect 17451 4573 17463 4576
rect 17405 4567 17463 4573
rect 18598 4564 18604 4576
rect 18656 4564 18662 4616
rect 19058 4564 19064 4616
rect 19116 4564 19122 4616
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19352 4604 19380 4632
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 19352 4576 19533 4604
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19705 4607 19763 4613
rect 19705 4573 19717 4607
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 16684 4536 16712 4564
rect 15396 4508 16712 4536
rect 17672 4539 17730 4545
rect 6880 4496 6886 4508
rect 17672 4505 17684 4539
rect 17718 4536 17730 4539
rect 17862 4536 17868 4548
rect 17718 4508 17868 4536
rect 17718 4505 17730 4508
rect 17672 4499 17730 4505
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 19720 4536 19748 4567
rect 19794 4564 19800 4616
rect 19852 4604 19858 4616
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19852 4576 19993 4604
rect 19852 4564 19858 4576
rect 19981 4573 19993 4576
rect 20027 4573 20039 4607
rect 19981 4567 20039 4573
rect 20070 4564 20076 4616
rect 20128 4564 20134 4616
rect 20272 4613 20300 4644
rect 20990 4632 20996 4684
rect 21048 4672 21054 4684
rect 22465 4675 22523 4681
rect 22465 4672 22477 4675
rect 21048 4644 21220 4672
rect 21048 4632 21054 4644
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 20530 4564 20536 4616
rect 20588 4564 20594 4616
rect 20622 4564 20628 4616
rect 20680 4604 20686 4616
rect 20809 4607 20867 4613
rect 20809 4604 20821 4607
rect 20680 4576 20821 4604
rect 20680 4564 20686 4576
rect 20809 4573 20821 4576
rect 20855 4573 20867 4607
rect 20809 4567 20867 4573
rect 20898 4564 20904 4616
rect 20956 4564 20962 4616
rect 21192 4613 21220 4644
rect 22296 4644 22477 4672
rect 22296 4616 22324 4644
rect 22465 4641 22477 4644
rect 22511 4641 22523 4675
rect 22465 4635 22523 4641
rect 21177 4607 21235 4613
rect 21177 4573 21189 4607
rect 21223 4573 21235 4607
rect 21177 4567 21235 4573
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4604 21419 4607
rect 21407 4576 21496 4604
rect 21407 4573 21419 4576
rect 21361 4567 21419 4573
rect 19720 4508 20668 4536
rect 8018 4468 8024 4480
rect 4262 4440 8024 4468
rect 4065 4431 4123 4437
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 9122 4468 9128 4480
rect 8720 4440 9128 4468
rect 8720 4428 8726 4440
rect 9122 4428 9128 4440
rect 9180 4468 9186 4480
rect 10410 4468 10416 4480
rect 9180 4440 10416 4468
rect 9180 4428 9186 4440
rect 10410 4428 10416 4440
rect 10468 4468 10474 4480
rect 11882 4468 11888 4480
rect 10468 4440 11888 4468
rect 10468 4428 10474 4440
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 19794 4428 19800 4480
rect 19852 4428 19858 4480
rect 20254 4428 20260 4480
rect 20312 4428 20318 4480
rect 20640 4477 20668 4508
rect 21468 4477 21496 4576
rect 21634 4564 21640 4616
rect 21692 4564 21698 4616
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4573 21971 4607
rect 21913 4567 21971 4573
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4573 22063 4607
rect 22005 4567 22063 4573
rect 20625 4471 20683 4477
rect 20625 4437 20637 4471
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 21453 4471 21511 4477
rect 21453 4437 21465 4471
rect 21499 4437 21511 4471
rect 21453 4431 21511 4437
rect 21726 4428 21732 4480
rect 21784 4428 21790 4480
rect 21928 4468 21956 4567
rect 22020 4536 22048 4567
rect 22278 4564 22284 4616
rect 22336 4564 22342 4616
rect 22738 4613 22744 4616
rect 22707 4607 22744 4613
rect 22707 4573 22719 4607
rect 22707 4567 22744 4573
rect 22738 4564 22744 4567
rect 22796 4564 22802 4616
rect 25222 4604 25228 4616
rect 23860 4576 25228 4604
rect 23860 4536 23888 4576
rect 25222 4564 25228 4576
rect 25280 4564 25286 4616
rect 22020 4508 23888 4536
rect 23937 4539 23995 4545
rect 23937 4505 23949 4539
rect 23983 4536 23995 4539
rect 24210 4536 24216 4548
rect 23983 4508 24216 4536
rect 23983 4505 23995 4508
rect 23937 4499 23995 4505
rect 24210 4496 24216 4508
rect 24268 4496 24274 4548
rect 22830 4468 22836 4480
rect 21928 4440 22836 4468
rect 22830 4428 22836 4440
rect 22888 4428 22894 4480
rect 22922 4428 22928 4480
rect 22980 4468 22986 4480
rect 23290 4468 23296 4480
rect 22980 4440 23296 4468
rect 22980 4428 22986 4440
rect 23290 4428 23296 4440
rect 23348 4468 23354 4480
rect 23477 4471 23535 4477
rect 23477 4468 23489 4471
rect 23348 4440 23489 4468
rect 23348 4428 23354 4440
rect 23477 4437 23489 4440
rect 23523 4437 23535 4471
rect 23477 4431 23535 4437
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 1504 4236 4353 4264
rect 1504 4205 1532 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 7742 4264 7748 4276
rect 4764 4236 7748 4264
rect 4764 4224 4770 4236
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 8996 4236 14596 4264
rect 8996 4224 9002 4236
rect 1489 4199 1547 4205
rect 1489 4165 1501 4199
rect 1535 4165 1547 4199
rect 10410 4196 10416 4208
rect 1489 4159 1547 4165
rect 9968 4168 10416 4196
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2293 4131 2351 4137
rect 2293 4128 2305 4131
rect 2188 4100 2305 4128
rect 2188 4088 2194 4100
rect 2293 4097 2305 4100
rect 2339 4097 2351 4131
rect 2293 4091 2351 4097
rect 2409 4131 2467 4137
rect 2409 4097 2421 4131
rect 2455 4128 2467 4131
rect 2455 4100 2542 4128
rect 2455 4097 2467 4100
rect 2409 4091 2467 4097
rect 1670 3952 1676 4004
rect 1728 3952 1734 4004
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2514 3992 2542 4100
rect 2590 4088 2596 4140
rect 2648 4088 2654 4140
rect 3326 4088 3332 4140
rect 3384 4088 3390 4140
rect 3510 4137 3516 4140
rect 3467 4131 3516 4137
rect 3467 4097 3479 4131
rect 3513 4097 3516 4131
rect 3467 4091 3516 4097
rect 3510 4088 3516 4091
rect 3568 4088 3574 4140
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4295 4100 4537 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4525 4091 4583 4097
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6730 4128 6736 4140
rect 6236 4100 6736 4128
rect 6236 4088 6242 4100
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 7007 4131 7065 4137
rect 7007 4097 7019 4131
rect 7053 4128 7065 4131
rect 8478 4128 8484 4140
rect 7053 4100 8484 4128
rect 7053 4097 7065 4100
rect 7007 4091 7065 4097
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9306 4088 9312 4140
rect 9364 4088 9370 4140
rect 8110 4020 8116 4072
rect 8168 4020 8174 4072
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4060 8355 4063
rect 8662 4060 8668 4072
rect 8343 4032 8668 4060
rect 8343 4029 8355 4032
rect 8297 4023 8355 4029
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9033 4063 9091 4069
rect 9033 4060 9045 4063
rect 8864 4032 9045 4060
rect 1912 3964 2542 3992
rect 3053 3995 3111 4001
rect 1912 3952 1918 3964
rect 3053 3961 3065 3995
rect 3099 3961 3111 3995
rect 3053 3955 3111 3961
rect 7745 3995 7803 4001
rect 7745 3961 7757 3995
rect 7791 3992 7803 3995
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 7791 3964 8769 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 8757 3961 8769 3964
rect 8803 3961 8815 3995
rect 8757 3955 8815 3961
rect 2130 3884 2136 3936
rect 2188 3884 2194 3936
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 3068 3924 3096 3955
rect 2556 3896 3096 3924
rect 8864 3924 8892 4032
rect 9033 4029 9045 4032
rect 9079 4029 9091 4063
rect 9033 4023 9091 4029
rect 9171 4063 9229 4069
rect 9171 4029 9183 4063
rect 9217 4060 9229 4063
rect 9674 4060 9680 4072
rect 9217 4032 9680 4060
rect 9217 4029 9229 4032
rect 9171 4023 9229 4029
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 9968 4060 9996 4168
rect 10410 4156 10416 4168
rect 10468 4156 10474 4208
rect 10594 4156 10600 4208
rect 10652 4156 10658 4208
rect 10319 4131 10377 4137
rect 10319 4097 10331 4131
rect 10365 4128 10377 4131
rect 10612 4128 10640 4156
rect 10365 4100 10640 4128
rect 10365 4097 10377 4100
rect 10319 4091 10377 4097
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 11514 4128 11520 4140
rect 10744 4100 11520 4128
rect 10744 4088 10750 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11791 4131 11849 4137
rect 11791 4097 11803 4131
rect 11837 4128 11849 4131
rect 12710 4128 12716 4140
rect 11837 4100 12716 4128
rect 11837 4097 11849 4100
rect 11791 4091 11849 4097
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 14568 4137 14596 4236
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 15344 4236 15577 4264
rect 15344 4224 15350 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 17678 4224 17684 4276
rect 17736 4224 17742 4276
rect 18325 4267 18383 4273
rect 18325 4233 18337 4267
rect 18371 4233 18383 4267
rect 18325 4227 18383 4233
rect 15470 4156 15476 4208
rect 15528 4156 15534 4208
rect 18340 4196 18368 4227
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 18874 4264 18880 4276
rect 18564 4236 18880 4264
rect 18564 4224 18570 4236
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 19153 4267 19211 4273
rect 19153 4233 19165 4267
rect 19199 4264 19211 4267
rect 19242 4264 19248 4276
rect 19199 4236 19248 4264
rect 19199 4233 19211 4236
rect 19153 4227 19211 4233
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 20254 4224 20260 4276
rect 20312 4224 20318 4276
rect 20530 4224 20536 4276
rect 20588 4264 20594 4276
rect 21266 4264 21272 4276
rect 20588 4236 21272 4264
rect 20588 4224 20594 4236
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 21453 4267 21511 4273
rect 21453 4233 21465 4267
rect 21499 4264 21511 4267
rect 21634 4264 21640 4276
rect 21499 4236 21640 4264
rect 21499 4233 21511 4236
rect 21453 4227 21511 4233
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 22278 4224 22284 4276
rect 22336 4264 22342 4276
rect 23198 4264 23204 4276
rect 22336 4236 23204 4264
rect 22336 4224 22342 4236
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 19613 4199 19671 4205
rect 19613 4196 19625 4199
rect 18340 4168 19625 4196
rect 19613 4165 19625 4168
rect 19659 4165 19671 4199
rect 20272 4196 20300 4224
rect 24305 4199 24363 4205
rect 20272 4168 24072 4196
rect 19613 4159 19671 4165
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4128 14611 4131
rect 14734 4128 14740 4140
rect 14599 4100 14740 4128
rect 14599 4097 14611 4100
rect 14553 4091 14611 4097
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 14827 4131 14885 4137
rect 14827 4097 14839 4131
rect 14873 4128 14885 4131
rect 15488 4128 15516 4156
rect 24044 4140 24072 4168
rect 24305 4165 24317 4199
rect 24351 4196 24363 4199
rect 24578 4196 24584 4208
rect 24351 4168 24584 4196
rect 24351 4165 24363 4168
rect 24305 4159 24363 4165
rect 24578 4156 24584 4168
rect 24636 4156 24642 4208
rect 14873 4100 15516 4128
rect 14873 4097 14885 4100
rect 14827 4091 14885 4097
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 18322 4088 18328 4140
rect 18380 4088 18386 4140
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4128 18567 4131
rect 18690 4128 18696 4140
rect 18555 4100 18696 4128
rect 18555 4097 18567 4100
rect 18509 4091 18567 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 18966 4128 18972 4140
rect 18831 4100 18972 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19061 4131 19119 4137
rect 19061 4097 19073 4131
rect 19107 4128 19119 4131
rect 19337 4131 19395 4137
rect 19107 4100 19196 4128
rect 19107 4097 19119 4100
rect 19061 4091 19119 4097
rect 9732 4032 9996 4060
rect 9732 4020 9738 4032
rect 10042 4020 10048 4072
rect 10100 4020 10106 4072
rect 9876 3964 10180 3992
rect 9674 3924 9680 3936
rect 8864 3896 9680 3924
rect 2556 3884 2562 3896
rect 9674 3884 9680 3896
rect 9732 3924 9738 3936
rect 9876 3924 9904 3964
rect 10152 3936 10180 3964
rect 9732 3896 9904 3924
rect 9732 3884 9738 3896
rect 9950 3884 9956 3936
rect 10008 3884 10014 3936
rect 10134 3884 10140 3936
rect 10192 3884 10198 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 11057 3927 11115 3933
rect 11057 3924 11069 3927
rect 10376 3896 11069 3924
rect 10376 3884 10382 3896
rect 11057 3893 11069 3896
rect 11103 3893 11115 3927
rect 11057 3887 11115 3893
rect 12526 3884 12532 3936
rect 12584 3884 12590 3936
rect 17880 3924 17908 4088
rect 18340 4060 18368 4088
rect 19168 4060 19196 4100
rect 19337 4097 19349 4131
rect 19383 4128 19395 4131
rect 19426 4128 19432 4140
rect 19383 4100 19432 4128
rect 19383 4097 19395 4100
rect 19337 4091 19395 4097
rect 19426 4088 19432 4100
rect 19484 4088 19490 4140
rect 20346 4137 20352 4140
rect 20340 4128 20352 4137
rect 20307 4100 20352 4128
rect 20340 4091 20352 4100
rect 20346 4088 20352 4091
rect 20404 4088 20410 4140
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4128 22431 4131
rect 22462 4128 22468 4140
rect 22419 4100 22468 4128
rect 22419 4097 22431 4100
rect 22373 4091 22431 4097
rect 22462 4088 22468 4100
rect 22520 4088 22526 4140
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 18340 4032 19196 4060
rect 20070 4020 20076 4072
rect 20128 4020 20134 4072
rect 22005 4063 22063 4069
rect 22005 4029 22017 4063
rect 22051 4060 22063 4063
rect 22094 4060 22100 4072
rect 22051 4032 22100 4060
rect 22051 4029 22063 4032
rect 22005 4023 22063 4029
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 22664 4060 22692 4091
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 23017 4131 23075 4137
rect 23017 4128 23029 4131
rect 22796 4100 23029 4128
rect 22796 4088 22802 4100
rect 23017 4097 23029 4100
rect 23063 4097 23075 4131
rect 23017 4091 23075 4097
rect 23382 4088 23388 4140
rect 23440 4128 23446 4140
rect 23440 4100 23980 4128
rect 23440 4088 23446 4100
rect 22244 4032 22692 4060
rect 23845 4063 23903 4069
rect 22244 4020 22250 4032
rect 23845 4029 23857 4063
rect 23891 4029 23903 4063
rect 23952 4060 23980 4100
rect 24026 4088 24032 4140
rect 24084 4088 24090 4140
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4097 24547 4131
rect 24489 4091 24547 4097
rect 24504 4060 24532 4091
rect 23952 4032 24532 4060
rect 23845 4023 23903 4029
rect 18966 3952 18972 4004
rect 19024 3992 19030 4004
rect 19024 3964 20116 3992
rect 19024 3952 19030 3964
rect 18601 3927 18659 3933
rect 18601 3924 18613 3927
rect 17880 3896 18613 3924
rect 18601 3893 18613 3896
rect 18647 3893 18659 3927
rect 18601 3887 18659 3893
rect 18877 3927 18935 3933
rect 18877 3893 18889 3927
rect 18923 3924 18935 3927
rect 19150 3924 19156 3936
rect 18923 3896 19156 3924
rect 18923 3893 18935 3896
rect 18877 3887 18935 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19705 3927 19763 3933
rect 19705 3924 19717 3927
rect 19300 3896 19717 3924
rect 19300 3884 19306 3896
rect 19705 3893 19717 3896
rect 19751 3893 19763 3927
rect 20088 3924 20116 3964
rect 22646 3952 22652 4004
rect 22704 3952 22710 4004
rect 23860 3992 23888 4023
rect 24302 3992 24308 4004
rect 23860 3964 24308 3992
rect 24302 3952 24308 3964
rect 24360 3952 24366 4004
rect 20438 3924 20444 3936
rect 20088 3896 20444 3924
rect 19705 3887 19763 3893
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 21450 3924 21456 3936
rect 20864 3896 21456 3924
rect 20864 3884 20870 3896
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 22278 3884 22284 3936
rect 22336 3924 22342 3936
rect 23934 3924 23940 3936
rect 22336 3896 23940 3924
rect 22336 3884 22342 3896
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 1762 3680 1768 3732
rect 1820 3680 1826 3732
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 5350 3720 5356 3732
rect 2188 3692 5356 3720
rect 2188 3680 2194 3692
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 9398 3720 9404 3732
rect 7208 3692 9404 3720
rect 1394 3612 1400 3664
rect 1452 3652 1458 3664
rect 2409 3655 2467 3661
rect 2409 3652 2421 3655
rect 1452 3624 2421 3652
rect 1452 3612 1458 3624
rect 2409 3621 2421 3624
rect 2455 3621 2467 3655
rect 2409 3615 2467 3621
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 2832 3624 2881 3652
rect 2832 3612 2838 3624
rect 2869 3621 2881 3624
rect 2915 3621 2927 3655
rect 2869 3615 2927 3621
rect 5074 3612 5080 3664
rect 5132 3612 5138 3664
rect 7208 3661 7236 3692
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9548 3692 10916 3720
rect 9548 3680 9554 3692
rect 7193 3655 7251 3661
rect 7193 3621 7205 3655
rect 7239 3621 7251 3655
rect 7193 3615 7251 3621
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 8527 3624 9536 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 3694 3584 3700 3596
rect 1688 3556 3700 3584
rect 1688 3525 1716 3556
rect 3694 3544 3700 3556
rect 3752 3544 3758 3596
rect 5092 3584 5120 3612
rect 4816 3556 5120 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1780 3488 2360 3516
rect 14 3408 20 3460
rect 72 3448 78 3460
rect 1780 3448 1808 3488
rect 72 3420 1808 3448
rect 72 3408 78 3420
rect 2222 3408 2228 3460
rect 2280 3408 2286 3460
rect 2332 3448 2360 3488
rect 2682 3476 2688 3528
rect 2740 3476 2746 3528
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 2832 3488 4568 3516
rect 2832 3476 2838 3488
rect 4540 3448 4568 3488
rect 4614 3476 4620 3528
rect 4672 3516 4678 3528
rect 4816 3525 4844 3556
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 7469 3587 7527 3593
rect 7469 3584 7481 3587
rect 6788 3556 7481 3584
rect 6788 3544 6794 3556
rect 7469 3553 7481 3556
rect 7515 3553 7527 3587
rect 9508 3584 9536 3624
rect 9674 3612 9680 3664
rect 9732 3612 9738 3664
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9508 3556 9597 3584
rect 7469 3547 7527 3553
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9692 3584 9720 3612
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9692 3556 9873 3584
rect 9585 3547 9643 3553
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 9861 3547 9919 3553
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4672 3488 4813 3516
rect 4672 3476 4678 3488
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5351 3519 5409 3525
rect 5351 3485 5363 3519
rect 5397 3516 5409 3519
rect 7282 3516 7288 3528
rect 5397 3488 7288 3516
rect 5397 3485 5409 3488
rect 5351 3479 5409 3485
rect 5092 3448 5120 3479
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7484 3516 7512 3547
rect 9950 3544 9956 3596
rect 10008 3593 10014 3596
rect 10008 3587 10036 3593
rect 10024 3553 10036 3587
rect 10008 3547 10036 3553
rect 10008 3544 10014 3547
rect 7650 3516 7656 3528
rect 7484 3488 7656 3516
rect 7377 3479 7435 3485
rect 5994 3448 6000 3460
rect 2332 3420 2774 3448
rect 4540 3420 5028 3448
rect 5092 3420 6000 3448
rect 2038 3340 2044 3392
rect 2096 3380 2102 3392
rect 2590 3380 2596 3392
rect 2096 3352 2596 3380
rect 2096 3340 2102 3352
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 2746 3380 2774 3420
rect 4522 3380 4528 3392
rect 2746 3352 4528 3380
rect 4522 3340 4528 3352
rect 4580 3340 4586 3392
rect 4890 3340 4896 3392
rect 4948 3340 4954 3392
rect 5000 3380 5028 3420
rect 5994 3408 6000 3420
rect 6052 3408 6058 3460
rect 6917 3451 6975 3457
rect 6917 3417 6929 3451
rect 6963 3448 6975 3451
rect 7392 3448 7420 3479
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 7743 3519 7801 3525
rect 7743 3485 7755 3519
rect 7789 3516 7801 3519
rect 7834 3516 7840 3528
rect 7789 3488 7840 3516
rect 7789 3485 7801 3488
rect 7743 3479 7801 3485
rect 7834 3476 7840 3488
rect 7892 3476 7898 3528
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8168 3488 8953 3516
rect 8168 3476 8174 3488
rect 8941 3485 8953 3488
rect 8987 3516 8999 3519
rect 9030 3516 9036 3528
rect 8987 3488 9036 3516
rect 8987 3485 8999 3488
rect 8941 3479 8999 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 8202 3448 8208 3460
rect 6963 3420 8208 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 5902 3380 5908 3392
rect 5000 3352 5908 3380
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6086 3340 6092 3392
rect 6144 3340 6150 3392
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 10781 3383 10839 3389
rect 10781 3380 10793 3383
rect 7340 3352 10793 3380
rect 7340 3340 7346 3352
rect 10781 3349 10793 3352
rect 10827 3349 10839 3383
rect 10888 3380 10916 3692
rect 13354 3680 13360 3732
rect 13412 3680 13418 3732
rect 13906 3680 13912 3732
rect 13964 3720 13970 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 13964 3692 15117 3720
rect 13964 3680 13970 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15105 3683 15163 3689
rect 17586 3680 17592 3732
rect 17644 3720 17650 3732
rect 17644 3692 18092 3720
rect 17644 3680 17650 3692
rect 18064 3652 18092 3692
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19978 3720 19984 3732
rect 18840 3692 19984 3720
rect 18840 3680 18846 3692
rect 18509 3655 18567 3661
rect 18064 3624 18451 3652
rect 12526 3544 12532 3596
rect 12584 3544 12590 3596
rect 18138 3584 18144 3596
rect 14752 3556 18144 3584
rect 13722 3516 13728 3528
rect 12084 3488 13728 3516
rect 12084 3457 12112 3488
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 12069 3451 12127 3457
rect 12069 3417 12081 3451
rect 12115 3417 12127 3451
rect 12069 3411 12127 3417
rect 12250 3408 12256 3460
rect 12308 3448 12314 3460
rect 12345 3451 12403 3457
rect 12345 3448 12357 3451
rect 12308 3420 12357 3448
rect 12308 3408 12314 3420
rect 12345 3417 12357 3420
rect 12391 3417 12403 3451
rect 12345 3411 12403 3417
rect 12434 3408 12440 3460
rect 12492 3408 12498 3460
rect 12526 3408 12532 3460
rect 12584 3448 12590 3460
rect 12805 3451 12863 3457
rect 12805 3448 12817 3451
rect 12584 3420 12817 3448
rect 12584 3408 12590 3420
rect 12805 3417 12817 3420
rect 12851 3417 12863 3451
rect 12805 3411 12863 3417
rect 12894 3408 12900 3460
rect 12952 3448 12958 3460
rect 14108 3448 14136 3479
rect 14366 3476 14372 3528
rect 14424 3476 14430 3528
rect 14752 3448 14780 3556
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18049 3519 18107 3525
rect 17954 3452 17960 3504
rect 18012 3452 18018 3504
rect 18049 3485 18061 3519
rect 18095 3486 18107 3519
rect 18325 3519 18383 3525
rect 18095 3485 18184 3486
rect 18049 3479 18184 3485
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 18423 3516 18451 3624
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 19150 3652 19156 3664
rect 18555 3624 19156 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 19260 3593 19288 3692
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 20622 3680 20628 3732
rect 20680 3680 20686 3732
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23256 3692 23949 3720
rect 23256 3680 23262 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 23937 3683 23995 3689
rect 23106 3612 23112 3664
rect 23164 3652 23170 3664
rect 23164 3624 23244 3652
rect 23164 3612 23170 3624
rect 19245 3587 19303 3593
rect 19245 3553 19257 3587
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 20898 3544 20904 3596
rect 20956 3584 20962 3596
rect 23216 3593 23244 3624
rect 21269 3587 21327 3593
rect 21269 3584 21281 3587
rect 20956 3556 21281 3584
rect 20956 3544 20962 3556
rect 21269 3553 21281 3556
rect 21315 3553 21327 3587
rect 21269 3547 21327 3553
rect 23201 3587 23259 3593
rect 23201 3553 23213 3587
rect 23247 3553 23259 3587
rect 23201 3547 23259 3553
rect 18371 3488 18451 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 18064 3458 18184 3479
rect 18782 3476 18788 3528
rect 18840 3476 18846 3528
rect 19058 3476 19064 3528
rect 19116 3476 19122 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20772 3488 20821 3516
rect 20772 3476 20778 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 21450 3476 21456 3528
rect 21508 3516 21514 3528
rect 21543 3519 21601 3525
rect 21543 3516 21555 3519
rect 21508 3488 21555 3516
rect 21508 3476 21514 3488
rect 21543 3485 21555 3488
rect 21589 3485 21601 3519
rect 21543 3479 21601 3485
rect 22278 3476 22284 3528
rect 22336 3516 22342 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22336 3488 22661 3516
rect 22336 3476 22342 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 23164 3488 23765 3516
rect 23164 3476 23170 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 12952 3420 14780 3448
rect 12952 3408 12958 3420
rect 13173 3383 13231 3389
rect 13173 3380 13185 3383
rect 10888 3352 13185 3380
rect 10781 3343 10839 3349
rect 13173 3349 13185 3352
rect 13219 3349 13231 3383
rect 13173 3343 13231 3349
rect 13538 3340 13544 3392
rect 13596 3340 13602 3392
rect 17770 3340 17776 3392
rect 17828 3340 17834 3392
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18156 3380 18184 3458
rect 19334 3448 19340 3460
rect 18248 3420 19340 3448
rect 18248 3389 18276 3420
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 19518 3457 19524 3460
rect 19512 3411 19524 3457
rect 19576 3448 19582 3460
rect 19576 3420 19612 3448
rect 19518 3408 19524 3411
rect 19576 3408 19582 3420
rect 20990 3408 20996 3460
rect 21048 3448 21054 3460
rect 24486 3448 24492 3460
rect 21048 3420 23336 3448
rect 21048 3408 21054 3420
rect 18104 3352 18184 3380
rect 18233 3383 18291 3389
rect 18104 3340 18110 3352
rect 18233 3349 18245 3383
rect 18279 3349 18291 3383
rect 18233 3343 18291 3349
rect 18598 3340 18604 3392
rect 18656 3340 18662 3392
rect 18690 3340 18696 3392
rect 18748 3380 18754 3392
rect 18877 3383 18935 3389
rect 18877 3380 18889 3383
rect 18748 3352 18889 3380
rect 18748 3340 18754 3352
rect 18877 3349 18889 3352
rect 18923 3349 18935 3383
rect 18877 3343 18935 3349
rect 19702 3340 19708 3392
rect 19760 3380 19766 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 19760 3352 20913 3380
rect 19760 3340 19766 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 22094 3340 22100 3392
rect 22152 3380 22158 3392
rect 22281 3383 22339 3389
rect 22281 3380 22293 3383
rect 22152 3352 22293 3380
rect 22152 3340 22158 3352
rect 22281 3349 22293 3352
rect 22327 3349 22339 3383
rect 23308 3380 23336 3420
rect 23584 3420 24492 3448
rect 23584 3380 23612 3420
rect 24486 3408 24492 3420
rect 24544 3408 24550 3460
rect 23308 3352 23612 3380
rect 22281 3343 22339 3349
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 1578 3136 1584 3188
rect 1636 3136 1642 3188
rect 2222 3136 2228 3188
rect 2280 3176 2286 3188
rect 2593 3179 2651 3185
rect 2593 3176 2605 3179
rect 2280 3148 2605 3176
rect 2280 3136 2286 3148
rect 2593 3145 2605 3148
rect 2639 3145 2651 3179
rect 2593 3139 2651 3145
rect 3326 3136 3332 3188
rect 3384 3136 3390 3188
rect 4522 3136 4528 3188
rect 4580 3136 4586 3188
rect 7282 3176 7288 3188
rect 6472 3148 7288 3176
rect 1026 3068 1032 3120
rect 1084 3108 1090 3120
rect 2314 3108 2320 3120
rect 1084 3080 2084 3108
rect 1084 3068 1090 3080
rect 2056 3049 2084 3080
rect 2240 3080 2320 3108
rect 2240 3049 2268 3080
rect 2314 3068 2320 3080
rect 2372 3068 2378 3120
rect 6472 3108 6500 3148
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7837 3179 7895 3185
rect 7837 3176 7849 3179
rect 7524 3148 7849 3176
rect 7524 3136 7530 3148
rect 7837 3145 7849 3148
rect 7883 3145 7895 3179
rect 7837 3139 7895 3145
rect 9125 3179 9183 3185
rect 9125 3145 9137 3179
rect 9171 3176 9183 3179
rect 9306 3176 9312 3188
rect 9171 3148 9312 3176
rect 9171 3145 9183 3148
rect 9125 3139 9183 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9953 3179 10011 3185
rect 9953 3145 9965 3179
rect 9999 3176 10011 3179
rect 11790 3176 11796 3188
rect 9999 3148 11796 3176
rect 9999 3145 10011 3148
rect 9953 3139 10011 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12066 3136 12072 3188
rect 12124 3136 12130 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 12492 3148 13185 3176
rect 12492 3136 12498 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 14366 3136 14372 3188
rect 14424 3136 14430 3188
rect 17129 3179 17187 3185
rect 17129 3145 17141 3179
rect 17175 3176 17187 3179
rect 17678 3176 17684 3188
rect 17175 3148 17684 3176
rect 17175 3145 17187 3148
rect 17129 3139 17187 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 17788 3148 18061 3176
rect 2516 3080 6500 3108
rect 2516 3049 2544 3080
rect 6546 3068 6552 3120
rect 6604 3068 6610 3120
rect 7653 3111 7711 3117
rect 7653 3108 7665 3111
rect 6654 3080 7665 3108
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3009 1547 3043
rect 1489 3003 1547 3009
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3009 2099 3043
rect 2041 3003 2099 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2501 3043 2559 3049
rect 2501 3009 2513 3043
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 1504 2972 1532 3003
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 1504 2944 2728 2972
rect 2700 2904 2728 2944
rect 3050 2932 3056 2984
rect 3108 2972 3114 2984
rect 3252 2972 3280 3003
rect 3326 3000 3332 3052
rect 3384 3040 3390 3052
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 3384 3012 4445 3040
rect 3384 3000 3390 3012
rect 4433 3009 4445 3012
rect 4479 3040 4491 3043
rect 6654 3040 6682 3080
rect 7653 3077 7665 3080
rect 7699 3077 7711 3111
rect 7653 3071 7711 3077
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 9582 3108 9588 3120
rect 7800 3080 9588 3108
rect 7800 3068 7806 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 10134 3068 10140 3120
rect 10192 3108 10198 3120
rect 10229 3111 10287 3117
rect 10229 3108 10241 3111
rect 10192 3080 10241 3108
rect 10192 3068 10198 3080
rect 10229 3077 10241 3080
rect 10275 3077 10287 3111
rect 10229 3071 10287 3077
rect 10318 3068 10324 3120
rect 10376 3068 10382 3120
rect 10410 3068 10416 3120
rect 10468 3108 10474 3120
rect 10468 3080 11008 3108
rect 10468 3068 10474 3080
rect 4479 3012 6682 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 6822 3000 6828 3052
rect 6880 3000 6886 3052
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7064 3012 7297 3040
rect 7064 3000 7070 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7285 3003 7343 3009
rect 7668 3012 8125 3040
rect 7668 2984 7696 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8387 3043 8445 3049
rect 8387 3009 8399 3043
rect 8433 3040 8445 3043
rect 8433 3012 9260 3040
rect 8433 3009 8445 3012
rect 8387 3003 8445 3009
rect 4062 2972 4068 2984
rect 3108 2944 4068 2972
rect 3108 2932 3114 2944
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 6144 2944 6394 2972
rect 6144 2932 6150 2944
rect 7650 2932 7656 2984
rect 7708 2932 7714 2984
rect 3418 2904 3424 2916
rect 2700 2876 3424 2904
rect 3418 2864 3424 2876
rect 3476 2864 3482 2916
rect 2317 2839 2375 2845
rect 2317 2805 2329 2839
rect 2363 2836 2375 2839
rect 3142 2836 3148 2848
rect 2363 2808 3148 2836
rect 2363 2805 2375 2808
rect 2317 2799 2375 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 8128 2836 8156 3003
rect 9232 2904 9260 3012
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9677 3043 9735 3049
rect 9677 3040 9689 3043
rect 9364 3012 9689 3040
rect 9364 3000 9370 3012
rect 9677 3009 9689 3012
rect 9723 3009 9735 3043
rect 9677 3003 9735 3009
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 10428 3040 10456 3068
rect 10100 3012 10456 3040
rect 10100 3000 10106 3012
rect 10502 3000 10508 3052
rect 10560 3040 10566 3052
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10560 3012 10701 3040
rect 10560 3000 10566 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10980 3040 11008 3080
rect 11054 3068 11060 3120
rect 11112 3068 11118 3120
rect 11514 3068 11520 3120
rect 11572 3068 11578 3120
rect 10980 3012 11284 3040
rect 10689 3003 10747 3009
rect 10778 2932 10784 2984
rect 10836 2932 10842 2984
rect 11256 2913 11284 3012
rect 11532 2972 11560 3068
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 11808 3040 11836 3136
rect 12084 3049 12112 3136
rect 12158 3068 12164 3120
rect 12216 3068 12222 3120
rect 11747 3012 11836 3040
rect 12069 3043 12127 3049
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12176 3040 12204 3068
rect 12435 3043 12493 3049
rect 12435 3040 12447 3043
rect 12176 3012 12447 3040
rect 12069 3003 12127 3009
rect 12435 3009 12447 3012
rect 12481 3040 12493 3043
rect 14384 3040 14412 3136
rect 16758 3068 16764 3120
rect 16816 3108 16822 3120
rect 17788 3108 17816 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 18785 3179 18843 3185
rect 18380 3148 18460 3176
rect 18380 3136 18386 3148
rect 16816 3080 17816 3108
rect 16816 3068 16822 3080
rect 18432 3064 18460 3148
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 19058 3176 19064 3188
rect 18831 3148 19064 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19518 3136 19524 3188
rect 19576 3136 19582 3188
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 20956 3148 21312 3176
rect 20956 3136 20962 3148
rect 18509 3067 18567 3073
rect 18966 3068 18972 3120
rect 19024 3108 19030 3120
rect 19536 3108 19564 3136
rect 20990 3108 20996 3120
rect 19024 3080 19564 3108
rect 19720 3080 20996 3108
rect 19024 3068 19030 3080
rect 18509 3064 18521 3067
rect 12481 3012 14412 3040
rect 16945 3043 17003 3049
rect 12481 3009 12493 3012
rect 12435 3003 12493 3009
rect 16945 3009 16957 3043
rect 16991 3009 17003 3043
rect 16945 3003 17003 3009
rect 12158 2972 12164 2984
rect 11532 2944 12164 2972
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 16960 2972 16988 3003
rect 17218 3000 17224 3052
rect 17276 3000 17282 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 17862 3040 17868 3052
rect 17543 3012 17868 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 17954 3000 17960 3052
rect 18012 3000 18018 3052
rect 18230 3000 18236 3052
rect 18288 3000 18294 3052
rect 18432 3036 18521 3064
rect 18509 3033 18521 3036
rect 18555 3033 18567 3067
rect 18509 3027 18567 3033
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19720 3049 19748 3080
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 21284 3108 21312 3148
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 21416 3148 23397 3176
rect 21416 3136 21422 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 21284 3080 22416 3108
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18932 3012 19257 3040
rect 18932 3000 18938 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 19794 3000 19800 3052
rect 19852 3040 19858 3052
rect 20809 3043 20867 3049
rect 19852 3012 20760 3040
rect 19852 3000 19858 3012
rect 16960 2944 17448 2972
rect 11241 2907 11299 2913
rect 9232 2876 9674 2904
rect 8938 2836 8944 2848
rect 8128 2808 8944 2836
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9272 2808 9505 2836
rect 9272 2796 9278 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9646 2836 9674 2876
rect 11241 2873 11253 2907
rect 11287 2873 11299 2907
rect 11241 2867 11299 2873
rect 11532 2876 12018 2904
rect 9950 2836 9956 2848
rect 9646 2808 9956 2836
rect 9493 2799 9551 2805
rect 9950 2796 9956 2808
rect 10008 2796 10014 2848
rect 11532 2845 11560 2876
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 11882 2796 11888 2848
rect 11940 2796 11946 2848
rect 11990 2836 12018 2876
rect 13814 2836 13820 2848
rect 11990 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 17420 2845 17448 2944
rect 17586 2932 17592 2984
rect 17644 2972 17650 2984
rect 19610 2972 19616 2984
rect 17644 2944 19616 2972
rect 17644 2932 17650 2944
rect 17696 2913 17724 2944
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 19886 2932 19892 2984
rect 19944 2972 19950 2984
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 19944 2944 19993 2972
rect 19944 2932 19950 2944
rect 19981 2941 19993 2944
rect 20027 2941 20039 2975
rect 20732 2972 20760 3012
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 21174 3040 21180 3052
rect 20855 3012 21180 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 21174 3000 21180 3012
rect 21232 3000 21238 3052
rect 22388 3049 22416 3080
rect 21913 3043 21971 3049
rect 21913 3040 21925 3043
rect 21376 3012 21925 3040
rect 21376 2972 21404 3012
rect 21913 3009 21925 3012
rect 21959 3009 21971 3043
rect 21913 3003 21971 3009
rect 22373 3043 22431 3049
rect 22373 3009 22385 3043
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 22647 3043 22705 3049
rect 22647 3009 22659 3043
rect 22693 3040 22705 3043
rect 23014 3040 23020 3052
rect 22693 3012 23020 3040
rect 22693 3009 22705 3012
rect 22647 3003 22705 3009
rect 23014 3000 23020 3012
rect 23072 3000 23078 3052
rect 23400 3040 23428 3139
rect 24026 3068 24032 3120
rect 24084 3108 24090 3120
rect 24305 3111 24363 3117
rect 24305 3108 24317 3111
rect 24084 3080 24317 3108
rect 24084 3068 24090 3080
rect 24305 3077 24317 3080
rect 24351 3077 24363 3111
rect 24305 3071 24363 3077
rect 23753 3043 23811 3049
rect 23753 3040 23765 3043
rect 23400 3012 23765 3040
rect 23753 3009 23765 3012
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 23842 3000 23848 3052
rect 23900 3040 23906 3052
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 23900 3012 23949 3040
rect 23900 3000 23906 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 20732 2944 21404 2972
rect 21453 2975 21511 2981
rect 19981 2935 20039 2941
rect 21453 2941 21465 2975
rect 21499 2972 21511 2975
rect 21542 2972 21548 2984
rect 21499 2944 21548 2972
rect 21499 2941 21511 2944
rect 21453 2935 21511 2941
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 17681 2907 17739 2913
rect 17681 2873 17693 2907
rect 17727 2873 17739 2907
rect 17681 2867 17739 2873
rect 17773 2907 17831 2913
rect 17773 2873 17785 2907
rect 17819 2873 17831 2907
rect 17773 2867 17831 2873
rect 18262 2876 18644 2904
rect 17405 2839 17463 2845
rect 17405 2805 17417 2839
rect 17451 2836 17463 2839
rect 17494 2836 17500 2848
rect 17451 2808 17500 2836
rect 17451 2805 17463 2808
rect 17405 2799 17463 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 17788 2836 17816 2867
rect 18262 2836 18290 2876
rect 17788 2808 18290 2836
rect 18322 2796 18328 2848
rect 18380 2796 18386 2848
rect 18616 2836 18644 2876
rect 18690 2864 18696 2916
rect 18748 2904 18754 2916
rect 20714 2904 20720 2916
rect 18748 2876 20720 2904
rect 18748 2864 18754 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 20806 2864 20812 2916
rect 20864 2904 20870 2916
rect 23937 2907 23995 2913
rect 23937 2904 23949 2907
rect 20864 2876 22508 2904
rect 20864 2864 20870 2876
rect 18966 2836 18972 2848
rect 18616 2808 18972 2836
rect 18966 2796 18972 2808
rect 19024 2796 19030 2848
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19337 2839 19395 2845
rect 19337 2836 19349 2839
rect 19208 2808 19349 2836
rect 19208 2796 19214 2808
rect 19337 2805 19349 2808
rect 19383 2805 19395 2839
rect 19337 2799 19395 2805
rect 19978 2796 19984 2848
rect 20036 2836 20042 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 20036 2808 22017 2836
rect 20036 2796 20042 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22480 2836 22508 2876
rect 23032 2876 23949 2904
rect 23032 2836 23060 2876
rect 23937 2873 23949 2876
rect 23983 2873 23995 2907
rect 23937 2867 23995 2873
rect 22480 2808 23060 2836
rect 22005 2799 22063 2805
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2130 2632 2136 2644
rect 1995 2604 2136 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2130 2592 2136 2604
rect 2188 2592 2194 2644
rect 2332 2604 2912 2632
rect 1673 2567 1731 2573
rect 1673 2533 1685 2567
rect 1719 2564 1731 2567
rect 2332 2564 2360 2604
rect 1719 2536 2360 2564
rect 1719 2533 1731 2536
rect 1673 2527 1731 2533
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 2225 2499 2283 2505
rect 2225 2496 2237 2499
rect 1360 2468 2237 2496
rect 1360 2456 1366 2468
rect 2225 2465 2237 2468
rect 2271 2465 2283 2499
rect 2884 2496 2912 2604
rect 2958 2592 2964 2644
rect 3016 2632 3022 2644
rect 3237 2635 3295 2641
rect 3237 2632 3249 2635
rect 3016 2604 3249 2632
rect 3016 2592 3022 2604
rect 3237 2601 3249 2604
rect 3283 2601 3295 2635
rect 3237 2595 3295 2601
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 5626 2632 5632 2644
rect 4663 2604 5632 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 5810 2592 5816 2644
rect 5868 2592 5874 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 6914 2632 6920 2644
rect 6871 2604 6920 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7926 2632 7932 2644
rect 7340 2604 7932 2632
rect 7340 2592 7346 2604
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8036 2604 8800 2632
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2564 4031 2567
rect 5074 2564 5080 2576
rect 4019 2536 5080 2564
rect 4019 2533 4031 2536
rect 3973 2527 4031 2533
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5828 2496 5856 2592
rect 8036 2576 8064 2604
rect 8018 2524 8024 2576
rect 8076 2524 8082 2576
rect 8772 2564 8800 2604
rect 9490 2592 9496 2644
rect 9548 2592 9554 2644
rect 9968 2604 10548 2632
rect 9968 2564 9996 2604
rect 8772 2536 9996 2564
rect 10520 2564 10548 2604
rect 10778 2592 10784 2644
rect 10836 2632 10842 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10836 2604 10885 2632
rect 10836 2592 10842 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 10980 2604 12020 2632
rect 10980 2564 11008 2604
rect 10520 2536 11008 2564
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11885 2567 11943 2573
rect 11885 2564 11897 2567
rect 11112 2536 11897 2564
rect 11112 2524 11118 2536
rect 11885 2533 11897 2536
rect 11931 2533 11943 2567
rect 11992 2564 12020 2604
rect 12250 2592 12256 2644
rect 12308 2632 12314 2644
rect 12308 2604 16574 2632
rect 12308 2592 12314 2604
rect 12526 2564 12532 2576
rect 11992 2536 12532 2564
rect 11885 2527 11943 2533
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 7742 2496 7748 2508
rect 2884 2468 5856 2496
rect 7392 2468 7748 2496
rect 2225 2459 2283 2465
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1596 2400 1777 2428
rect 474 2320 480 2372
rect 532 2360 538 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 532 2332 1501 2360
rect 532 2320 538 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 1596 2292 1624 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 2499 2431 2557 2437
rect 2499 2397 2511 2431
rect 2545 2428 2557 2431
rect 2590 2428 2596 2440
rect 2545 2400 2596 2428
rect 2545 2397 2557 2400
rect 2499 2391 2557 2397
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2746 2400 3801 2428
rect 2746 2372 2774 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 4430 2388 4436 2440
rect 4488 2388 4494 2440
rect 4890 2388 4896 2440
rect 4948 2388 4954 2440
rect 5718 2388 5724 2440
rect 5776 2388 5782 2440
rect 5810 2388 5816 2440
rect 5868 2388 5874 2440
rect 6087 2431 6145 2437
rect 6087 2397 6099 2431
rect 6133 2428 6145 2431
rect 6730 2428 6736 2440
rect 6133 2400 6736 2428
rect 6133 2397 6145 2400
rect 6087 2391 6145 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7392 2437 7420 2468
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 8628 2468 9076 2496
rect 8628 2456 8634 2468
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7650 2388 7656 2440
rect 7708 2388 7714 2440
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8402 2400 8493 2428
rect 2682 2320 2688 2372
rect 2740 2332 2774 2372
rect 7852 2360 7880 2388
rect 8402 2360 8430 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 8754 2388 8760 2440
rect 8812 2388 8818 2440
rect 9048 2360 9076 2468
rect 10686 2456 10692 2508
rect 10744 2456 10750 2508
rect 11238 2456 11244 2508
rect 11296 2496 11302 2508
rect 11296 2468 11836 2496
rect 11296 2456 11302 2468
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9490 2428 9496 2440
rect 9355 2400 9496 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10103 2431 10161 2437
rect 10103 2428 10115 2431
rect 9968 2400 10115 2428
rect 9968 2360 9996 2400
rect 10103 2397 10115 2400
rect 10149 2397 10161 2431
rect 10103 2391 10161 2397
rect 10704 2360 10732 2456
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11808 2437 11836 2468
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 14148 2468 15148 2496
rect 14148 2456 14154 2468
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11204 2400 11529 2428
rect 11204 2388 11210 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11793 2431 11851 2437
rect 11793 2397 11805 2431
rect 11839 2397 11851 2431
rect 11793 2391 11851 2397
rect 12066 2388 12072 2440
rect 12124 2388 12130 2440
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12345 2431 12403 2437
rect 12345 2428 12357 2431
rect 12216 2400 12357 2428
rect 12216 2388 12222 2400
rect 12345 2397 12357 2400
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12894 2388 12900 2440
rect 12952 2388 12958 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 14826 2388 14832 2440
rect 14884 2388 14890 2440
rect 15120 2437 15148 2468
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2428 15439 2431
rect 15562 2428 15568 2440
rect 15427 2400 15568 2428
rect 15427 2397 15439 2400
rect 15381 2391 15439 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15654 2388 15660 2440
rect 15712 2388 15718 2440
rect 16390 2388 16396 2440
rect 16448 2388 16454 2440
rect 16546 2360 16574 2604
rect 17034 2592 17040 2644
rect 17092 2632 17098 2644
rect 17681 2635 17739 2641
rect 17681 2632 17693 2635
rect 17092 2604 17693 2632
rect 17092 2592 17098 2604
rect 17681 2601 17693 2604
rect 17727 2601 17739 2635
rect 17681 2595 17739 2601
rect 17862 2592 17868 2644
rect 17920 2632 17926 2644
rect 23474 2632 23480 2644
rect 17920 2604 23480 2632
rect 17920 2592 17926 2604
rect 23474 2592 23480 2604
rect 23532 2592 23538 2644
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 24213 2635 24271 2641
rect 24213 2632 24225 2635
rect 23624 2604 24225 2632
rect 23624 2592 23630 2604
rect 24213 2601 24225 2604
rect 24259 2601 24271 2635
rect 24213 2595 24271 2601
rect 16761 2567 16819 2573
rect 16761 2533 16773 2567
rect 16807 2564 16819 2567
rect 18874 2564 18880 2576
rect 16807 2536 18880 2564
rect 16807 2533 16819 2536
rect 16761 2527 16819 2533
rect 18874 2524 18880 2536
rect 18932 2524 18938 2576
rect 19610 2524 19616 2576
rect 19668 2564 19674 2576
rect 19668 2536 22582 2564
rect 19668 2524 19674 2536
rect 17310 2496 17316 2508
rect 16684 2468 17316 2496
rect 16684 2437 16712 2468
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18012 2468 19656 2496
rect 18012 2456 18018 2468
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 16942 2388 16948 2440
rect 17000 2388 17006 2440
rect 17218 2388 17224 2440
rect 17276 2388 17282 2440
rect 18141 2431 18199 2437
rect 17512 2400 18092 2428
rect 17512 2360 17540 2400
rect 5552 2332 7880 2360
rect 8220 2332 8430 2360
rect 8496 2332 8984 2360
rect 9048 2332 9996 2360
rect 10060 2332 10732 2360
rect 11716 2332 15240 2360
rect 16546 2332 17540 2360
rect 17589 2363 17647 2369
rect 2740 2320 2746 2332
rect 584 2264 1624 2292
rect 4709 2295 4767 2301
rect 474 2184 480 2236
rect 532 2224 538 2236
rect 584 2224 612 2264
rect 4709 2261 4721 2295
rect 4755 2292 4767 2295
rect 5442 2292 5448 2304
rect 4755 2264 5448 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 5552 2301 5580 2332
rect 8220 2304 8248 2332
rect 8496 2304 8524 2332
rect 5537 2295 5595 2301
rect 5537 2261 5549 2295
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 6086 2292 6092 2304
rect 5868 2264 6092 2292
rect 5868 2252 5874 2264
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 6270 2252 6276 2304
rect 6328 2292 6334 2304
rect 7006 2292 7012 2304
rect 6328 2264 7012 2292
rect 6328 2252 6334 2264
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7190 2252 7196 2304
rect 7248 2252 7254 2304
rect 7466 2252 7472 2304
rect 7524 2252 7530 2304
rect 7558 2252 7564 2304
rect 7616 2292 7622 2304
rect 7745 2295 7803 2301
rect 7745 2292 7757 2295
rect 7616 2264 7757 2292
rect 7616 2252 7622 2264
rect 7745 2261 7757 2264
rect 7791 2261 7803 2295
rect 7745 2255 7803 2261
rect 7834 2252 7840 2304
rect 7892 2292 7898 2304
rect 8021 2295 8079 2301
rect 8021 2292 8033 2295
rect 7892 2264 8033 2292
rect 7892 2252 7898 2264
rect 8021 2261 8033 2264
rect 8067 2261 8079 2295
rect 8021 2255 8079 2261
rect 8202 2252 8208 2304
rect 8260 2252 8266 2304
rect 8294 2252 8300 2304
rect 8352 2252 8358 2304
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 8570 2252 8576 2304
rect 8628 2252 8634 2304
rect 8956 2301 8984 2332
rect 8941 2295 8999 2301
rect 8941 2261 8953 2295
rect 8987 2261 8999 2295
rect 8941 2255 8999 2261
rect 9858 2252 9864 2304
rect 9916 2292 9922 2304
rect 10060 2292 10088 2332
rect 11716 2304 11744 2332
rect 9916 2264 10088 2292
rect 9916 2252 9922 2264
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 11333 2295 11391 2301
rect 11333 2292 11345 2295
rect 10468 2264 11345 2292
rect 10468 2252 10474 2264
rect 11333 2261 11345 2264
rect 11379 2261 11391 2295
rect 11333 2255 11391 2261
rect 11606 2252 11612 2304
rect 11664 2252 11670 2304
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 12158 2252 12164 2304
rect 12216 2252 12222 2304
rect 12434 2252 12440 2304
rect 12492 2252 12498 2304
rect 12526 2252 12532 2304
rect 12584 2292 12590 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 12584 2264 12725 2292
rect 12584 2252 12590 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 13081 2295 13139 2301
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 13906 2292 13912 2304
rect 13127 2264 13912 2292
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 13906 2252 13912 2264
rect 13964 2252 13970 2304
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 14645 2295 14703 2301
rect 14645 2292 14657 2295
rect 14516 2264 14657 2292
rect 14516 2252 14522 2264
rect 14645 2261 14657 2264
rect 14691 2261 14703 2295
rect 14645 2255 14703 2261
rect 14918 2252 14924 2304
rect 14976 2252 14982 2304
rect 15212 2301 15240 2332
rect 17589 2329 17601 2363
rect 17635 2360 17647 2363
rect 17954 2360 17960 2372
rect 17635 2332 17960 2360
rect 17635 2329 17647 2332
rect 17589 2323 17647 2329
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 18064 2360 18092 2400
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18414 2428 18420 2440
rect 18187 2400 18420 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 18598 2388 18604 2440
rect 18656 2428 18662 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18656 2400 18705 2428
rect 18656 2388 18662 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 18693 2391 18751 2397
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19518 2388 19524 2440
rect 19576 2388 19582 2440
rect 19628 2428 19656 2468
rect 19794 2456 19800 2508
rect 19852 2456 19858 2508
rect 22462 2496 22468 2508
rect 20640 2468 22468 2496
rect 20640 2437 20668 2468
rect 22462 2456 22468 2468
rect 22520 2456 22526 2508
rect 22554 2496 22582 2536
rect 22554 2468 22968 2496
rect 20625 2431 20683 2437
rect 19628 2400 20024 2428
rect 19886 2360 19892 2372
rect 18064 2332 19892 2360
rect 19886 2320 19892 2332
rect 19944 2320 19950 2372
rect 15197 2295 15255 2301
rect 15197 2261 15209 2295
rect 15243 2261 15255 2295
rect 15197 2255 15255 2261
rect 15470 2252 15476 2304
rect 15528 2252 15534 2304
rect 16206 2252 16212 2304
rect 16264 2252 16270 2304
rect 16482 2252 16488 2304
rect 16540 2252 16546 2304
rect 17037 2295 17095 2301
rect 17037 2261 17049 2295
rect 17083 2292 17095 2295
rect 17494 2292 17500 2304
rect 17083 2264 17500 2292
rect 17083 2261 17095 2264
rect 17037 2255 17095 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 18414 2252 18420 2304
rect 18472 2292 18478 2304
rect 18785 2295 18843 2301
rect 18785 2292 18797 2295
rect 18472 2264 18797 2292
rect 18472 2252 18478 2264
rect 18785 2261 18797 2264
rect 18831 2261 18843 2295
rect 18785 2255 18843 2261
rect 19242 2252 19248 2304
rect 19300 2252 19306 2304
rect 19996 2292 20024 2400
rect 20625 2397 20637 2431
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20714 2388 20720 2440
rect 20772 2388 20778 2440
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 20956 2400 21281 2428
rect 20956 2388 20962 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21542 2388 21548 2440
rect 21600 2388 21606 2440
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22646 2428 22652 2440
rect 21876 2400 22652 2428
rect 21876 2388 21882 2400
rect 22646 2388 22652 2400
rect 22704 2428 22710 2440
rect 22833 2431 22891 2437
rect 22833 2428 22845 2431
rect 22704 2400 22845 2428
rect 22704 2388 22710 2400
rect 22833 2397 22845 2400
rect 22879 2397 22891 2431
rect 22940 2428 22968 2468
rect 23089 2431 23147 2437
rect 23089 2428 23101 2431
rect 22940 2400 23101 2428
rect 22833 2391 22891 2397
rect 23089 2397 23101 2400
rect 23135 2397 23147 2431
rect 23089 2391 23147 2397
rect 20732 2360 20760 2388
rect 22373 2363 22431 2369
rect 22373 2360 22385 2363
rect 20732 2332 22385 2360
rect 22373 2329 22385 2332
rect 22419 2329 22431 2363
rect 22373 2323 22431 2329
rect 21542 2292 21548 2304
rect 19996 2264 21548 2292
rect 21542 2252 21548 2264
rect 21600 2252 21606 2304
rect 23474 2252 23480 2304
rect 23532 2292 23538 2304
rect 25590 2292 25596 2304
rect 23532 2264 25596 2292
rect 23532 2252 23538 2264
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 532 2196 612 2224
rect 1104 2202 25000 2224
rect 532 2184 538 2196
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 842 2048 848 2100
rect 900 2088 906 2100
rect 900 2060 2268 2088
rect 900 2048 906 2060
rect 2240 2020 2268 2060
rect 2406 2048 2412 2100
rect 2464 2088 2470 2100
rect 2685 2091 2743 2097
rect 2685 2088 2697 2091
rect 2464 2060 2697 2088
rect 2464 2048 2470 2060
rect 2685 2057 2697 2060
rect 2731 2057 2743 2091
rect 2685 2051 2743 2057
rect 3513 2091 3571 2097
rect 3513 2057 3525 2091
rect 3559 2088 3571 2091
rect 3559 2060 4476 2088
rect 3559 2057 3571 2060
rect 3513 2051 3571 2057
rect 3881 2023 3939 2029
rect 3881 2020 3893 2023
rect 2240 1992 3893 2020
rect 1931 1985 1989 1991
rect 1302 1912 1308 1964
rect 1360 1912 1366 1964
rect 1394 1912 1400 1964
rect 1452 1912 1458 1964
rect 1931 1951 1943 1985
rect 1977 1982 1989 1985
rect 3881 1989 3893 1992
rect 3927 1989 3939 2023
rect 4448 2020 4476 2060
rect 4522 2048 4528 2100
rect 4580 2048 4586 2100
rect 5077 2091 5135 2097
rect 5077 2057 5089 2091
rect 5123 2057 5135 2091
rect 5077 2051 5135 2057
rect 5092 2020 5120 2051
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 5500 2060 6500 2088
rect 5500 2048 5506 2060
rect 5997 2023 6055 2029
rect 5997 2020 6009 2023
rect 4448 1992 4936 2020
rect 5092 1992 6009 2020
rect 3881 1983 3939 1989
rect 1977 1952 1992 1982
rect 2038 1952 2044 1964
rect 1977 1951 2044 1952
rect 1931 1945 2044 1951
rect 1964 1924 2044 1945
rect 2038 1912 2044 1924
rect 2096 1912 2102 1964
rect 3234 1912 3240 1964
rect 3292 1912 3298 1964
rect 3694 1912 3700 1964
rect 3752 1912 3758 1964
rect 4433 1955 4491 1961
rect 4433 1952 4445 1955
rect 3988 1924 4445 1952
rect 1320 1884 1348 1912
rect 1673 1887 1731 1893
rect 1673 1884 1685 1887
rect 1320 1856 1685 1884
rect 1673 1853 1685 1856
rect 1719 1853 1731 1887
rect 1673 1847 1731 1853
rect 3786 1844 3792 1896
rect 3844 1884 3850 1896
rect 3988 1884 4016 1924
rect 4433 1921 4445 1924
rect 4479 1921 4491 1955
rect 4706 1952 4712 1964
rect 4433 1915 4491 1921
rect 4540 1924 4712 1952
rect 3844 1856 4016 1884
rect 4157 1887 4215 1893
rect 3844 1844 3850 1856
rect 4157 1853 4169 1887
rect 4203 1884 4215 1887
rect 4540 1884 4568 1924
rect 4706 1912 4712 1924
rect 4764 1912 4770 1964
rect 4798 1912 4804 1964
rect 4856 1912 4862 1964
rect 4203 1856 4568 1884
rect 4203 1853 4215 1856
rect 4157 1847 4215 1853
rect 4614 1844 4620 1896
rect 4672 1844 4678 1896
rect 3421 1819 3479 1825
rect 3421 1785 3433 1819
rect 3467 1816 3479 1819
rect 4632 1816 4660 1844
rect 3467 1788 4660 1816
rect 3467 1785 3479 1788
rect 3421 1779 3479 1785
rect 1581 1751 1639 1757
rect 1581 1717 1593 1751
rect 1627 1748 1639 1751
rect 3050 1748 3056 1760
rect 1627 1720 3056 1748
rect 1627 1717 1639 1720
rect 1581 1711 1639 1717
rect 3050 1708 3056 1720
rect 3108 1708 3114 1760
rect 4908 1748 4936 1992
rect 5997 1989 6009 1992
rect 6043 1989 6055 2023
rect 5997 1983 6055 1989
rect 6178 1980 6184 2032
rect 6236 1980 6242 2032
rect 6472 2029 6500 2060
rect 6546 2048 6552 2100
rect 6604 2048 6610 2100
rect 7558 2088 7564 2100
rect 6748 2060 7564 2088
rect 6457 2023 6515 2029
rect 6457 1989 6469 2023
rect 6503 1989 6515 2023
rect 6457 1983 6515 1989
rect 5261 1955 5319 1961
rect 5261 1921 5273 1955
rect 5307 1921 5319 1955
rect 5261 1915 5319 1921
rect 5445 1955 5503 1961
rect 5445 1921 5457 1955
rect 5491 1952 5503 1955
rect 5718 1952 5724 1964
rect 5491 1924 5724 1952
rect 5491 1921 5503 1924
rect 5445 1915 5503 1921
rect 5276 1884 5304 1915
rect 5718 1912 5724 1924
rect 5776 1912 5782 1964
rect 5902 1912 5908 1964
rect 5960 1912 5966 1964
rect 6748 1961 6776 2060
rect 7558 2048 7564 2060
rect 7616 2048 7622 2100
rect 7653 2091 7711 2097
rect 7653 2057 7665 2091
rect 7699 2088 7711 2091
rect 7742 2088 7748 2100
rect 7699 2060 7748 2088
rect 7699 2057 7711 2060
rect 7653 2051 7711 2057
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 7834 2048 7840 2100
rect 7892 2048 7898 2100
rect 8021 2091 8079 2097
rect 8021 2057 8033 2091
rect 8067 2088 8079 2091
rect 8110 2088 8116 2100
rect 8067 2060 8116 2088
rect 8067 2057 8079 2060
rect 8021 2051 8079 2057
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 8386 2048 8392 2100
rect 8444 2048 8450 2100
rect 8478 2048 8484 2100
rect 8536 2048 8542 2100
rect 8570 2048 8576 2100
rect 8628 2048 8634 2100
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2088 8815 2091
rect 8846 2088 8852 2100
rect 8803 2060 8852 2088
rect 8803 2057 8815 2060
rect 8757 2051 8815 2057
rect 8846 2048 8852 2060
rect 8904 2048 8910 2100
rect 9953 2091 10011 2097
rect 9953 2057 9965 2091
rect 9999 2088 10011 2091
rect 10226 2088 10232 2100
rect 9999 2060 10232 2088
rect 9999 2057 10011 2060
rect 9953 2051 10011 2057
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 11606 2048 11612 2100
rect 11664 2088 11670 2100
rect 11664 2060 12020 2088
rect 11664 2048 11670 2060
rect 7852 2020 7880 2048
rect 7116 1992 7880 2020
rect 7929 2023 7987 2029
rect 7116 1961 7144 1992
rect 7929 1989 7941 2023
rect 7975 2020 7987 2023
rect 8496 2020 8524 2048
rect 7975 1992 8524 2020
rect 7975 1989 7987 1992
rect 7929 1983 7987 1989
rect 6733 1955 6791 1961
rect 6733 1921 6745 1955
rect 6779 1921 6791 1955
rect 6733 1915 6791 1921
rect 7101 1955 7159 1961
rect 7101 1921 7113 1955
rect 7147 1921 7159 1955
rect 7561 1955 7619 1961
rect 7101 1915 7159 1921
rect 7208 1924 7512 1952
rect 5810 1884 5816 1896
rect 5276 1856 5816 1884
rect 5810 1844 5816 1856
rect 5868 1844 5874 1896
rect 4985 1819 5043 1825
rect 4985 1785 4997 1819
rect 5031 1816 5043 1819
rect 5920 1816 5948 1912
rect 6454 1844 6460 1896
rect 6512 1844 6518 1896
rect 6472 1816 6500 1844
rect 5031 1788 5948 1816
rect 6012 1788 6500 1816
rect 6917 1819 6975 1825
rect 5031 1785 5043 1788
rect 4985 1779 5043 1785
rect 5534 1748 5540 1760
rect 4908 1720 5540 1748
rect 5534 1708 5540 1720
rect 5592 1708 5598 1760
rect 5721 1751 5779 1757
rect 5721 1717 5733 1751
rect 5767 1748 5779 1751
rect 6012 1748 6040 1788
rect 6917 1785 6929 1819
rect 6963 1816 6975 1819
rect 7208 1816 7236 1924
rect 6963 1788 7236 1816
rect 6963 1785 6975 1788
rect 6917 1779 6975 1785
rect 7282 1776 7288 1828
rect 7340 1776 7346 1828
rect 7484 1816 7512 1924
rect 7561 1921 7573 1955
rect 7607 1921 7619 1955
rect 7561 1915 7619 1921
rect 8205 1955 8263 1961
rect 8205 1921 8217 1955
rect 8251 1952 8263 1955
rect 8478 1952 8484 1964
rect 8251 1924 8484 1952
rect 8251 1921 8263 1924
rect 8205 1915 8263 1921
rect 7576 1884 7604 1915
rect 8478 1912 8484 1924
rect 8536 1912 8542 1964
rect 8588 1884 8616 2048
rect 8662 1980 8668 2032
rect 8720 1980 8726 2032
rect 9214 1991 9220 2032
rect 9199 1985 9220 1991
rect 8938 1912 8944 1964
rect 8996 1912 9002 1964
rect 9199 1951 9211 1985
rect 9272 1980 9278 2032
rect 9398 1980 9404 2032
rect 9456 2020 9462 2032
rect 10413 2023 10471 2029
rect 10413 2020 10425 2023
rect 9456 1992 10425 2020
rect 9456 1980 9462 1992
rect 10413 1989 10425 1992
rect 10459 1989 10471 2023
rect 10413 1983 10471 1989
rect 10965 2023 11023 2029
rect 10965 1989 10977 2023
rect 11011 2020 11023 2023
rect 11698 2020 11704 2032
rect 11011 1992 11704 2020
rect 11011 1989 11023 1992
rect 10965 1983 11023 1989
rect 11698 1980 11704 1992
rect 11756 1980 11762 2032
rect 11992 2029 12020 2060
rect 12434 2048 12440 2100
rect 12492 2048 12498 2100
rect 13538 2048 13544 2100
rect 13596 2048 13602 2100
rect 14734 2088 14740 2100
rect 13832 2060 14740 2088
rect 11977 2023 12035 2029
rect 11977 1989 11989 2023
rect 12023 1989 12035 2023
rect 12452 2020 12480 2048
rect 12805 2023 12863 2029
rect 12805 2020 12817 2023
rect 12452 1992 12817 2020
rect 11977 1983 12035 1989
rect 12805 1989 12817 1992
rect 12851 1989 12863 2023
rect 13556 2020 13584 2048
rect 12805 1983 12863 1989
rect 13096 1992 13584 2020
rect 9245 1954 9260 1980
rect 9245 1951 9257 1954
rect 9199 1945 9257 1951
rect 11790 1912 11796 1964
rect 11848 1912 11854 1964
rect 12621 1955 12679 1961
rect 12621 1921 12633 1955
rect 12667 1952 12679 1955
rect 13096 1952 13124 1992
rect 12667 1924 13124 1952
rect 12667 1921 12679 1924
rect 12621 1915 12679 1921
rect 13538 1912 13544 1964
rect 13596 1912 13602 1964
rect 13832 1961 13860 2060
rect 14734 2048 14740 2060
rect 14792 2048 14798 2100
rect 14918 2048 14924 2100
rect 14976 2048 14982 2100
rect 15197 2091 15255 2097
rect 15197 2057 15209 2091
rect 15243 2057 15255 2091
rect 15197 2051 15255 2057
rect 14936 2020 14964 2048
rect 14476 1992 14964 2020
rect 14476 1961 14504 1992
rect 13817 1955 13875 1961
rect 13817 1921 13829 1955
rect 13863 1921 13875 1955
rect 13817 1915 13875 1921
rect 14277 1955 14335 1961
rect 14277 1921 14289 1955
rect 14323 1921 14335 1955
rect 14277 1915 14335 1921
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1952 14887 1955
rect 15212 1952 15240 2051
rect 15470 2048 15476 2100
rect 15528 2048 15534 2100
rect 17954 2048 17960 2100
rect 18012 2088 18018 2100
rect 18325 2091 18383 2097
rect 18325 2088 18337 2091
rect 18012 2060 18337 2088
rect 18012 2048 18018 2060
rect 18325 2057 18337 2060
rect 18371 2057 18383 2091
rect 18325 2051 18383 2057
rect 19242 2048 19248 2100
rect 19300 2048 19306 2100
rect 19518 2048 19524 2100
rect 19576 2088 19582 2100
rect 19576 2060 22784 2088
rect 19576 2048 19582 2060
rect 15488 2020 15516 2048
rect 15488 1992 16160 2020
rect 14875 1924 15240 1952
rect 14875 1921 14887 1924
rect 14829 1915 14887 1921
rect 7576 1856 8616 1884
rect 9674 1844 9680 1896
rect 9732 1884 9738 1896
rect 10502 1884 10508 1896
rect 9732 1856 10508 1884
rect 9732 1844 9738 1856
rect 10502 1844 10508 1856
rect 10560 1844 10566 1896
rect 14292 1884 14320 1915
rect 15378 1912 15384 1964
rect 15436 1912 15442 1964
rect 16132 1961 16160 1992
rect 16758 1980 16764 2032
rect 16816 1980 16822 2032
rect 17770 1980 17776 2032
rect 17828 2020 17834 2032
rect 17865 2023 17923 2029
rect 17865 2020 17877 2023
rect 17828 1992 17877 2020
rect 17828 1980 17834 1992
rect 17865 1989 17877 1992
rect 17911 1989 17923 2023
rect 19260 2020 19288 2048
rect 17865 1983 17923 1989
rect 18248 1992 19288 2020
rect 19628 1992 21312 2020
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1921 15715 1955
rect 15657 1915 15715 1921
rect 16117 1955 16175 1961
rect 16117 1921 16129 1955
rect 16163 1921 16175 1955
rect 16117 1915 16175 1921
rect 17313 1955 17371 1961
rect 17313 1921 17325 1955
rect 17359 1952 17371 1955
rect 18248 1952 18276 1992
rect 17359 1924 18276 1952
rect 17359 1921 17371 1924
rect 17313 1915 17371 1921
rect 15010 1884 15016 1896
rect 14292 1856 15016 1884
rect 15010 1844 15016 1856
rect 15068 1844 15074 1896
rect 15672 1884 15700 1915
rect 18506 1912 18512 1964
rect 18564 1912 18570 1964
rect 19628 1952 19656 1992
rect 18616 1924 19656 1952
rect 19705 1955 19763 1961
rect 16298 1884 16304 1896
rect 15672 1856 16304 1884
rect 16298 1844 16304 1856
rect 16356 1844 16362 1896
rect 18616 1893 18644 1924
rect 19705 1921 19717 1955
rect 19751 1921 19763 1955
rect 19705 1915 19763 1921
rect 18601 1887 18659 1893
rect 18601 1853 18613 1887
rect 18647 1853 18659 1887
rect 18601 1847 18659 1853
rect 18877 1887 18935 1893
rect 18877 1853 18889 1887
rect 18923 1884 18935 1887
rect 19426 1884 19432 1896
rect 18923 1856 19432 1884
rect 18923 1853 18935 1856
rect 18877 1847 18935 1853
rect 19426 1844 19432 1856
rect 19484 1844 19490 1896
rect 7650 1816 7656 1828
rect 7484 1788 7656 1816
rect 7650 1776 7656 1788
rect 7708 1776 7714 1828
rect 8478 1776 8484 1828
rect 8536 1816 8542 1828
rect 8846 1816 8852 1828
rect 8536 1788 8852 1816
rect 8536 1776 8542 1788
rect 8846 1776 8852 1788
rect 8904 1776 8910 1828
rect 13357 1819 13415 1825
rect 13357 1785 13369 1819
rect 13403 1816 13415 1819
rect 13998 1816 14004 1828
rect 13403 1788 14004 1816
rect 13403 1785 13415 1788
rect 13357 1779 13415 1785
rect 13998 1776 14004 1788
rect 14056 1776 14062 1828
rect 15378 1776 15384 1828
rect 15436 1816 15442 1828
rect 15436 1788 16344 1816
rect 15436 1776 15442 1788
rect 5767 1720 6040 1748
rect 5767 1717 5779 1720
rect 5721 1711 5779 1717
rect 6086 1708 6092 1760
rect 6144 1748 6150 1760
rect 9858 1748 9864 1760
rect 6144 1720 9864 1748
rect 6144 1708 6150 1720
rect 9858 1708 9864 1720
rect 9916 1708 9922 1760
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 10962 1708 10968 1760
rect 11020 1748 11026 1760
rect 11057 1751 11115 1757
rect 11057 1748 11069 1751
rect 11020 1720 11069 1748
rect 11020 1708 11026 1720
rect 11057 1717 11069 1720
rect 11103 1717 11115 1751
rect 11057 1711 11115 1717
rect 11609 1751 11667 1757
rect 11609 1717 11621 1751
rect 11655 1748 11667 1751
rect 11790 1748 11796 1760
rect 11655 1720 11796 1748
rect 11655 1717 11667 1720
rect 11609 1711 11667 1717
rect 11790 1708 11796 1720
rect 11848 1708 11854 1760
rect 12066 1708 12072 1760
rect 12124 1708 12130 1760
rect 12434 1708 12440 1760
rect 12492 1708 12498 1760
rect 12618 1708 12624 1760
rect 12676 1748 12682 1760
rect 12897 1751 12955 1757
rect 12897 1748 12909 1751
rect 12676 1720 12909 1748
rect 12676 1708 12682 1720
rect 12897 1717 12909 1720
rect 12943 1717 12955 1751
rect 12897 1711 12955 1717
rect 13630 1708 13636 1760
rect 13688 1708 13694 1760
rect 14090 1708 14096 1760
rect 14148 1708 14154 1760
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14645 1751 14703 1757
rect 14645 1748 14657 1751
rect 14332 1720 14657 1748
rect 14332 1708 14338 1720
rect 14645 1717 14657 1720
rect 14691 1717 14703 1751
rect 14645 1711 14703 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15746 1708 15752 1760
rect 15804 1708 15810 1760
rect 16316 1757 16344 1788
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1717 16359 1751
rect 16301 1711 16359 1717
rect 16850 1708 16856 1760
rect 16908 1708 16914 1760
rect 17402 1708 17408 1760
rect 17460 1708 17466 1760
rect 17586 1708 17592 1760
rect 17644 1748 17650 1760
rect 17957 1751 18015 1757
rect 17957 1748 17969 1751
rect 17644 1720 17969 1748
rect 17644 1708 17650 1720
rect 17957 1717 17969 1720
rect 18003 1717 18015 1751
rect 19720 1748 19748 1915
rect 19886 1912 19892 1964
rect 19944 1912 19950 1964
rect 20809 1955 20867 1961
rect 20809 1921 20821 1955
rect 20855 1952 20867 1955
rect 20898 1952 20904 1964
rect 20855 1924 20904 1952
rect 20855 1921 20867 1924
rect 20809 1915 20867 1921
rect 20898 1912 20904 1924
rect 20956 1912 20962 1964
rect 21284 1952 21312 1992
rect 21358 1980 21364 2032
rect 21416 2020 21422 2032
rect 21453 2023 21511 2029
rect 21453 2020 21465 2023
rect 21416 1992 21465 2020
rect 21416 1980 21422 1992
rect 21453 1989 21465 1992
rect 21499 1989 21511 2023
rect 21453 1983 21511 1989
rect 21542 1980 21548 2032
rect 21600 2020 21606 2032
rect 22066 2023 22124 2029
rect 22066 2020 22078 2023
rect 21600 1992 22078 2020
rect 21600 1980 21606 1992
rect 22066 1989 22078 1992
rect 22112 1989 22124 2023
rect 22756 2020 22784 2060
rect 22830 2048 22836 2100
rect 22888 2088 22894 2100
rect 23201 2091 23259 2097
rect 23201 2088 23213 2091
rect 22888 2060 23213 2088
rect 22888 2048 22894 2060
rect 23201 2057 23213 2060
rect 23247 2057 23259 2091
rect 23201 2051 23259 2057
rect 23014 2020 23020 2032
rect 22756 1992 23020 2020
rect 22066 1983 22124 1989
rect 23014 1980 23020 1992
rect 23072 1980 23078 2032
rect 25130 2020 25136 2032
rect 23216 1992 25136 2020
rect 23216 1952 23244 1992
rect 25130 1980 25136 1992
rect 25188 1980 25194 2032
rect 21284 1924 23244 1952
rect 23293 1955 23351 1961
rect 23293 1921 23305 1955
rect 23339 1921 23351 1955
rect 23293 1915 23351 1921
rect 19904 1884 19932 1912
rect 19981 1887 20039 1893
rect 19981 1884 19993 1887
rect 19904 1856 19993 1884
rect 19981 1853 19993 1856
rect 20027 1853 20039 1887
rect 19981 1847 20039 1853
rect 20070 1844 20076 1896
rect 20128 1844 20134 1896
rect 21266 1844 21272 1896
rect 21324 1884 21330 1896
rect 21542 1884 21548 1896
rect 21324 1856 21548 1884
rect 21324 1844 21330 1856
rect 21542 1844 21548 1856
rect 21600 1844 21606 1896
rect 21818 1844 21824 1896
rect 21876 1844 21882 1896
rect 20088 1816 20116 1844
rect 21836 1816 21864 1844
rect 23308 1816 23336 1915
rect 23658 1912 23664 1964
rect 23716 1912 23722 1964
rect 23676 1884 23704 1912
rect 23753 1887 23811 1893
rect 23753 1884 23765 1887
rect 23676 1856 23765 1884
rect 23753 1853 23765 1856
rect 23799 1853 23811 1887
rect 23753 1847 23811 1853
rect 20088 1788 21864 1816
rect 22756 1788 23336 1816
rect 20346 1748 20352 1760
rect 19720 1720 20352 1748
rect 17957 1711 18015 1717
rect 20346 1708 20352 1720
rect 20404 1708 20410 1760
rect 20622 1708 20628 1760
rect 20680 1748 20686 1760
rect 22756 1748 22784 1788
rect 20680 1720 22784 1748
rect 20680 1708 20686 1720
rect 23014 1708 23020 1760
rect 23072 1748 23078 1760
rect 24854 1748 24860 1760
rect 23072 1720 24860 1748
rect 23072 1708 23078 1720
rect 24854 1708 24860 1720
rect 24912 1708 24918 1760
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 1581 1547 1639 1553
rect 1581 1513 1593 1547
rect 1627 1544 1639 1547
rect 3326 1544 3332 1556
rect 1627 1516 3332 1544
rect 1627 1513 1639 1516
rect 1581 1507 1639 1513
rect 3326 1504 3332 1516
rect 3384 1504 3390 1556
rect 4890 1504 4896 1556
rect 4948 1544 4954 1556
rect 7282 1544 7288 1556
rect 4948 1516 7288 1544
rect 4948 1504 4954 1516
rect 7282 1504 7288 1516
rect 7340 1504 7346 1556
rect 8662 1504 8668 1556
rect 8720 1504 8726 1556
rect 8846 1504 8852 1556
rect 8904 1544 8910 1556
rect 9490 1544 9496 1556
rect 8904 1516 9496 1544
rect 8904 1504 8910 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 13722 1504 13728 1556
rect 13780 1544 13786 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13780 1516 14289 1544
rect 13780 1504 13786 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 15102 1504 15108 1556
rect 15160 1544 15166 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 15160 1516 15393 1544
rect 15160 1504 15166 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 750 1436 756 1488
rect 808 1476 814 1488
rect 2501 1479 2559 1485
rect 2501 1476 2513 1479
rect 808 1448 2513 1476
rect 808 1436 814 1448
rect 2501 1445 2513 1448
rect 2547 1445 2559 1479
rect 2501 1439 2559 1445
rect 5810 1436 5816 1488
rect 5868 1476 5874 1488
rect 6638 1476 6644 1488
rect 5868 1448 6644 1476
rect 5868 1436 5874 1448
rect 6638 1436 6644 1448
rect 6696 1436 6702 1488
rect 6730 1436 6736 1488
rect 6788 1476 6794 1488
rect 11422 1476 11428 1488
rect 6788 1448 11428 1476
rect 6788 1436 6794 1448
rect 11422 1436 11428 1448
rect 11480 1436 11486 1488
rect 11517 1479 11575 1485
rect 11517 1445 11529 1479
rect 11563 1445 11575 1479
rect 11517 1439 11575 1445
rect 9585 1411 9643 1417
rect 9585 1377 9597 1411
rect 9631 1408 9643 1411
rect 10042 1408 10048 1420
rect 9631 1380 10048 1408
rect 9631 1377 9643 1380
rect 9585 1371 9643 1377
rect 10042 1368 10048 1380
rect 10100 1368 10106 1420
rect 10873 1411 10931 1417
rect 10873 1377 10885 1411
rect 10919 1408 10931 1411
rect 11146 1408 11152 1420
rect 10919 1380 11152 1408
rect 10919 1377 10931 1380
rect 10873 1371 10931 1377
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 1394 1300 1400 1352
rect 1452 1300 1458 1352
rect 1946 1300 1952 1352
rect 2004 1300 2010 1352
rect 2038 1300 2044 1352
rect 2096 1340 2102 1352
rect 2096 1312 2728 1340
rect 2096 1300 2102 1312
rect 1762 1232 1768 1284
rect 1820 1232 1826 1284
rect 2314 1232 2320 1284
rect 2372 1232 2378 1284
rect 2700 1281 2728 1312
rect 3050 1300 3056 1352
rect 3108 1300 3114 1352
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1309 3663 1343
rect 3605 1303 3663 1309
rect 2685 1275 2743 1281
rect 2685 1241 2697 1275
rect 2731 1241 2743 1275
rect 3620 1272 3648 1303
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4062 1300 4068 1352
rect 4120 1300 4126 1352
rect 5258 1300 5264 1352
rect 5316 1300 5322 1352
rect 5534 1300 5540 1352
rect 5592 1300 5598 1352
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 7009 1343 7067 1349
rect 7009 1309 7021 1343
rect 7055 1340 7067 1343
rect 7466 1340 7472 1352
rect 7055 1312 7472 1340
rect 7055 1309 7067 1312
rect 7009 1303 7067 1309
rect 7466 1300 7472 1312
rect 7524 1300 7530 1352
rect 7926 1300 7932 1352
rect 7984 1300 7990 1352
rect 8294 1300 8300 1352
rect 8352 1300 8358 1352
rect 8386 1300 8392 1352
rect 8444 1300 8450 1352
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 9125 1343 9183 1349
rect 8527 1312 8984 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 4522 1272 4528 1284
rect 2685 1235 2743 1241
rect 3252 1244 3556 1272
rect 3620 1244 4528 1272
rect 2774 1164 2780 1216
rect 2832 1164 2838 1216
rect 3252 1213 3280 1244
rect 3237 1207 3295 1213
rect 3237 1173 3249 1207
rect 3283 1173 3295 1207
rect 3237 1167 3295 1173
rect 3418 1164 3424 1216
rect 3476 1164 3482 1216
rect 3528 1204 3556 1244
rect 4522 1232 4528 1244
rect 4580 1232 4586 1284
rect 4985 1275 5043 1281
rect 4985 1241 4997 1275
rect 5031 1272 5043 1275
rect 5626 1272 5632 1284
rect 5031 1244 5632 1272
rect 5031 1241 5043 1244
rect 4985 1235 5043 1241
rect 5626 1232 5632 1244
rect 5684 1232 5690 1284
rect 6454 1232 6460 1284
rect 6512 1272 6518 1284
rect 7377 1275 7435 1281
rect 7377 1272 7389 1275
rect 6512 1244 7389 1272
rect 6512 1232 6518 1244
rect 7377 1241 7389 1244
rect 7423 1241 7435 1275
rect 7377 1235 7435 1241
rect 7745 1275 7803 1281
rect 7745 1241 7757 1275
rect 7791 1272 7803 1275
rect 8312 1272 8340 1300
rect 7791 1244 8340 1272
rect 7791 1241 7803 1244
rect 7745 1235 7803 1241
rect 8846 1232 8852 1284
rect 8904 1232 8910 1284
rect 3970 1204 3976 1216
rect 3528 1176 3976 1204
rect 3970 1164 3976 1176
rect 4028 1164 4034 1216
rect 5077 1207 5135 1213
rect 5077 1173 5089 1207
rect 5123 1204 5135 1207
rect 5166 1204 5172 1216
rect 5123 1176 5172 1204
rect 5123 1173 5135 1176
rect 5077 1167 5135 1173
rect 5166 1164 5172 1176
rect 5224 1164 5230 1216
rect 6546 1164 6552 1216
rect 6604 1164 6610 1216
rect 6730 1164 6736 1216
rect 6788 1204 6794 1216
rect 7101 1207 7159 1213
rect 7101 1204 7113 1207
rect 6788 1176 7113 1204
rect 6788 1164 6794 1176
rect 7101 1173 7113 1176
rect 7147 1173 7159 1207
rect 7101 1167 7159 1173
rect 7466 1164 7472 1216
rect 7524 1164 7530 1216
rect 8205 1207 8263 1213
rect 8205 1173 8217 1207
rect 8251 1204 8263 1207
rect 8864 1204 8892 1232
rect 8956 1213 8984 1312
rect 9125 1309 9137 1343
rect 9171 1340 9183 1343
rect 9674 1340 9680 1352
rect 9171 1312 9680 1340
rect 9171 1309 9183 1312
rect 9125 1303 9183 1309
rect 9674 1300 9680 1312
rect 9732 1300 9738 1352
rect 9769 1343 9827 1349
rect 9769 1309 9781 1343
rect 9815 1340 9827 1343
rect 9950 1340 9956 1352
rect 9815 1312 9956 1340
rect 9815 1309 9827 1312
rect 9769 1303 9827 1309
rect 9950 1300 9956 1312
rect 10008 1300 10014 1352
rect 10137 1343 10195 1349
rect 10137 1309 10149 1343
rect 10183 1340 10195 1343
rect 10410 1340 10416 1352
rect 10183 1312 10416 1340
rect 10183 1309 10195 1312
rect 10137 1303 10195 1309
rect 10410 1300 10416 1312
rect 10468 1300 10474 1352
rect 10597 1343 10655 1349
rect 10597 1309 10609 1343
rect 10643 1309 10655 1343
rect 10597 1303 10655 1309
rect 11057 1343 11115 1349
rect 11057 1309 11069 1343
rect 11103 1340 11115 1343
rect 11532 1340 11560 1439
rect 14090 1436 14096 1488
rect 14148 1436 14154 1488
rect 15194 1436 15200 1488
rect 15252 1476 15258 1488
rect 15948 1476 15976 1507
rect 16298 1504 16304 1556
rect 16356 1504 16362 1556
rect 16666 1504 16672 1556
rect 16724 1544 16730 1556
rect 17957 1547 18015 1553
rect 17957 1544 17969 1547
rect 16724 1516 17969 1544
rect 16724 1504 16730 1516
rect 17957 1513 17969 1516
rect 18003 1513 18015 1547
rect 17957 1507 18015 1513
rect 18509 1547 18567 1553
rect 18509 1513 18521 1547
rect 18555 1513 18567 1547
rect 18509 1507 18567 1513
rect 15252 1448 15976 1476
rect 15252 1436 15258 1448
rect 16114 1436 16120 1488
rect 16172 1476 16178 1488
rect 16945 1479 17003 1485
rect 16945 1476 16957 1479
rect 16172 1448 16957 1476
rect 16172 1436 16178 1448
rect 16945 1445 16957 1448
rect 16991 1445 17003 1479
rect 16945 1439 17003 1445
rect 17497 1479 17555 1485
rect 17497 1445 17509 1479
rect 17543 1445 17555 1479
rect 17497 1439 17555 1445
rect 14108 1408 14136 1436
rect 12084 1380 13032 1408
rect 14108 1380 14780 1408
rect 11103 1312 11560 1340
rect 11103 1309 11115 1312
rect 11057 1303 11115 1309
rect 9309 1275 9367 1281
rect 9309 1241 9321 1275
rect 9355 1241 9367 1275
rect 10612 1272 10640 1303
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 12084 1340 12112 1380
rect 11900 1312 12112 1340
rect 11900 1272 11928 1312
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 12253 1343 12311 1349
rect 12253 1340 12265 1343
rect 12216 1312 12265 1340
rect 12216 1300 12222 1312
rect 12253 1309 12265 1312
rect 12299 1309 12311 1343
rect 12253 1303 12311 1309
rect 12434 1300 12440 1352
rect 12492 1340 12498 1352
rect 12897 1343 12955 1349
rect 12897 1340 12909 1343
rect 12492 1312 12909 1340
rect 12492 1300 12498 1312
rect 12897 1309 12909 1312
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 12710 1272 12716 1284
rect 9309 1235 9367 1241
rect 9968 1244 10548 1272
rect 10612 1244 11928 1272
rect 11992 1244 12716 1272
rect 8251 1176 8892 1204
rect 8941 1207 8999 1213
rect 8251 1173 8263 1176
rect 8205 1167 8263 1173
rect 8941 1173 8953 1207
rect 8987 1173 8999 1207
rect 9324 1204 9352 1235
rect 9766 1204 9772 1216
rect 9324 1176 9772 1204
rect 8941 1167 8999 1173
rect 9766 1164 9772 1176
rect 9824 1164 9830 1216
rect 9968 1213 9996 1244
rect 9953 1207 10011 1213
rect 9953 1173 9965 1207
rect 9999 1173 10011 1207
rect 9953 1167 10011 1173
rect 10318 1164 10324 1216
rect 10376 1164 10382 1216
rect 10520 1204 10548 1244
rect 10686 1204 10692 1216
rect 10520 1176 10692 1204
rect 10686 1164 10692 1176
rect 10744 1164 10750 1216
rect 11238 1164 11244 1216
rect 11296 1164 11302 1216
rect 11992 1213 12020 1244
rect 12710 1232 12716 1244
rect 12768 1232 12774 1284
rect 13004 1272 13032 1380
rect 13265 1343 13323 1349
rect 13265 1309 13277 1343
rect 13311 1340 13323 1343
rect 13630 1340 13636 1352
rect 13311 1312 13636 1340
rect 13311 1309 13323 1312
rect 13265 1303 13323 1309
rect 13630 1300 13636 1312
rect 13688 1300 13694 1352
rect 13814 1300 13820 1352
rect 13872 1300 13878 1352
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 13998 1300 14004 1352
rect 14056 1340 14062 1352
rect 14645 1343 14703 1349
rect 14645 1340 14657 1343
rect 14056 1312 14657 1340
rect 14056 1300 14062 1312
rect 14645 1309 14657 1312
rect 14691 1309 14703 1343
rect 14752 1340 14780 1380
rect 16390 1368 16396 1420
rect 16448 1408 16454 1420
rect 17512 1408 17540 1439
rect 17862 1436 17868 1488
rect 17920 1476 17926 1488
rect 18524 1476 18552 1507
rect 19426 1504 19432 1556
rect 19484 1544 19490 1556
rect 20162 1544 20168 1556
rect 19484 1516 20168 1544
rect 19484 1504 19490 1516
rect 20162 1504 20168 1516
rect 20220 1504 20226 1556
rect 20530 1504 20536 1556
rect 20588 1504 20594 1556
rect 22370 1504 22376 1556
rect 22428 1504 22434 1556
rect 22462 1504 22468 1556
rect 22520 1544 22526 1556
rect 22830 1544 22836 1556
rect 22520 1516 22836 1544
rect 22520 1504 22526 1516
rect 22830 1504 22836 1516
rect 22888 1504 22894 1556
rect 22094 1476 22100 1488
rect 17920 1448 18552 1476
rect 21560 1448 22100 1476
rect 17920 1436 17926 1448
rect 16448 1380 17540 1408
rect 16448 1368 16454 1380
rect 17678 1368 17684 1420
rect 17736 1408 17742 1420
rect 21358 1408 21364 1420
rect 17736 1380 21364 1408
rect 17736 1368 17742 1380
rect 21358 1368 21364 1380
rect 21416 1368 21422 1420
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 14752 1312 15301 1340
rect 14645 1303 14703 1309
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 16482 1300 16488 1352
rect 16540 1300 16546 1352
rect 16574 1300 16580 1352
rect 16632 1340 16638 1352
rect 17313 1343 17371 1349
rect 17313 1340 17325 1343
rect 16632 1312 17325 1340
rect 16632 1300 16638 1312
rect 17313 1309 17325 1312
rect 17359 1309 17371 1343
rect 17313 1303 17371 1309
rect 17494 1300 17500 1352
rect 17552 1340 17558 1352
rect 17865 1343 17923 1349
rect 17865 1340 17877 1343
rect 17552 1312 17877 1340
rect 17552 1300 17558 1312
rect 17865 1309 17877 1312
rect 17911 1309 17923 1343
rect 17865 1303 17923 1309
rect 18322 1300 18328 1352
rect 18380 1340 18386 1352
rect 18417 1343 18475 1349
rect 18417 1340 18429 1343
rect 18380 1312 18429 1340
rect 18380 1300 18386 1312
rect 18417 1309 18429 1312
rect 18463 1309 18475 1343
rect 18417 1303 18475 1309
rect 18877 1343 18935 1349
rect 18877 1309 18889 1343
rect 18923 1340 18935 1343
rect 20530 1340 20536 1352
rect 18923 1312 20536 1340
rect 18923 1309 18935 1312
rect 18877 1303 18935 1309
rect 20530 1300 20536 1312
rect 20588 1300 20594 1352
rect 21453 1343 21511 1349
rect 21453 1309 21465 1343
rect 21499 1340 21511 1343
rect 21560 1340 21588 1448
rect 22094 1436 22100 1448
rect 22152 1436 22158 1488
rect 22388 1476 22416 1504
rect 22296 1448 22416 1476
rect 21499 1312 21588 1340
rect 21499 1309 21511 1312
rect 21453 1303 21511 1309
rect 21634 1300 21640 1352
rect 21692 1300 21698 1352
rect 22189 1343 22247 1349
rect 22189 1309 22201 1343
rect 22235 1309 22247 1343
rect 22296 1340 22324 1448
rect 25038 1368 25044 1420
rect 25096 1368 25102 1420
rect 22364 1343 22422 1349
rect 22364 1340 22376 1343
rect 22296 1312 22376 1340
rect 22189 1303 22247 1309
rect 22364 1309 22376 1312
rect 22410 1309 22422 1343
rect 22364 1303 22422 1309
rect 13924 1272 13952 1300
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 13004 1244 13676 1272
rect 13924 1244 14197 1272
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 12342 1164 12348 1216
rect 12400 1164 12406 1216
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13648 1213 13676 1244
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14185 1235 14243 1241
rect 14458 1232 14464 1284
rect 14516 1272 14522 1284
rect 15841 1275 15899 1281
rect 15841 1272 15853 1275
rect 14516 1244 15853 1272
rect 14516 1232 14522 1244
rect 15841 1241 15853 1244
rect 15887 1241 15899 1275
rect 15841 1235 15899 1241
rect 16206 1232 16212 1284
rect 16264 1272 16270 1284
rect 16761 1275 16819 1281
rect 16761 1272 16773 1275
rect 16264 1244 16773 1272
rect 16264 1232 16270 1244
rect 16761 1241 16773 1244
rect 16807 1241 16819 1275
rect 16761 1235 16819 1241
rect 19245 1275 19303 1281
rect 19245 1241 19257 1275
rect 19291 1272 19303 1275
rect 20990 1272 20996 1284
rect 19291 1244 20996 1272
rect 19291 1241 19303 1244
rect 19245 1235 19303 1241
rect 20990 1232 20996 1244
rect 21048 1232 21054 1284
rect 21174 1232 21180 1284
rect 21232 1232 21238 1284
rect 21910 1232 21916 1284
rect 21968 1232 21974 1284
rect 22094 1232 22100 1284
rect 22152 1232 22158 1284
rect 22204 1272 22232 1303
rect 22462 1300 22468 1352
rect 22520 1300 22526 1352
rect 23750 1300 23756 1352
rect 23808 1300 23814 1352
rect 24213 1343 24271 1349
rect 24213 1309 24225 1343
rect 24259 1340 24271 1343
rect 25056 1340 25084 1368
rect 24259 1312 25084 1340
rect 24259 1309 24271 1312
rect 24213 1303 24271 1309
rect 22922 1272 22928 1284
rect 22204 1244 22928 1272
rect 22922 1232 22928 1244
rect 22980 1232 22986 1284
rect 13633 1207 13691 1213
rect 13633 1173 13645 1207
rect 13679 1173 13691 1207
rect 13633 1167 13691 1173
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 14829 1167 14887 1173
rect 19061 1207 19119 1213
rect 19061 1173 19073 1207
rect 19107 1204 19119 1207
rect 21082 1204 21088 1216
rect 19107 1176 21088 1204
rect 19107 1173 19119 1176
rect 19061 1167 19119 1173
rect 21082 1164 21088 1176
rect 21140 1164 21146 1216
rect 21266 1164 21272 1216
rect 21324 1164 21330 1216
rect 21637 1207 21695 1213
rect 21637 1173 21649 1207
rect 21683 1204 21695 1207
rect 22186 1204 22192 1216
rect 21683 1176 22192 1204
rect 21683 1173 21695 1176
rect 21637 1167 21695 1173
rect 22186 1164 22192 1176
rect 22244 1164 22250 1216
rect 22373 1207 22431 1213
rect 22373 1173 22385 1207
rect 22419 1204 22431 1207
rect 23768 1204 23796 1300
rect 22419 1176 23796 1204
rect 22419 1173 22431 1176
rect 22373 1167 22431 1173
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 566 960 572 1012
rect 624 1000 630 1012
rect 2774 1000 2780 1012
rect 624 972 2780 1000
rect 624 960 630 972
rect 2774 960 2780 972
rect 2832 960 2838 1012
rect 3418 960 3424 1012
rect 3476 1000 3482 1012
rect 6270 1000 6276 1012
rect 3476 972 6276 1000
rect 3476 960 3482 972
rect 6270 960 6276 972
rect 6328 960 6334 1012
rect 9950 960 9956 1012
rect 10008 1000 10014 1012
rect 12526 1000 12532 1012
rect 10008 972 12532 1000
rect 10008 960 10014 972
rect 12526 960 12532 972
rect 12584 960 12590 1012
rect 21174 960 21180 1012
rect 21232 1000 21238 1012
rect 25590 1000 25596 1012
rect 21232 972 25596 1000
rect 21232 960 21238 972
rect 25590 960 25596 972
rect 25648 960 25654 1012
rect 9766 892 9772 944
rect 9824 932 9830 944
rect 11054 932 11060 944
rect 9824 904 11060 932
rect 9824 892 9830 904
rect 11054 892 11060 904
rect 11112 892 11118 944
rect 12250 892 12256 944
rect 12308 892 12314 944
rect 21082 892 21088 944
rect 21140 932 21146 944
rect 24210 932 24216 944
rect 21140 904 24216 932
rect 21140 892 21146 904
rect 24210 892 24216 904
rect 24268 892 24274 944
rect 5166 824 5172 876
rect 5224 864 5230 876
rect 12268 864 12296 892
rect 5224 836 12296 864
rect 5224 824 5230 836
rect 21266 824 21272 876
rect 21324 864 21330 876
rect 25498 864 25504 876
rect 21324 836 25504 864
rect 21324 824 21330 836
rect 25498 824 25504 836
rect 25556 824 25562 876
rect 7466 756 7472 808
rect 7524 796 7530 808
rect 14182 796 14188 808
rect 7524 768 14188 796
rect 7524 756 7530 768
rect 14182 756 14188 768
rect 14240 756 14246 808
rect 22094 756 22100 808
rect 22152 796 22158 808
rect 25222 796 25228 808
rect 22152 768 25228 796
rect 22152 756 22158 768
rect 25222 756 25228 768
rect 25280 756 25286 808
rect 1394 688 1400 740
rect 1452 728 1458 740
rect 2406 728 2412 740
rect 1452 700 2412 728
rect 1452 688 1458 700
rect 2406 688 2412 700
rect 2464 688 2470 740
rect 10318 688 10324 740
rect 10376 728 10382 740
rect 11330 728 11336 740
rect 10376 700 11336 728
rect 10376 688 10382 700
rect 11330 688 11336 700
rect 11388 688 11394 740
rect 20530 688 20536 740
rect 20588 728 20594 740
rect 23198 728 23204 740
rect 20588 700 23204 728
rect 20588 688 20594 700
rect 23198 688 23204 700
rect 23256 688 23262 740
rect 11238 620 11244 672
rect 11296 660 11302 672
rect 12066 660 12072 672
rect 11296 632 12072 660
rect 11296 620 11302 632
rect 12066 620 12072 632
rect 12124 620 12130 672
rect 20990 620 20996 672
rect 21048 660 21054 672
rect 22002 660 22008 672
rect 21048 632 22008 660
rect 21048 620 21054 632
rect 22002 620 22008 632
rect 22060 620 22066 672
rect 21910 552 21916 604
rect 21968 592 21974 604
rect 23750 592 23756 604
rect 21968 564 23756 592
rect 21968 552 21974 564
rect 23750 552 23756 564
rect 23808 552 23814 604
rect 18046 484 18052 536
rect 18104 524 18110 536
rect 24210 524 24216 536
rect 18104 496 24216 524
rect 18104 484 18110 496
rect 24210 484 24216 496
rect 24268 484 24274 536
rect 21174 416 21180 468
rect 21232 456 21238 468
rect 22462 456 22468 468
rect 21232 428 22468 456
rect 21232 416 21238 428
rect 22462 416 22468 428
rect 22520 416 22526 468
rect 8386 76 8392 128
rect 8444 116 8450 128
rect 9398 116 9404 128
rect 8444 88 9404 116
rect 8444 76 8450 88
rect 9398 76 9404 88
rect 9456 76 9462 128
<< via1 >>
rect 18604 43800 18656 43852
rect 20720 43800 20772 43852
rect 19432 43732 19484 43784
rect 19800 43732 19852 43784
rect 15292 43664 15344 43716
rect 5356 43596 5408 43648
rect 10508 43596 10560 43648
rect 17500 43596 17552 43648
rect 21272 43596 21324 43648
rect 24400 43596 24452 43648
rect 6884 43494 6936 43546
rect 6948 43494 7000 43546
rect 7012 43494 7064 43546
rect 7076 43494 7128 43546
rect 7140 43494 7192 43546
rect 12818 43494 12870 43546
rect 12882 43494 12934 43546
rect 12946 43494 12998 43546
rect 13010 43494 13062 43546
rect 13074 43494 13126 43546
rect 18752 43494 18804 43546
rect 18816 43494 18868 43546
rect 18880 43494 18932 43546
rect 18944 43494 18996 43546
rect 19008 43494 19060 43546
rect 24686 43494 24738 43546
rect 24750 43494 24802 43546
rect 24814 43494 24866 43546
rect 24878 43494 24930 43546
rect 24942 43494 24994 43546
rect 1860 43435 1912 43444
rect 1860 43401 1869 43435
rect 1869 43401 1903 43435
rect 1903 43401 1912 43435
rect 1860 43392 1912 43401
rect 2964 43392 3016 43444
rect 388 43324 440 43376
rect 4344 43392 4396 43444
rect 5540 43435 5592 43444
rect 5540 43401 5549 43435
rect 5549 43401 5583 43435
rect 5583 43401 5592 43435
rect 5540 43392 5592 43401
rect 6276 43392 6328 43444
rect 3424 43324 3476 43376
rect 6828 43435 6880 43444
rect 6828 43401 6837 43435
rect 6837 43401 6871 43435
rect 6871 43401 6880 43435
rect 6828 43392 6880 43401
rect 7656 43392 7708 43444
rect 7932 43392 7984 43444
rect 8484 43392 8536 43444
rect 9036 43392 9088 43444
rect 9588 43392 9640 43444
rect 9864 43392 9916 43444
rect 10508 43435 10560 43444
rect 10508 43401 10517 43435
rect 10517 43401 10551 43435
rect 10551 43401 10560 43435
rect 10508 43392 10560 43401
rect 13360 43392 13412 43444
rect 8576 43324 8628 43376
rect 1216 43256 1268 43308
rect 1768 43299 1820 43308
rect 1768 43265 1777 43299
rect 1777 43265 1811 43299
rect 1811 43265 1820 43299
rect 1768 43256 1820 43265
rect 2504 43299 2556 43308
rect 2504 43265 2513 43299
rect 2513 43265 2547 43299
rect 2547 43265 2556 43299
rect 2504 43256 2556 43265
rect 3056 43299 3108 43308
rect 3056 43265 3065 43299
rect 3065 43265 3099 43299
rect 3099 43265 3108 43299
rect 3056 43256 3108 43265
rect 5264 43299 5316 43308
rect 5264 43265 5273 43299
rect 5273 43265 5307 43299
rect 5307 43265 5316 43299
rect 5264 43256 5316 43265
rect 6000 43256 6052 43308
rect 6276 43256 6328 43308
rect 7288 43256 7340 43308
rect 8116 43256 8168 43308
rect 9404 43324 9456 43376
rect 4804 43188 4856 43240
rect 9956 43299 10008 43308
rect 9956 43265 9965 43299
rect 9965 43265 9999 43299
rect 9999 43265 10008 43299
rect 9956 43256 10008 43265
rect 10324 43299 10376 43308
rect 10324 43265 10333 43299
rect 10333 43265 10367 43299
rect 10367 43265 10376 43299
rect 10324 43256 10376 43265
rect 10692 43299 10744 43308
rect 10692 43265 10701 43299
rect 10701 43265 10735 43299
rect 10735 43265 10744 43299
rect 10692 43256 10744 43265
rect 11060 43299 11112 43308
rect 11060 43265 11069 43299
rect 11069 43265 11103 43299
rect 11103 43265 11112 43299
rect 11060 43256 11112 43265
rect 11244 43256 11296 43308
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 12440 43367 12492 43376
rect 12440 43333 12449 43367
rect 12449 43333 12483 43367
rect 12483 43333 12492 43367
rect 12440 43324 12492 43333
rect 12808 43367 12860 43376
rect 12808 43333 12817 43367
rect 12817 43333 12851 43367
rect 12851 43333 12860 43367
rect 12808 43324 12860 43333
rect 13452 43324 13504 43376
rect 15292 43392 15344 43444
rect 17040 43392 17092 43444
rect 14740 43367 14792 43376
rect 14740 43333 14749 43367
rect 14749 43333 14783 43367
rect 14783 43333 14792 43367
rect 14740 43324 14792 43333
rect 14832 43324 14884 43376
rect 15568 43367 15620 43376
rect 15568 43333 15577 43367
rect 15577 43333 15611 43367
rect 15611 43333 15620 43367
rect 15568 43324 15620 43333
rect 15936 43324 15988 43376
rect 16396 43324 16448 43376
rect 16856 43324 16908 43376
rect 13636 43256 13688 43308
rect 15844 43299 15896 43308
rect 15844 43265 15853 43299
rect 15853 43265 15887 43299
rect 15887 43265 15896 43299
rect 15844 43256 15896 43265
rect 9680 43188 9732 43240
rect 4712 43120 4764 43172
rect 9128 43120 9180 43172
rect 14924 43163 14976 43172
rect 14924 43129 14933 43163
rect 14933 43129 14967 43163
rect 14967 43129 14976 43163
rect 14924 43120 14976 43129
rect 15568 43120 15620 43172
rect 1676 43052 1728 43104
rect 3608 43052 3660 43104
rect 4436 43052 4488 43104
rect 9404 43052 9456 43104
rect 10600 43052 10652 43104
rect 10876 43095 10928 43104
rect 10876 43061 10885 43095
rect 10885 43061 10919 43095
rect 10919 43061 10928 43095
rect 10876 43052 10928 43061
rect 11244 43095 11296 43104
rect 11244 43061 11253 43095
rect 11253 43061 11287 43095
rect 11287 43061 11296 43095
rect 11244 43052 11296 43061
rect 11704 43095 11756 43104
rect 11704 43061 11713 43095
rect 11713 43061 11747 43095
rect 11747 43061 11756 43095
rect 11704 43052 11756 43061
rect 12256 43095 12308 43104
rect 12256 43061 12265 43095
rect 12265 43061 12299 43095
rect 12299 43061 12308 43095
rect 12256 43052 12308 43061
rect 12532 43095 12584 43104
rect 12532 43061 12541 43095
rect 12541 43061 12575 43095
rect 12575 43061 12584 43095
rect 12532 43052 12584 43061
rect 12624 43052 12676 43104
rect 13820 43095 13872 43104
rect 13820 43061 13829 43095
rect 13829 43061 13863 43095
rect 13863 43061 13872 43095
rect 13820 43052 13872 43061
rect 14280 43095 14332 43104
rect 14280 43061 14289 43095
rect 14289 43061 14323 43095
rect 14323 43061 14332 43095
rect 14280 43052 14332 43061
rect 14740 43052 14792 43104
rect 15660 43095 15712 43104
rect 15660 43061 15669 43095
rect 15669 43061 15703 43095
rect 15703 43061 15712 43095
rect 15660 43052 15712 43061
rect 16304 43120 16356 43172
rect 18144 43392 18196 43444
rect 18236 43324 18288 43376
rect 17408 43188 17460 43240
rect 19340 43256 19392 43308
rect 20352 43392 20404 43444
rect 20628 43392 20680 43444
rect 21180 43392 21232 43444
rect 19984 43324 20036 43376
rect 19708 43299 19760 43308
rect 19708 43265 19717 43299
rect 19717 43265 19751 43299
rect 19751 43265 19760 43299
rect 19708 43256 19760 43265
rect 19892 43299 19944 43308
rect 19892 43265 19901 43299
rect 19901 43265 19935 43299
rect 19935 43265 19944 43299
rect 19892 43256 19944 43265
rect 17776 43120 17828 43172
rect 18236 43120 18288 43172
rect 19156 43120 19208 43172
rect 19708 43120 19760 43172
rect 16856 43095 16908 43104
rect 16856 43061 16865 43095
rect 16865 43061 16899 43095
rect 16899 43061 16908 43095
rect 16856 43052 16908 43061
rect 17500 43052 17552 43104
rect 17592 43095 17644 43104
rect 17592 43061 17601 43095
rect 17601 43061 17635 43095
rect 17635 43061 17644 43095
rect 17592 43052 17644 43061
rect 17868 43095 17920 43104
rect 17868 43061 17877 43095
rect 17877 43061 17911 43095
rect 17911 43061 17920 43095
rect 17868 43052 17920 43061
rect 18052 43052 18104 43104
rect 18604 43052 18656 43104
rect 19524 43095 19576 43104
rect 19524 43061 19533 43095
rect 19533 43061 19567 43095
rect 19567 43061 19576 43095
rect 19524 43052 19576 43061
rect 20444 43256 20496 43308
rect 21548 43324 21600 43376
rect 23112 43392 23164 43444
rect 21640 43256 21692 43308
rect 22376 43256 22428 43308
rect 22652 43256 22704 43308
rect 22560 43188 22612 43240
rect 20904 43120 20956 43172
rect 22192 43120 22244 43172
rect 23480 43256 23532 43308
rect 21364 43052 21416 43104
rect 21916 43052 21968 43104
rect 24124 43095 24176 43104
rect 24124 43061 24133 43095
rect 24133 43061 24167 43095
rect 24167 43061 24176 43095
rect 24124 43052 24176 43061
rect 3917 42950 3969 43002
rect 3981 42950 4033 43002
rect 4045 42950 4097 43002
rect 4109 42950 4161 43002
rect 4173 42950 4225 43002
rect 9851 42950 9903 43002
rect 9915 42950 9967 43002
rect 9979 42950 10031 43002
rect 10043 42950 10095 43002
rect 10107 42950 10159 43002
rect 15785 42950 15837 43002
rect 15849 42950 15901 43002
rect 15913 42950 15965 43002
rect 15977 42950 16029 43002
rect 16041 42950 16093 43002
rect 21719 42950 21771 43002
rect 21783 42950 21835 43002
rect 21847 42950 21899 43002
rect 21911 42950 21963 43002
rect 21975 42950 22027 43002
rect 2228 42891 2280 42900
rect 2228 42857 2237 42891
rect 2237 42857 2271 42891
rect 2271 42857 2280 42891
rect 2228 42848 2280 42857
rect 3332 42891 3384 42900
rect 3332 42857 3341 42891
rect 3341 42857 3375 42891
rect 3375 42857 3384 42891
rect 3332 42848 3384 42857
rect 6092 42891 6144 42900
rect 6092 42857 6101 42891
rect 6101 42857 6135 42891
rect 6135 42857 6144 42891
rect 6092 42848 6144 42857
rect 6828 42891 6880 42900
rect 6828 42857 6837 42891
rect 6837 42857 6871 42891
rect 6871 42857 6880 42891
rect 6828 42848 6880 42857
rect 7380 42891 7432 42900
rect 7380 42857 7389 42891
rect 7389 42857 7423 42891
rect 7423 42857 7432 42891
rect 7380 42848 7432 42857
rect 1400 42712 1452 42764
rect 20 42644 72 42696
rect 3700 42712 3752 42764
rect 4344 42755 4396 42764
rect 4344 42721 4353 42755
rect 4353 42721 4387 42755
rect 4387 42721 4396 42755
rect 4344 42712 4396 42721
rect 4896 42712 4948 42764
rect 5540 42780 5592 42832
rect 9128 42848 9180 42900
rect 9680 42848 9732 42900
rect 10600 42891 10652 42900
rect 10600 42857 10609 42891
rect 10609 42857 10643 42891
rect 10643 42857 10652 42891
rect 10600 42848 10652 42857
rect 9220 42780 9272 42832
rect 16856 42848 16908 42900
rect 17868 42848 17920 42900
rect 18144 42848 18196 42900
rect 8484 42712 8536 42764
rect 8760 42712 8812 42764
rect 9312 42712 9364 42764
rect 4252 42644 4304 42696
rect 4712 42644 4764 42696
rect 5540 42687 5592 42696
rect 5540 42653 5549 42687
rect 5549 42653 5583 42687
rect 5583 42653 5592 42687
rect 5540 42644 5592 42653
rect 7564 42644 7616 42696
rect 8392 42687 8444 42696
rect 8392 42653 8401 42687
rect 8401 42653 8435 42687
rect 8435 42653 8444 42687
rect 8392 42644 8444 42653
rect 9036 42644 9088 42696
rect 9404 42644 9456 42696
rect 9956 42644 10008 42696
rect 12256 42712 12308 42764
rect 12440 42712 12492 42764
rect 14740 42780 14792 42832
rect 17132 42780 17184 42832
rect 13820 42712 13872 42764
rect 2320 42576 2372 42628
rect 2872 42576 2924 42628
rect 3240 42619 3292 42628
rect 3240 42585 3249 42619
rect 3249 42585 3283 42619
rect 3283 42585 3292 42619
rect 3240 42576 3292 42585
rect 4436 42576 4488 42628
rect 6000 42619 6052 42628
rect 6000 42585 6009 42619
rect 6009 42585 6043 42619
rect 6043 42585 6052 42619
rect 6000 42576 6052 42585
rect 2780 42551 2832 42560
rect 2780 42517 2789 42551
rect 2789 42517 2823 42551
rect 2823 42517 2832 42551
rect 2780 42508 2832 42517
rect 4620 42508 4672 42560
rect 5724 42551 5776 42560
rect 5724 42517 5733 42551
rect 5733 42517 5767 42551
rect 5767 42517 5776 42551
rect 5724 42508 5776 42517
rect 5908 42508 5960 42560
rect 7288 42619 7340 42628
rect 7288 42585 7297 42619
rect 7297 42585 7331 42619
rect 7331 42585 7340 42619
rect 7288 42576 7340 42585
rect 7472 42508 7524 42560
rect 9588 42576 9640 42628
rect 10416 42576 10468 42628
rect 11612 42687 11664 42696
rect 11612 42653 11621 42687
rect 11621 42653 11655 42687
rect 11655 42653 11664 42687
rect 11612 42644 11664 42653
rect 11888 42687 11940 42696
rect 11888 42653 11897 42687
rect 11897 42653 11931 42687
rect 11931 42653 11940 42687
rect 11888 42644 11940 42653
rect 11336 42576 11388 42628
rect 12992 42687 13044 42696
rect 12992 42653 13001 42687
rect 13001 42653 13035 42687
rect 13035 42653 13044 42687
rect 12992 42644 13044 42653
rect 14096 42687 14148 42696
rect 14096 42653 14105 42687
rect 14105 42653 14139 42687
rect 14139 42653 14148 42687
rect 14096 42644 14148 42653
rect 14372 42687 14424 42696
rect 14372 42653 14381 42687
rect 14381 42653 14415 42687
rect 14415 42653 14424 42687
rect 14372 42644 14424 42653
rect 15200 42712 15252 42764
rect 18328 42780 18380 42832
rect 15292 42687 15344 42696
rect 15292 42653 15301 42687
rect 15301 42653 15335 42687
rect 15335 42653 15344 42687
rect 15292 42644 15344 42653
rect 16488 42687 16540 42696
rect 16488 42653 16497 42687
rect 16497 42653 16531 42687
rect 16531 42653 16540 42687
rect 16488 42644 16540 42653
rect 16580 42687 16632 42696
rect 16580 42653 16589 42687
rect 16589 42653 16623 42687
rect 16623 42653 16632 42687
rect 16580 42644 16632 42653
rect 9128 42508 9180 42560
rect 11796 42551 11848 42560
rect 11796 42517 11805 42551
rect 11805 42517 11839 42551
rect 11839 42517 11848 42551
rect 11796 42508 11848 42517
rect 13268 42576 13320 42628
rect 14740 42576 14792 42628
rect 17592 42644 17644 42696
rect 17776 42644 17828 42696
rect 18052 42644 18104 42696
rect 18604 42712 18656 42764
rect 18788 42683 18840 42696
rect 18788 42649 18797 42683
rect 18797 42649 18831 42683
rect 18831 42649 18840 42683
rect 18788 42644 18840 42649
rect 19064 42687 19116 42696
rect 19064 42653 19073 42687
rect 19073 42653 19107 42687
rect 19107 42653 19116 42687
rect 19064 42644 19116 42653
rect 21272 42780 21324 42832
rect 12164 42508 12216 42560
rect 13452 42508 13504 42560
rect 14556 42551 14608 42560
rect 14556 42517 14565 42551
rect 14565 42517 14599 42551
rect 14599 42517 14608 42551
rect 14556 42508 14608 42517
rect 14832 42551 14884 42560
rect 14832 42517 14841 42551
rect 14841 42517 14875 42551
rect 14875 42517 14884 42551
rect 14832 42508 14884 42517
rect 15476 42551 15528 42560
rect 15476 42517 15485 42551
rect 15485 42517 15519 42551
rect 15519 42517 15528 42551
rect 15476 42508 15528 42517
rect 19248 42619 19300 42628
rect 19248 42585 19257 42619
rect 19257 42585 19291 42619
rect 19291 42585 19300 42619
rect 19248 42576 19300 42585
rect 15844 42508 15896 42560
rect 16764 42551 16816 42560
rect 16764 42517 16773 42551
rect 16773 42517 16807 42551
rect 16807 42517 16816 42551
rect 16764 42508 16816 42517
rect 16948 42551 17000 42560
rect 16948 42517 16957 42551
rect 16957 42517 16991 42551
rect 16991 42517 17000 42551
rect 16948 42508 17000 42517
rect 17224 42551 17276 42560
rect 17224 42517 17233 42551
rect 17233 42517 17267 42551
rect 17267 42517 17276 42551
rect 17224 42508 17276 42517
rect 17316 42508 17368 42560
rect 17776 42551 17828 42560
rect 17776 42517 17785 42551
rect 17785 42517 17819 42551
rect 17819 42517 17828 42551
rect 17776 42508 17828 42517
rect 18052 42551 18104 42560
rect 18052 42517 18061 42551
rect 18061 42517 18095 42551
rect 18095 42517 18104 42551
rect 18052 42508 18104 42517
rect 18328 42551 18380 42560
rect 18328 42517 18337 42551
rect 18337 42517 18371 42551
rect 18371 42517 18380 42551
rect 18328 42508 18380 42517
rect 18604 42551 18656 42560
rect 18604 42517 18613 42551
rect 18613 42517 18647 42551
rect 18647 42517 18656 42551
rect 18604 42508 18656 42517
rect 18972 42508 19024 42560
rect 20812 42576 20864 42628
rect 21088 42576 21140 42628
rect 21548 42619 21600 42628
rect 21548 42585 21557 42619
rect 21557 42585 21591 42619
rect 21591 42585 21600 42619
rect 21548 42576 21600 42585
rect 21916 42687 21968 42696
rect 21916 42653 21925 42687
rect 21925 42653 21959 42687
rect 21959 42653 21968 42687
rect 21916 42644 21968 42653
rect 22376 42780 22428 42832
rect 23020 42780 23072 42832
rect 22284 42712 22336 42764
rect 25136 42712 25188 42764
rect 20536 42551 20588 42560
rect 20536 42517 20545 42551
rect 20545 42517 20579 42551
rect 20579 42517 20588 42551
rect 20536 42508 20588 42517
rect 20996 42508 21048 42560
rect 21916 42508 21968 42560
rect 22192 42508 22244 42560
rect 23756 42619 23808 42628
rect 23756 42585 23765 42619
rect 23765 42585 23799 42619
rect 23799 42585 23808 42619
rect 23756 42576 23808 42585
rect 24216 42644 24268 42696
rect 24584 42644 24636 42696
rect 6884 42406 6936 42458
rect 6948 42406 7000 42458
rect 7012 42406 7064 42458
rect 7076 42406 7128 42458
rect 7140 42406 7192 42458
rect 12818 42406 12870 42458
rect 12882 42406 12934 42458
rect 12946 42406 12998 42458
rect 13010 42406 13062 42458
rect 13074 42406 13126 42458
rect 18752 42406 18804 42458
rect 18816 42406 18868 42458
rect 18880 42406 18932 42458
rect 18944 42406 18996 42458
rect 19008 42406 19060 42458
rect 24686 42406 24738 42458
rect 24750 42406 24802 42458
rect 24814 42406 24866 42458
rect 24878 42406 24930 42458
rect 24942 42406 24994 42458
rect 480 42304 532 42356
rect 1768 42304 1820 42356
rect 3240 42304 3292 42356
rect 3608 42304 3660 42356
rect 2412 42168 2464 42220
rect 2780 42211 2832 42220
rect 2780 42177 2789 42211
rect 2789 42177 2823 42211
rect 2823 42177 2832 42211
rect 2780 42168 2832 42177
rect 3792 42304 3844 42356
rect 3884 42211 3936 42220
rect 3884 42177 3893 42211
rect 3893 42177 3927 42211
rect 3927 42177 3936 42211
rect 3884 42168 3936 42177
rect 1216 41964 1268 42016
rect 3148 42100 3200 42152
rect 3516 42032 3568 42084
rect 3608 42032 3660 42084
rect 4712 42211 4764 42220
rect 4712 42177 4721 42211
rect 4721 42177 4755 42211
rect 4755 42177 4764 42211
rect 4712 42168 4764 42177
rect 5172 42304 5224 42356
rect 6276 42304 6328 42356
rect 7012 42304 7064 42356
rect 7380 42304 7432 42356
rect 8208 42304 8260 42356
rect 8576 42304 8628 42356
rect 9128 42304 9180 42356
rect 9496 42304 9548 42356
rect 9956 42347 10008 42356
rect 9956 42313 9965 42347
rect 9965 42313 9999 42347
rect 9999 42313 10008 42347
rect 9956 42304 10008 42313
rect 15476 42304 15528 42356
rect 5080 42032 5132 42084
rect 5724 42168 5776 42220
rect 6184 42211 6236 42220
rect 6184 42177 6193 42211
rect 6193 42177 6227 42211
rect 6227 42177 6236 42211
rect 6184 42168 6236 42177
rect 6552 42211 6604 42220
rect 6552 42177 6561 42211
rect 6561 42177 6595 42211
rect 6595 42177 6604 42211
rect 6552 42168 6604 42177
rect 7380 42211 7432 42220
rect 7380 42177 7389 42211
rect 7389 42177 7423 42211
rect 7423 42177 7432 42211
rect 7380 42168 7432 42177
rect 7656 42211 7708 42220
rect 7656 42177 7665 42211
rect 7665 42177 7699 42211
rect 7699 42177 7708 42211
rect 7656 42168 7708 42177
rect 7932 42211 7984 42220
rect 7932 42177 7941 42211
rect 7941 42177 7975 42211
rect 7975 42177 7984 42211
rect 7932 42168 7984 42177
rect 8208 42211 8260 42220
rect 8208 42177 8217 42211
rect 8217 42177 8251 42211
rect 8251 42177 8260 42211
rect 8208 42168 8260 42177
rect 7196 42100 7248 42152
rect 7840 42100 7892 42152
rect 9128 42211 9180 42220
rect 9128 42177 9137 42211
rect 9137 42177 9171 42211
rect 9171 42177 9180 42211
rect 9128 42168 9180 42177
rect 9404 42211 9456 42220
rect 9404 42177 9413 42211
rect 9413 42177 9447 42211
rect 9447 42177 9456 42211
rect 9404 42168 9456 42177
rect 13636 42236 13688 42288
rect 15844 42236 15896 42288
rect 17224 42304 17276 42356
rect 17316 42304 17368 42356
rect 17776 42304 17828 42356
rect 18052 42304 18104 42356
rect 16948 42236 17000 42288
rect 18144 42236 18196 42288
rect 18328 42304 18380 42356
rect 19064 42304 19116 42356
rect 19432 42304 19484 42356
rect 18604 42279 18656 42288
rect 18604 42245 18613 42279
rect 18613 42245 18647 42279
rect 18647 42245 18656 42279
rect 18604 42236 18656 42245
rect 9864 42211 9916 42220
rect 9864 42177 9873 42211
rect 9873 42177 9907 42211
rect 9907 42177 9916 42211
rect 9864 42168 9916 42177
rect 9496 42100 9548 42152
rect 5632 42032 5684 42084
rect 6460 42032 6512 42084
rect 5724 42007 5776 42016
rect 5724 41973 5733 42007
rect 5733 41973 5767 42007
rect 5767 41973 5776 42007
rect 5724 41964 5776 41973
rect 6920 42007 6972 42016
rect 6920 41973 6929 42007
rect 6929 41973 6963 42007
rect 6963 41973 6972 42007
rect 6920 41964 6972 41973
rect 7380 41964 7432 42016
rect 7472 42007 7524 42016
rect 7472 41973 7481 42007
rect 7481 41973 7515 42007
rect 7515 41973 7524 42007
rect 7472 41964 7524 41973
rect 7748 42007 7800 42016
rect 7748 41973 7757 42007
rect 7757 41973 7791 42007
rect 7791 41973 7800 42007
rect 7748 41964 7800 41973
rect 8024 42007 8076 42016
rect 8024 41973 8033 42007
rect 8033 41973 8067 42007
rect 8067 41973 8076 42007
rect 8024 41964 8076 41973
rect 8300 42032 8352 42084
rect 12164 42168 12216 42220
rect 19524 42236 19576 42288
rect 18880 42168 18932 42220
rect 20812 42347 20864 42356
rect 20812 42313 20821 42347
rect 20821 42313 20855 42347
rect 20855 42313 20864 42347
rect 20812 42304 20864 42313
rect 21640 42304 21692 42356
rect 22836 42304 22888 42356
rect 23204 42304 23256 42356
rect 24492 42304 24544 42356
rect 15292 42032 15344 42084
rect 16120 42032 16172 42084
rect 16396 42075 16448 42084
rect 16396 42041 16405 42075
rect 16405 42041 16439 42075
rect 16439 42041 16448 42075
rect 16396 42032 16448 42041
rect 17316 42075 17368 42084
rect 17316 42041 17325 42075
rect 17325 42041 17359 42075
rect 17359 42041 17368 42075
rect 17316 42032 17368 42041
rect 18420 42075 18472 42084
rect 18420 42041 18429 42075
rect 18429 42041 18463 42075
rect 18463 42041 18472 42075
rect 18420 42032 18472 42041
rect 15200 41964 15252 42016
rect 15384 41964 15436 42016
rect 16488 41964 16540 42016
rect 16856 42007 16908 42016
rect 16856 41973 16865 42007
rect 16865 41973 16899 42007
rect 16899 41973 16908 42007
rect 16856 41964 16908 41973
rect 17592 42007 17644 42016
rect 17592 41973 17601 42007
rect 17601 41973 17635 42007
rect 17635 41973 17644 42007
rect 17592 41964 17644 41973
rect 18144 41964 18196 42016
rect 18972 42032 19024 42084
rect 19892 42032 19944 42084
rect 20260 42100 20312 42152
rect 20812 42168 20864 42220
rect 21272 42211 21324 42220
rect 21272 42177 21281 42211
rect 21281 42177 21315 42211
rect 21315 42177 21324 42211
rect 21272 42168 21324 42177
rect 20904 42100 20956 42152
rect 22192 42168 22244 42220
rect 18696 42007 18748 42016
rect 18696 41973 18705 42007
rect 18705 41973 18739 42007
rect 18739 41973 18748 42007
rect 18696 41964 18748 41973
rect 18788 41964 18840 42016
rect 19432 42007 19484 42016
rect 19432 41973 19441 42007
rect 19441 41973 19475 42007
rect 19475 41973 19484 42007
rect 19432 41964 19484 41973
rect 20444 42032 20496 42084
rect 21916 42032 21968 42084
rect 22008 42032 22060 42084
rect 22836 42211 22888 42220
rect 22836 42177 22845 42211
rect 22845 42177 22879 42211
rect 22879 42177 22888 42211
rect 22836 42168 22888 42177
rect 24584 42236 24636 42288
rect 24032 42211 24084 42220
rect 24032 42177 24041 42211
rect 24041 42177 24075 42211
rect 24075 42177 24084 42211
rect 24032 42168 24084 42177
rect 25596 42100 25648 42152
rect 24216 42032 24268 42084
rect 21180 41964 21232 42016
rect 23480 41964 23532 42016
rect 25228 41964 25280 42016
rect 3917 41862 3969 41914
rect 3981 41862 4033 41914
rect 4045 41862 4097 41914
rect 4109 41862 4161 41914
rect 4173 41862 4225 41914
rect 9851 41862 9903 41914
rect 9915 41862 9967 41914
rect 9979 41862 10031 41914
rect 10043 41862 10095 41914
rect 10107 41862 10159 41914
rect 15785 41862 15837 41914
rect 15849 41862 15901 41914
rect 15913 41862 15965 41914
rect 15977 41862 16029 41914
rect 16041 41862 16093 41914
rect 21719 41862 21771 41914
rect 21783 41862 21835 41914
rect 21847 41862 21899 41914
rect 21911 41862 21963 41914
rect 21975 41862 22027 41914
rect 940 41760 992 41812
rect 2596 41760 2648 41812
rect 2780 41760 2832 41812
rect 3332 41760 3384 41812
rect 3608 41760 3660 41812
rect 4252 41760 4304 41812
rect 4436 41803 4488 41812
rect 4436 41769 4445 41803
rect 4445 41769 4479 41803
rect 4479 41769 4488 41803
rect 4436 41760 4488 41769
rect 5264 41760 5316 41812
rect 5540 41760 5592 41812
rect 5908 41760 5960 41812
rect 6000 41760 6052 41812
rect 6920 41760 6972 41812
rect 7288 41760 7340 41812
rect 7380 41760 7432 41812
rect 7472 41760 7524 41812
rect 7564 41803 7616 41812
rect 7564 41769 7573 41803
rect 7573 41769 7607 41803
rect 7607 41769 7616 41803
rect 7564 41760 7616 41769
rect 7748 41760 7800 41812
rect 3792 41624 3844 41676
rect 4988 41624 5040 41676
rect 5080 41624 5132 41676
rect 1492 41599 1544 41608
rect 1492 41565 1501 41599
rect 1501 41565 1535 41599
rect 1535 41565 1544 41599
rect 1492 41556 1544 41565
rect 1676 41488 1728 41540
rect 2320 41488 2372 41540
rect 2964 41488 3016 41540
rect 3332 41599 3384 41608
rect 3332 41565 3341 41599
rect 3341 41565 3375 41599
rect 3375 41565 3384 41599
rect 3332 41556 3384 41565
rect 3608 41599 3660 41608
rect 3608 41565 3617 41599
rect 3617 41565 3651 41599
rect 3651 41565 3660 41599
rect 3608 41556 3660 41565
rect 3700 41556 3752 41608
rect 4252 41599 4304 41608
rect 4252 41565 4261 41599
rect 4261 41565 4295 41599
rect 4295 41565 4304 41599
rect 4252 41556 4304 41565
rect 4620 41599 4672 41608
rect 4620 41565 4629 41599
rect 4629 41565 4663 41599
rect 4663 41565 4672 41599
rect 4620 41556 4672 41565
rect 3424 41488 3476 41540
rect 4160 41488 4212 41540
rect 5632 41599 5684 41608
rect 5632 41565 5641 41599
rect 5641 41565 5675 41599
rect 5675 41565 5684 41599
rect 5632 41556 5684 41565
rect 5724 41556 5776 41608
rect 6736 41599 6788 41608
rect 6736 41565 6745 41599
rect 6745 41565 6779 41599
rect 6779 41565 6788 41599
rect 6736 41556 6788 41565
rect 8116 41735 8168 41744
rect 8116 41701 8125 41735
rect 8125 41701 8159 41735
rect 8159 41701 8168 41735
rect 8116 41692 8168 41701
rect 8484 41760 8536 41812
rect 10048 41760 10100 41812
rect 17960 41803 18012 41812
rect 17960 41769 17969 41803
rect 17969 41769 18003 41803
rect 18003 41769 18012 41803
rect 17960 41760 18012 41769
rect 18052 41760 18104 41812
rect 18512 41760 18564 41812
rect 18880 41760 18932 41812
rect 19524 41760 19576 41812
rect 20260 41803 20312 41812
rect 20260 41769 20269 41803
rect 20269 41769 20303 41803
rect 20303 41769 20312 41803
rect 20260 41760 20312 41769
rect 20536 41760 20588 41812
rect 20352 41692 20404 41744
rect 20720 41803 20772 41812
rect 20720 41769 20729 41803
rect 20729 41769 20763 41803
rect 20763 41769 20772 41803
rect 20720 41760 20772 41769
rect 21180 41803 21232 41812
rect 21180 41769 21189 41803
rect 21189 41769 21223 41803
rect 21223 41769 21232 41803
rect 21180 41760 21232 41769
rect 21364 41760 21416 41812
rect 22284 41760 22336 41812
rect 23940 41760 23992 41812
rect 25320 41760 25372 41812
rect 25412 41760 25464 41812
rect 8852 41556 8904 41608
rect 10324 41556 10376 41608
rect 17960 41556 18012 41608
rect 1584 41420 1636 41472
rect 6092 41420 6144 41472
rect 7012 41488 7064 41540
rect 7288 41420 7340 41472
rect 15476 41488 15528 41540
rect 17776 41488 17828 41540
rect 18144 41599 18196 41608
rect 18144 41565 18153 41599
rect 18153 41565 18187 41599
rect 18187 41565 18196 41599
rect 18144 41556 18196 41565
rect 18236 41556 18288 41608
rect 18420 41556 18472 41608
rect 19708 41556 19760 41608
rect 20260 41556 20312 41608
rect 19340 41488 19392 41540
rect 10692 41463 10744 41472
rect 10692 41429 10701 41463
rect 10701 41429 10735 41463
rect 10735 41429 10744 41463
rect 10692 41420 10744 41429
rect 15200 41420 15252 41472
rect 21180 41556 21232 41608
rect 21364 41599 21416 41608
rect 21364 41565 21373 41599
rect 21373 41565 21407 41599
rect 21407 41565 21416 41599
rect 21364 41556 21416 41565
rect 21640 41599 21692 41608
rect 21640 41565 21649 41599
rect 21649 41565 21683 41599
rect 21683 41565 21692 41599
rect 21640 41556 21692 41565
rect 21824 41488 21876 41540
rect 23572 41556 23624 41608
rect 25780 41556 25832 41608
rect 21456 41463 21508 41472
rect 21456 41429 21465 41463
rect 21465 41429 21499 41463
rect 21499 41429 21508 41463
rect 21456 41420 21508 41429
rect 22376 41420 22428 41472
rect 23664 41420 23716 41472
rect 23848 41531 23900 41540
rect 23848 41497 23857 41531
rect 23857 41497 23891 41531
rect 23891 41497 23900 41531
rect 23848 41488 23900 41497
rect 23940 41420 23992 41472
rect 6884 41318 6936 41370
rect 6948 41318 7000 41370
rect 7012 41318 7064 41370
rect 7076 41318 7128 41370
rect 7140 41318 7192 41370
rect 12818 41318 12870 41370
rect 12882 41318 12934 41370
rect 12946 41318 12998 41370
rect 13010 41318 13062 41370
rect 13074 41318 13126 41370
rect 18752 41318 18804 41370
rect 18816 41318 18868 41370
rect 18880 41318 18932 41370
rect 18944 41318 18996 41370
rect 19008 41318 19060 41370
rect 24686 41318 24738 41370
rect 24750 41318 24802 41370
rect 24814 41318 24866 41370
rect 24878 41318 24930 41370
rect 24942 41318 24994 41370
rect 2504 41259 2556 41268
rect 2504 41225 2513 41259
rect 2513 41225 2547 41259
rect 2547 41225 2556 41259
rect 2504 41216 2556 41225
rect 2780 41259 2832 41268
rect 2780 41225 2789 41259
rect 2789 41225 2823 41259
rect 2823 41225 2832 41259
rect 2780 41216 2832 41225
rect 2964 41216 3016 41268
rect 7840 41216 7892 41268
rect 15108 41216 15160 41268
rect 1400 41123 1452 41132
rect 1400 41089 1409 41123
rect 1409 41089 1443 41123
rect 1443 41089 1452 41123
rect 1400 41080 1452 41089
rect 480 41012 532 41064
rect 388 40944 440 40996
rect 3240 41123 3292 41132
rect 3240 41089 3249 41123
rect 3249 41089 3283 41123
rect 3283 41089 3292 41123
rect 3240 41080 3292 41089
rect 3424 41080 3476 41132
rect 3516 41055 3568 41064
rect 3516 41021 3525 41055
rect 3525 41021 3559 41055
rect 3559 41021 3568 41055
rect 3516 41012 3568 41021
rect 1032 40876 1084 40928
rect 3332 40876 3384 40928
rect 4528 40919 4580 40928
rect 4528 40885 4537 40919
rect 4537 40885 4571 40919
rect 4571 40885 4580 40919
rect 4528 40876 4580 40885
rect 5264 41080 5316 41132
rect 7932 41123 7984 41132
rect 7932 41089 7941 41123
rect 7941 41089 7975 41123
rect 7975 41089 7984 41123
rect 7932 41080 7984 41089
rect 12532 41148 12584 41200
rect 4896 41055 4948 41064
rect 4896 41021 4905 41055
rect 4905 41021 4939 41055
rect 4939 41021 4948 41055
rect 4896 41012 4948 41021
rect 8576 41055 8628 41064
rect 8576 41021 8585 41055
rect 8585 41021 8619 41055
rect 8619 41021 8628 41055
rect 8576 41012 8628 41021
rect 10048 41055 10100 41064
rect 5816 40876 5868 40928
rect 6000 40876 6052 40928
rect 10048 41021 10057 41055
rect 10057 41021 10091 41055
rect 10091 41021 10100 41055
rect 10048 41012 10100 41021
rect 20260 41216 20312 41268
rect 21088 41216 21140 41268
rect 21180 41216 21232 41268
rect 21272 41216 21324 41268
rect 21732 41216 21784 41268
rect 19708 41123 19760 41132
rect 19708 41089 19717 41123
rect 19717 41089 19751 41123
rect 19751 41089 19760 41123
rect 19708 41080 19760 41089
rect 19892 41080 19944 41132
rect 16304 41012 16356 41064
rect 20536 41123 20588 41132
rect 20536 41089 20545 41123
rect 20545 41089 20579 41123
rect 20579 41089 20588 41123
rect 20536 41080 20588 41089
rect 20444 41012 20496 41064
rect 21088 41123 21140 41132
rect 21088 41089 21097 41123
rect 21097 41089 21131 41123
rect 21131 41089 21140 41123
rect 21088 41080 21140 41089
rect 21180 41080 21232 41132
rect 21364 41123 21416 41132
rect 21364 41089 21373 41123
rect 21373 41089 21407 41123
rect 21407 41089 21416 41123
rect 21364 41080 21416 41089
rect 21548 41080 21600 41132
rect 21916 41080 21968 41132
rect 22284 41216 22336 41268
rect 23388 41216 23440 41268
rect 25044 41216 25096 41268
rect 22100 41148 22152 41200
rect 22192 41080 22244 41132
rect 22560 41123 22612 41132
rect 22560 41089 22569 41123
rect 22569 41089 22603 41123
rect 22603 41089 22612 41123
rect 22560 41080 22612 41089
rect 23112 41080 23164 41132
rect 9588 40919 9640 40928
rect 9588 40885 9597 40919
rect 9597 40885 9631 40919
rect 9631 40885 9640 40919
rect 9588 40876 9640 40885
rect 9680 40876 9732 40928
rect 19708 40944 19760 40996
rect 19984 40944 20036 40996
rect 20812 40944 20864 40996
rect 22744 41012 22796 41064
rect 23204 41012 23256 41064
rect 22008 40944 22060 40996
rect 22652 40944 22704 40996
rect 11060 40919 11112 40928
rect 11060 40885 11069 40919
rect 11069 40885 11103 40919
rect 11103 40885 11112 40919
rect 11060 40876 11112 40885
rect 19064 40919 19116 40928
rect 19064 40885 19073 40919
rect 19073 40885 19107 40919
rect 19107 40885 19116 40919
rect 19064 40876 19116 40885
rect 20628 40876 20680 40928
rect 20720 40876 20772 40928
rect 21916 40876 21968 40928
rect 22284 40876 22336 40928
rect 23664 40919 23716 40928
rect 23664 40885 23673 40919
rect 23673 40885 23707 40919
rect 23707 40885 23716 40919
rect 23664 40876 23716 40885
rect 3917 40774 3969 40826
rect 3981 40774 4033 40826
rect 4045 40774 4097 40826
rect 4109 40774 4161 40826
rect 4173 40774 4225 40826
rect 9851 40774 9903 40826
rect 9915 40774 9967 40826
rect 9979 40774 10031 40826
rect 10043 40774 10095 40826
rect 10107 40774 10159 40826
rect 15785 40774 15837 40826
rect 15849 40774 15901 40826
rect 15913 40774 15965 40826
rect 15977 40774 16029 40826
rect 16041 40774 16093 40826
rect 21719 40774 21771 40826
rect 21783 40774 21835 40826
rect 21847 40774 21899 40826
rect 21911 40774 21963 40826
rect 21975 40774 22027 40826
rect 3056 40672 3108 40724
rect 3148 40604 3200 40656
rect 3516 40536 3568 40588
rect 3792 40579 3844 40588
rect 3792 40545 3801 40579
rect 3801 40545 3835 40579
rect 3835 40545 3844 40579
rect 3792 40536 3844 40545
rect 3332 40468 3384 40520
rect 3976 40468 4028 40520
rect 5264 40672 5316 40724
rect 7656 40672 7708 40724
rect 9680 40672 9732 40724
rect 9772 40672 9824 40724
rect 11796 40672 11848 40724
rect 4896 40536 4948 40588
rect 1400 40443 1452 40452
rect 1400 40409 1409 40443
rect 1409 40409 1443 40443
rect 1443 40409 1452 40443
rect 1400 40400 1452 40409
rect 2228 40443 2280 40452
rect 2228 40409 2237 40443
rect 2237 40409 2271 40443
rect 2271 40409 2280 40443
rect 2228 40400 2280 40409
rect 2780 40400 2832 40452
rect 3516 40400 3568 40452
rect 3792 40332 3844 40384
rect 5816 40511 5868 40520
rect 5816 40477 5823 40511
rect 5823 40477 5857 40511
rect 5857 40477 5868 40511
rect 5816 40468 5868 40477
rect 6828 40468 6880 40520
rect 9312 40536 9364 40588
rect 10324 40604 10376 40656
rect 10508 40647 10560 40656
rect 10508 40613 10517 40647
rect 10517 40613 10551 40647
rect 10551 40613 10560 40647
rect 10508 40604 10560 40613
rect 16304 40672 16356 40724
rect 16396 40672 16448 40724
rect 19800 40672 19852 40724
rect 20812 40715 20864 40724
rect 20812 40681 20821 40715
rect 20821 40681 20855 40715
rect 20855 40681 20864 40715
rect 20812 40672 20864 40681
rect 20996 40672 21048 40724
rect 22100 40672 22152 40724
rect 22560 40672 22612 40724
rect 22744 40715 22796 40724
rect 22744 40681 22753 40715
rect 22753 40681 22787 40715
rect 22787 40681 22796 40715
rect 22744 40672 22796 40681
rect 23020 40715 23072 40724
rect 23020 40681 23029 40715
rect 23029 40681 23063 40715
rect 23063 40681 23072 40715
rect 23020 40672 23072 40681
rect 24032 40672 24084 40724
rect 10048 40579 10100 40588
rect 10048 40545 10057 40579
rect 10057 40545 10091 40579
rect 10091 40545 10100 40579
rect 10048 40536 10100 40545
rect 10876 40579 10928 40588
rect 7656 40468 7708 40520
rect 6092 40400 6144 40452
rect 6368 40400 6420 40452
rect 9772 40468 9824 40520
rect 6644 40332 6696 40384
rect 7932 40375 7984 40384
rect 7932 40341 7941 40375
rect 7941 40341 7975 40375
rect 7975 40341 7984 40375
rect 7932 40332 7984 40341
rect 9128 40332 9180 40384
rect 9772 40332 9824 40384
rect 9956 40468 10008 40520
rect 10876 40545 10910 40579
rect 10910 40545 10928 40579
rect 10876 40536 10928 40545
rect 11060 40579 11112 40588
rect 11060 40545 11069 40579
rect 11069 40545 11103 40579
rect 11103 40545 11112 40579
rect 11060 40536 11112 40545
rect 10784 40511 10836 40520
rect 10784 40477 10793 40511
rect 10793 40477 10827 40511
rect 10827 40477 10836 40511
rect 10784 40468 10836 40477
rect 11704 40468 11756 40520
rect 20260 40647 20312 40656
rect 20260 40613 20269 40647
rect 20269 40613 20303 40647
rect 20303 40613 20312 40647
rect 20260 40604 20312 40613
rect 19064 40536 19116 40588
rect 12532 40468 12584 40520
rect 12716 40468 12768 40520
rect 19524 40468 19576 40520
rect 20168 40511 20220 40520
rect 20168 40477 20177 40511
rect 20177 40477 20211 40511
rect 20211 40477 20220 40511
rect 20168 40468 20220 40477
rect 21180 40536 21232 40588
rect 21364 40536 21416 40588
rect 25320 40604 25372 40656
rect 13544 40400 13596 40452
rect 19156 40400 19208 40452
rect 20996 40511 21048 40520
rect 20996 40477 21005 40511
rect 21005 40477 21039 40511
rect 21039 40477 21048 40511
rect 20996 40468 21048 40477
rect 21272 40511 21324 40520
rect 21272 40477 21281 40511
rect 21281 40477 21315 40511
rect 21315 40477 21324 40511
rect 21272 40468 21324 40477
rect 11520 40332 11572 40384
rect 12348 40332 12400 40384
rect 12532 40332 12584 40384
rect 19432 40375 19484 40384
rect 19432 40341 19441 40375
rect 19441 40341 19475 40375
rect 19475 40341 19484 40375
rect 19432 40332 19484 40341
rect 19616 40375 19668 40384
rect 19616 40341 19625 40375
rect 19625 40341 19659 40375
rect 19659 40341 19668 40375
rect 19616 40332 19668 40341
rect 19800 40332 19852 40384
rect 21732 40400 21784 40452
rect 21640 40332 21692 40384
rect 22744 40536 22796 40588
rect 22376 40511 22428 40520
rect 22376 40477 22385 40511
rect 22385 40477 22419 40511
rect 22419 40477 22428 40511
rect 22376 40468 22428 40477
rect 22652 40511 22704 40520
rect 22652 40477 22661 40511
rect 22661 40477 22695 40511
rect 22695 40477 22704 40511
rect 22652 40468 22704 40477
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 23664 40468 23716 40477
rect 22284 40400 22336 40452
rect 25136 40400 25188 40452
rect 22928 40332 22980 40384
rect 6884 40230 6936 40282
rect 6948 40230 7000 40282
rect 7012 40230 7064 40282
rect 7076 40230 7128 40282
rect 7140 40230 7192 40282
rect 12818 40230 12870 40282
rect 12882 40230 12934 40282
rect 12946 40230 12998 40282
rect 13010 40230 13062 40282
rect 13074 40230 13126 40282
rect 18752 40230 18804 40282
rect 18816 40230 18868 40282
rect 18880 40230 18932 40282
rect 18944 40230 18996 40282
rect 19008 40230 19060 40282
rect 24686 40230 24738 40282
rect 24750 40230 24802 40282
rect 24814 40230 24866 40282
rect 24878 40230 24930 40282
rect 24942 40230 24994 40282
rect 3148 40128 3200 40180
rect 3516 40128 3568 40180
rect 7472 40171 7524 40180
rect 7472 40137 7481 40171
rect 7481 40137 7515 40171
rect 7515 40137 7524 40171
rect 7472 40128 7524 40137
rect 8024 40128 8076 40180
rect 9312 40128 9364 40180
rect 1584 39992 1636 40044
rect 3148 39992 3200 40044
rect 3424 39992 3476 40044
rect 1860 39924 1912 39976
rect 3056 39924 3108 39976
rect 7564 40060 7616 40112
rect 8392 40060 8444 40112
rect 7656 39992 7708 40044
rect 8024 39992 8076 40044
rect 8116 39992 8168 40044
rect 9128 40103 9180 40112
rect 9128 40069 9137 40103
rect 9137 40069 9171 40103
rect 9171 40069 9180 40103
rect 9128 40060 9180 40069
rect 9220 40060 9272 40112
rect 9496 40103 9548 40112
rect 9496 40069 9505 40103
rect 9505 40069 9539 40103
rect 9539 40069 9548 40103
rect 9496 40060 9548 40069
rect 9772 40060 9824 40112
rect 10048 40060 10100 40112
rect 10324 40060 10376 40112
rect 10692 40060 10744 40112
rect 10784 40060 10836 40112
rect 9680 39992 9732 40044
rect 12716 40035 12768 40044
rect 12716 40001 12725 40035
rect 12725 40001 12759 40035
rect 12759 40001 12768 40035
rect 12716 39992 12768 40001
rect 19616 40128 19668 40180
rect 19800 40171 19852 40180
rect 19800 40137 19809 40171
rect 19809 40137 19843 40171
rect 19843 40137 19852 40171
rect 19800 40128 19852 40137
rect 20076 40171 20128 40180
rect 20076 40137 20085 40171
rect 20085 40137 20119 40171
rect 20119 40137 20128 40171
rect 20076 40128 20128 40137
rect 4344 39924 4396 39976
rect 4804 39924 4856 39976
rect 4896 39967 4948 39976
rect 4896 39933 4905 39967
rect 4905 39933 4939 39967
rect 4939 39933 4948 39967
rect 4896 39924 4948 39933
rect 7932 39924 7984 39976
rect 9588 39924 9640 39976
rect 11428 39924 11480 39976
rect 11888 39924 11940 39976
rect 12348 39924 12400 39976
rect 13360 39924 13412 39976
rect 19984 40035 20036 40044
rect 19984 40001 19993 40035
rect 19993 40001 20027 40035
rect 20027 40001 20036 40035
rect 19984 39992 20036 40001
rect 20720 40060 20772 40112
rect 21548 40060 21600 40112
rect 20812 40035 20864 40044
rect 20812 40001 20821 40035
rect 20821 40001 20855 40035
rect 20855 40001 20864 40035
rect 20812 39992 20864 40001
rect 21088 40035 21140 40044
rect 21088 40001 21097 40035
rect 21097 40001 21131 40035
rect 21131 40001 21140 40035
rect 21088 39992 21140 40001
rect 21364 40035 21416 40044
rect 21364 40001 21373 40035
rect 21373 40001 21407 40035
rect 21407 40001 21416 40035
rect 21364 39992 21416 40001
rect 21732 39992 21784 40044
rect 22468 39992 22520 40044
rect 2872 39856 2924 39908
rect 3976 39856 4028 39908
rect 12532 39856 12584 39908
rect 19432 39899 19484 39908
rect 19432 39865 19441 39899
rect 19441 39865 19475 39899
rect 19475 39865 19484 39899
rect 19432 39856 19484 39865
rect 20812 39856 20864 39908
rect 23020 39992 23072 40044
rect 23848 40128 23900 40180
rect 2320 39788 2372 39840
rect 3424 39788 3476 39840
rect 4252 39788 4304 39840
rect 5356 39788 5408 39840
rect 5908 39831 5960 39840
rect 5908 39797 5917 39831
rect 5917 39797 5951 39831
rect 5951 39797 5960 39831
rect 5908 39788 5960 39797
rect 8668 39788 8720 39840
rect 10324 39788 10376 39840
rect 13636 39831 13688 39840
rect 13636 39797 13645 39831
rect 13645 39797 13679 39831
rect 13679 39797 13688 39831
rect 13636 39788 13688 39797
rect 22836 39856 22888 39908
rect 23020 39856 23072 39908
rect 23756 39992 23808 40044
rect 24032 39992 24084 40044
rect 21088 39788 21140 39840
rect 21640 39788 21692 39840
rect 22284 39788 22336 39840
rect 22928 39831 22980 39840
rect 22928 39797 22937 39831
rect 22937 39797 22971 39831
rect 22971 39797 22980 39831
rect 22928 39788 22980 39797
rect 23940 39788 23992 39840
rect 24400 39831 24452 39840
rect 24400 39797 24409 39831
rect 24409 39797 24443 39831
rect 24443 39797 24452 39831
rect 24400 39788 24452 39797
rect 3917 39686 3969 39738
rect 3981 39686 4033 39738
rect 4045 39686 4097 39738
rect 4109 39686 4161 39738
rect 4173 39686 4225 39738
rect 9851 39686 9903 39738
rect 9915 39686 9967 39738
rect 9979 39686 10031 39738
rect 10043 39686 10095 39738
rect 10107 39686 10159 39738
rect 15785 39686 15837 39738
rect 15849 39686 15901 39738
rect 15913 39686 15965 39738
rect 15977 39686 16029 39738
rect 16041 39686 16093 39738
rect 21719 39686 21771 39738
rect 21783 39686 21835 39738
rect 21847 39686 21899 39738
rect 21911 39686 21963 39738
rect 21975 39686 22027 39738
rect 3424 39584 3476 39636
rect 5908 39584 5960 39636
rect 3240 39559 3292 39568
rect 3240 39525 3249 39559
rect 3249 39525 3283 39559
rect 3283 39525 3292 39559
rect 3240 39516 3292 39525
rect 2688 39448 2740 39500
rect 3792 39448 3844 39500
rect 5080 39448 5132 39500
rect 5448 39491 5500 39500
rect 5448 39457 5457 39491
rect 5457 39457 5491 39491
rect 5491 39457 5500 39491
rect 5448 39448 5500 39457
rect 6736 39584 6788 39636
rect 8392 39627 8444 39636
rect 8392 39593 8401 39627
rect 8401 39593 8435 39627
rect 8435 39593 8444 39627
rect 8392 39584 8444 39593
rect 9496 39584 9548 39636
rect 13360 39627 13412 39636
rect 13360 39593 13369 39627
rect 13369 39593 13403 39627
rect 13403 39593 13412 39627
rect 13360 39584 13412 39593
rect 13636 39584 13688 39636
rect 20904 39584 20956 39636
rect 20996 39584 21048 39636
rect 22192 39584 22244 39636
rect 22376 39627 22428 39636
rect 22376 39593 22385 39627
rect 22385 39593 22419 39627
rect 22419 39593 22428 39627
rect 22376 39584 22428 39593
rect 22836 39627 22888 39636
rect 22836 39593 22845 39627
rect 22845 39593 22879 39627
rect 22879 39593 22888 39627
rect 22836 39584 22888 39593
rect 8668 39516 8720 39568
rect 21180 39516 21232 39568
rect 21364 39516 21416 39568
rect 6644 39491 6696 39500
rect 6644 39457 6653 39491
rect 6653 39457 6687 39491
rect 6687 39457 6696 39491
rect 6644 39448 6696 39457
rect 6828 39448 6880 39500
rect 7380 39491 7432 39500
rect 7380 39457 7389 39491
rect 7389 39457 7423 39491
rect 7423 39457 7432 39491
rect 7380 39448 7432 39457
rect 11704 39448 11756 39500
rect 20444 39448 20496 39500
rect 20720 39448 20772 39500
rect 4528 39380 4580 39432
rect 1492 39355 1544 39364
rect 1492 39321 1501 39355
rect 1501 39321 1535 39355
rect 1535 39321 1544 39355
rect 1492 39312 1544 39321
rect 1676 39355 1728 39364
rect 1676 39321 1685 39355
rect 1685 39321 1719 39355
rect 1719 39321 1728 39355
rect 1676 39312 1728 39321
rect 2320 39355 2372 39364
rect 2320 39321 2329 39355
rect 2329 39321 2363 39355
rect 2363 39321 2372 39355
rect 2320 39312 2372 39321
rect 2596 39312 2648 39364
rect 4252 39355 4304 39364
rect 4252 39321 4261 39355
rect 4261 39321 4295 39355
rect 4295 39321 4304 39355
rect 4252 39312 4304 39321
rect 6368 39423 6420 39432
rect 6368 39389 6377 39423
rect 6377 39389 6411 39423
rect 6411 39389 6420 39423
rect 6368 39380 6420 39389
rect 7564 39380 7616 39432
rect 8576 39380 8628 39432
rect 10232 39380 10284 39432
rect 16488 39380 16540 39432
rect 20904 39423 20956 39432
rect 20904 39389 20913 39423
rect 20913 39389 20947 39423
rect 20947 39389 20956 39423
rect 20904 39380 20956 39389
rect 3608 39244 3660 39296
rect 4068 39244 4120 39296
rect 4160 39244 4212 39296
rect 4528 39244 4580 39296
rect 8024 39312 8076 39364
rect 10324 39312 10376 39364
rect 11980 39312 12032 39364
rect 20076 39312 20128 39364
rect 20812 39312 20864 39364
rect 4896 39244 4948 39296
rect 5356 39244 5408 39296
rect 20444 39244 20496 39296
rect 21456 39380 21508 39432
rect 22008 39423 22060 39432
rect 22008 39389 22017 39423
rect 22017 39389 22051 39423
rect 22051 39389 22060 39423
rect 22008 39380 22060 39389
rect 22284 39423 22336 39432
rect 22284 39389 22293 39423
rect 22293 39389 22327 39423
rect 22327 39389 22336 39423
rect 22284 39380 22336 39389
rect 22560 39423 22612 39432
rect 22560 39389 22569 39423
rect 22569 39389 22603 39423
rect 22603 39389 22612 39423
rect 22560 39380 22612 39389
rect 21456 39244 21508 39296
rect 23848 39423 23900 39432
rect 23848 39389 23857 39423
rect 23857 39389 23891 39423
rect 23891 39389 23900 39423
rect 23848 39380 23900 39389
rect 23940 39423 23992 39432
rect 23940 39389 23949 39423
rect 23949 39389 23983 39423
rect 23983 39389 23992 39423
rect 23940 39380 23992 39389
rect 23940 39244 23992 39296
rect 25228 39244 25280 39296
rect 6884 39142 6936 39194
rect 6948 39142 7000 39194
rect 7012 39142 7064 39194
rect 7076 39142 7128 39194
rect 7140 39142 7192 39194
rect 12818 39142 12870 39194
rect 12882 39142 12934 39194
rect 12946 39142 12998 39194
rect 13010 39142 13062 39194
rect 13074 39142 13126 39194
rect 18752 39142 18804 39194
rect 18816 39142 18868 39194
rect 18880 39142 18932 39194
rect 18944 39142 18996 39194
rect 19008 39142 19060 39194
rect 24686 39142 24738 39194
rect 24750 39142 24802 39194
rect 24814 39142 24866 39194
rect 24878 39142 24930 39194
rect 24942 39142 24994 39194
rect 1492 39040 1544 39092
rect 4160 39040 4212 39092
rect 4896 39040 4948 39092
rect 5356 39040 5408 39092
rect 6368 39040 6420 39092
rect 8024 39040 8076 39092
rect 11704 39040 11756 39092
rect 20444 39083 20496 39092
rect 20444 39049 20453 39083
rect 20453 39049 20487 39083
rect 20487 39049 20496 39083
rect 20444 39040 20496 39049
rect 20904 39040 20956 39092
rect 21456 39040 21508 39092
rect 1860 38904 1912 38956
rect 2872 38904 2924 38956
rect 3056 38947 3108 38956
rect 3056 38913 3065 38947
rect 3065 38913 3099 38947
rect 3099 38913 3108 38947
rect 3056 38904 3108 38913
rect 3424 38904 3476 38956
rect 2688 38836 2740 38888
rect 3516 38836 3568 38888
rect 3884 38836 3936 38888
rect 5264 38904 5316 38956
rect 7380 38904 7432 38956
rect 5908 38836 5960 38888
rect 6828 38836 6880 38888
rect 8300 38972 8352 39024
rect 8668 38972 8720 39024
rect 16488 38972 16540 39024
rect 21180 38972 21232 39024
rect 8392 38947 8444 38956
rect 8392 38913 8399 38947
rect 8399 38913 8433 38947
rect 8433 38913 8444 38947
rect 8392 38904 8444 38913
rect 19248 38904 19300 38956
rect 11520 38879 11572 38888
rect 11520 38845 11529 38879
rect 11529 38845 11563 38879
rect 11563 38845 11572 38879
rect 11520 38836 11572 38845
rect 20628 38931 20680 38940
rect 20628 38897 20637 38931
rect 20637 38897 20671 38931
rect 20671 38897 20680 38931
rect 20628 38888 20680 38897
rect 20904 38947 20956 38956
rect 20904 38913 20913 38947
rect 20913 38913 20947 38947
rect 20947 38913 20956 38947
rect 20904 38904 20956 38913
rect 20444 38836 20496 38888
rect 21824 38879 21876 38888
rect 21824 38845 21833 38879
rect 21833 38845 21867 38879
rect 21867 38845 21876 38879
rect 21824 38836 21876 38845
rect 23848 39040 23900 39092
rect 23572 38947 23624 38956
rect 23572 38913 23581 38947
rect 23581 38913 23615 38947
rect 23615 38913 23624 38947
rect 23572 38904 23624 38913
rect 23664 38904 23716 38956
rect 24032 38904 24084 38956
rect 16672 38768 16724 38820
rect 20076 38768 20128 38820
rect 23480 38768 23532 38820
rect 5264 38700 5316 38752
rect 8576 38700 8628 38752
rect 9128 38743 9180 38752
rect 9128 38709 9137 38743
rect 9137 38709 9171 38743
rect 9171 38709 9180 38743
rect 9128 38700 9180 38709
rect 12532 38743 12584 38752
rect 12532 38709 12541 38743
rect 12541 38709 12575 38743
rect 12575 38709 12584 38743
rect 12532 38700 12584 38709
rect 17132 38700 17184 38752
rect 20904 38700 20956 38752
rect 22100 38700 22152 38752
rect 24400 38743 24452 38752
rect 24400 38709 24409 38743
rect 24409 38709 24443 38743
rect 24443 38709 24452 38743
rect 24400 38700 24452 38709
rect 3917 38598 3969 38650
rect 3981 38598 4033 38650
rect 4045 38598 4097 38650
rect 4109 38598 4161 38650
rect 4173 38598 4225 38650
rect 9851 38598 9903 38650
rect 9915 38598 9967 38650
rect 9979 38598 10031 38650
rect 10043 38598 10095 38650
rect 10107 38598 10159 38650
rect 15785 38598 15837 38650
rect 15849 38598 15901 38650
rect 15913 38598 15965 38650
rect 15977 38598 16029 38650
rect 16041 38598 16093 38650
rect 21719 38598 21771 38650
rect 21783 38598 21835 38650
rect 21847 38598 21899 38650
rect 21911 38598 21963 38650
rect 21975 38598 22027 38650
rect 1860 38292 1912 38344
rect 5264 38496 5316 38548
rect 756 38224 808 38276
rect 2228 38267 2280 38276
rect 2228 38233 2237 38267
rect 2237 38233 2271 38267
rect 2271 38233 2280 38267
rect 2228 38224 2280 38233
rect 1216 38156 1268 38208
rect 2872 38224 2924 38276
rect 3056 38224 3108 38276
rect 5080 38292 5132 38344
rect 9220 38496 9272 38548
rect 11704 38496 11756 38548
rect 6000 38471 6052 38480
rect 6000 38437 6009 38471
rect 6009 38437 6043 38471
rect 6043 38437 6052 38471
rect 6000 38428 6052 38437
rect 11336 38428 11388 38480
rect 11888 38428 11940 38480
rect 8300 38360 8352 38412
rect 8668 38360 8720 38412
rect 5540 38335 5592 38344
rect 5540 38301 5549 38335
rect 5549 38301 5583 38335
rect 5583 38301 5592 38335
rect 5540 38292 5592 38301
rect 6276 38335 6328 38344
rect 6276 38301 6285 38335
rect 6285 38301 6319 38335
rect 6319 38301 6328 38335
rect 6276 38292 6328 38301
rect 6552 38335 6604 38344
rect 6552 38301 6561 38335
rect 6561 38301 6595 38335
rect 6595 38301 6604 38335
rect 6552 38292 6604 38301
rect 7656 38292 7708 38344
rect 9496 38292 9548 38344
rect 4804 38199 4856 38208
rect 4804 38165 4813 38199
rect 4813 38165 4847 38199
rect 4847 38165 4856 38199
rect 4804 38156 4856 38165
rect 5356 38156 5408 38208
rect 6828 38156 6880 38208
rect 7472 38156 7524 38208
rect 7932 38224 7984 38276
rect 12532 38496 12584 38548
rect 13268 38539 13320 38548
rect 13268 38505 13277 38539
rect 13277 38505 13311 38539
rect 13311 38505 13320 38539
rect 13268 38496 13320 38505
rect 20628 38496 20680 38548
rect 21088 38496 21140 38548
rect 22928 38496 22980 38548
rect 23572 38496 23624 38548
rect 23756 38496 23808 38548
rect 20720 38428 20772 38480
rect 22744 38428 22796 38480
rect 11980 38360 12032 38412
rect 23112 38360 23164 38412
rect 11336 38292 11388 38344
rect 12348 38335 12400 38344
rect 12348 38301 12357 38335
rect 12357 38301 12391 38335
rect 12391 38301 12400 38335
rect 12348 38292 12400 38301
rect 12624 38335 12676 38344
rect 12624 38301 12633 38335
rect 12633 38301 12667 38335
rect 12667 38301 12676 38335
rect 12624 38292 12676 38301
rect 10140 38199 10192 38208
rect 10140 38165 10149 38199
rect 10149 38165 10183 38199
rect 10183 38165 10192 38199
rect 10140 38156 10192 38165
rect 22100 38335 22152 38344
rect 22100 38301 22109 38335
rect 22109 38301 22143 38335
rect 22143 38301 22152 38335
rect 22100 38292 22152 38301
rect 22652 38335 22704 38344
rect 22652 38301 22661 38335
rect 22661 38301 22695 38335
rect 22695 38301 22704 38335
rect 22652 38292 22704 38301
rect 22928 38335 22980 38344
rect 22928 38301 22937 38335
rect 22937 38301 22971 38335
rect 22971 38301 22980 38335
rect 22928 38292 22980 38301
rect 23020 38224 23072 38276
rect 23480 38335 23532 38344
rect 23480 38301 23489 38335
rect 23489 38301 23523 38335
rect 23523 38301 23532 38335
rect 23480 38292 23532 38301
rect 23940 38335 23992 38344
rect 23940 38301 23949 38335
rect 23949 38301 23983 38335
rect 23983 38301 23992 38335
rect 23940 38292 23992 38301
rect 22192 38199 22244 38208
rect 22192 38165 22201 38199
rect 22201 38165 22235 38199
rect 22235 38165 22244 38199
rect 22192 38156 22244 38165
rect 22836 38156 22888 38208
rect 22928 38199 22980 38208
rect 22928 38165 22937 38199
rect 22937 38165 22971 38199
rect 22971 38165 22980 38199
rect 22928 38156 22980 38165
rect 25228 38156 25280 38208
rect 6884 38054 6936 38106
rect 6948 38054 7000 38106
rect 7012 38054 7064 38106
rect 7076 38054 7128 38106
rect 7140 38054 7192 38106
rect 12818 38054 12870 38106
rect 12882 38054 12934 38106
rect 12946 38054 12998 38106
rect 13010 38054 13062 38106
rect 13074 38054 13126 38106
rect 18752 38054 18804 38106
rect 18816 38054 18868 38106
rect 18880 38054 18932 38106
rect 18944 38054 18996 38106
rect 19008 38054 19060 38106
rect 24686 38054 24738 38106
rect 24750 38054 24802 38106
rect 24814 38054 24866 38106
rect 24878 38054 24930 38106
rect 24942 38054 24994 38106
rect 2044 37884 2096 37936
rect 3516 37927 3568 37936
rect 3516 37893 3525 37927
rect 3525 37893 3559 37927
rect 3559 37893 3568 37927
rect 3516 37884 3568 37893
rect 4804 37952 4856 38004
rect 6552 37952 6604 38004
rect 8300 37952 8352 38004
rect 8944 37995 8996 38004
rect 8944 37961 8953 37995
rect 8953 37961 8987 37995
rect 8987 37961 8996 37995
rect 8944 37952 8996 37961
rect 1400 37859 1452 37868
rect 1400 37825 1409 37859
rect 1409 37825 1443 37859
rect 1443 37825 1452 37859
rect 1400 37816 1452 37825
rect 1124 37748 1176 37800
rect 3608 37816 3660 37868
rect 4160 37816 4212 37868
rect 4528 37884 4580 37936
rect 7840 37884 7892 37936
rect 8116 37884 8168 37936
rect 8760 37884 8812 37936
rect 9220 37927 9272 37936
rect 9220 37893 9229 37927
rect 9229 37893 9263 37927
rect 9263 37893 9272 37927
rect 9220 37884 9272 37893
rect 10140 37952 10192 38004
rect 11980 37952 12032 38004
rect 12348 37952 12400 38004
rect 12624 37952 12676 38004
rect 20168 37952 20220 38004
rect 22192 37952 22244 38004
rect 9496 37884 9548 37936
rect 4804 37816 4856 37868
rect 4988 37859 5040 37868
rect 4988 37825 4997 37859
rect 4997 37825 5031 37859
rect 5031 37825 5040 37859
rect 4988 37816 5040 37825
rect 1860 37748 1912 37800
rect 4896 37748 4948 37800
rect 7564 37816 7616 37868
rect 9680 37859 9732 37868
rect 9680 37825 9689 37859
rect 9689 37825 9723 37859
rect 9723 37825 9732 37859
rect 9680 37816 9732 37825
rect 9772 37816 9824 37868
rect 11520 37816 11572 37868
rect 6092 37748 6144 37800
rect 9128 37748 9180 37800
rect 5264 37612 5316 37664
rect 6276 37612 6328 37664
rect 7380 37612 7432 37664
rect 8668 37612 8720 37664
rect 8944 37612 8996 37664
rect 10600 37612 10652 37664
rect 13636 37816 13688 37868
rect 15292 37816 15344 37868
rect 20260 37748 20312 37800
rect 22560 37884 22612 37936
rect 22744 37952 22796 38004
rect 22928 37952 22980 38004
rect 24032 37859 24084 37868
rect 24032 37825 24041 37859
rect 24041 37825 24075 37859
rect 24075 37825 24084 37859
rect 24032 37816 24084 37825
rect 22928 37748 22980 37800
rect 22836 37723 22888 37732
rect 22836 37689 22845 37723
rect 22845 37689 22879 37723
rect 22879 37689 22888 37723
rect 22836 37680 22888 37689
rect 14096 37612 14148 37664
rect 21640 37612 21692 37664
rect 24400 37655 24452 37664
rect 24400 37621 24409 37655
rect 24409 37621 24443 37655
rect 24443 37621 24452 37655
rect 24400 37612 24452 37621
rect 25412 37612 25464 37664
rect 3917 37510 3969 37562
rect 3981 37510 4033 37562
rect 4045 37510 4097 37562
rect 4109 37510 4161 37562
rect 4173 37510 4225 37562
rect 9851 37510 9903 37562
rect 9915 37510 9967 37562
rect 9979 37510 10031 37562
rect 10043 37510 10095 37562
rect 10107 37510 10159 37562
rect 15785 37510 15837 37562
rect 15849 37510 15901 37562
rect 15913 37510 15965 37562
rect 15977 37510 16029 37562
rect 16041 37510 16093 37562
rect 21719 37510 21771 37562
rect 21783 37510 21835 37562
rect 21847 37510 21899 37562
rect 21911 37510 21963 37562
rect 21975 37510 22027 37562
rect 3884 37408 3936 37460
rect 4988 37408 5040 37460
rect 5632 37408 5684 37460
rect 6552 37408 6604 37460
rect 7380 37340 7432 37392
rect 8116 37340 8168 37392
rect 21640 37451 21692 37460
rect 21640 37417 21649 37451
rect 21649 37417 21683 37451
rect 21683 37417 21692 37451
rect 21640 37408 21692 37417
rect 22652 37408 22704 37460
rect 23112 37408 23164 37460
rect 1952 37272 2004 37324
rect 2872 37204 2924 37256
rect 4988 37247 5040 37256
rect 1492 37136 1544 37188
rect 2228 37179 2280 37188
rect 2228 37145 2237 37179
rect 2237 37145 2271 37179
rect 2271 37145 2280 37179
rect 2228 37136 2280 37145
rect 2780 37179 2832 37188
rect 2780 37145 2789 37179
rect 2789 37145 2823 37179
rect 2823 37145 2832 37179
rect 2780 37136 2832 37145
rect 1676 37068 1728 37120
rect 4068 37179 4120 37188
rect 2964 37068 3016 37120
rect 4068 37145 4077 37179
rect 4077 37145 4111 37179
rect 4111 37145 4120 37179
rect 4068 37136 4120 37145
rect 4988 37213 4995 37247
rect 4995 37213 5029 37247
rect 5029 37213 5040 37247
rect 4988 37204 5040 37213
rect 5356 37204 5408 37256
rect 5724 37204 5776 37256
rect 3424 37111 3476 37120
rect 3424 37077 3433 37111
rect 3433 37077 3467 37111
rect 3467 37077 3476 37111
rect 3424 37068 3476 37077
rect 4620 37068 4672 37120
rect 5448 37068 5500 37120
rect 5908 37068 5960 37120
rect 8024 37247 8076 37256
rect 8024 37213 8033 37247
rect 8033 37213 8067 37247
rect 8067 37213 8076 37247
rect 8024 37204 8076 37213
rect 8484 37247 8536 37256
rect 8484 37213 8493 37247
rect 8493 37213 8527 37247
rect 8527 37213 8536 37247
rect 8484 37204 8536 37213
rect 9036 37204 9088 37256
rect 10048 37247 10100 37256
rect 10048 37213 10057 37247
rect 10057 37213 10091 37247
rect 10091 37213 10100 37247
rect 10048 37204 10100 37213
rect 9772 37136 9824 37188
rect 16396 37272 16448 37324
rect 16764 37272 16816 37324
rect 18512 37272 18564 37324
rect 19340 37272 19392 37324
rect 23020 37340 23072 37392
rect 14372 37204 14424 37256
rect 17224 37204 17276 37256
rect 20720 37247 20772 37256
rect 20720 37213 20729 37247
rect 20729 37213 20763 37247
rect 20763 37213 20772 37247
rect 20720 37204 20772 37213
rect 21824 37247 21876 37256
rect 21824 37213 21833 37247
rect 21833 37213 21867 37247
rect 21867 37213 21876 37247
rect 21824 37204 21876 37213
rect 22284 37272 22336 37324
rect 22100 37247 22152 37256
rect 22100 37213 22109 37247
rect 22109 37213 22143 37247
rect 22143 37213 22152 37247
rect 22100 37204 22152 37213
rect 22192 37204 22244 37256
rect 22744 37247 22796 37256
rect 22744 37213 22753 37247
rect 22753 37213 22787 37247
rect 22787 37213 22796 37247
rect 22744 37204 22796 37213
rect 24124 37315 24176 37324
rect 24124 37281 24133 37315
rect 24133 37281 24167 37315
rect 24167 37281 24176 37315
rect 24124 37272 24176 37281
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 23664 37204 23716 37256
rect 23940 37204 23992 37256
rect 11060 37111 11112 37120
rect 11060 37077 11069 37111
rect 11069 37077 11103 37111
rect 11103 37077 11112 37111
rect 11060 37068 11112 37077
rect 11244 37068 11296 37120
rect 18144 37068 18196 37120
rect 20536 37111 20588 37120
rect 20536 37077 20545 37111
rect 20545 37077 20579 37111
rect 20579 37077 20588 37111
rect 20536 37068 20588 37077
rect 22192 37068 22244 37120
rect 23848 37179 23900 37188
rect 23848 37145 23857 37179
rect 23857 37145 23891 37179
rect 23891 37145 23900 37179
rect 23848 37136 23900 37145
rect 6884 36966 6936 37018
rect 6948 36966 7000 37018
rect 7012 36966 7064 37018
rect 7076 36966 7128 37018
rect 7140 36966 7192 37018
rect 12818 36966 12870 37018
rect 12882 36966 12934 37018
rect 12946 36966 12998 37018
rect 13010 36966 13062 37018
rect 13074 36966 13126 37018
rect 18752 36966 18804 37018
rect 18816 36966 18868 37018
rect 18880 36966 18932 37018
rect 18944 36966 18996 37018
rect 19008 36966 19060 37018
rect 24686 36966 24738 37018
rect 24750 36966 24802 37018
rect 24814 36966 24866 37018
rect 24878 36966 24930 37018
rect 24942 36966 24994 37018
rect 2504 36728 2556 36780
rect 3516 36796 3568 36848
rect 3608 36796 3660 36848
rect 8024 36864 8076 36916
rect 8208 36864 8260 36916
rect 8484 36864 8536 36916
rect 7472 36796 7524 36848
rect 9772 36796 9824 36848
rect 4344 36728 4396 36780
rect 4712 36728 4764 36780
rect 1768 36635 1820 36644
rect 1768 36601 1777 36635
rect 1777 36601 1811 36635
rect 1811 36601 1820 36635
rect 1768 36592 1820 36601
rect 4804 36660 4856 36712
rect 6920 36771 6972 36780
rect 6920 36737 6929 36771
rect 6929 36737 6963 36771
rect 6963 36737 6972 36771
rect 6920 36728 6972 36737
rect 7012 36728 7064 36780
rect 7104 36728 7156 36780
rect 7748 36771 7800 36780
rect 7748 36737 7755 36771
rect 7755 36737 7789 36771
rect 7789 36737 7800 36771
rect 7748 36728 7800 36737
rect 9128 36728 9180 36780
rect 9312 36728 9364 36780
rect 17224 36864 17276 36916
rect 14372 36796 14424 36848
rect 19340 36796 19392 36848
rect 20720 36864 20772 36916
rect 21824 36864 21876 36916
rect 16672 36728 16724 36780
rect 7472 36703 7524 36712
rect 2320 36524 2372 36576
rect 4620 36524 4672 36576
rect 4804 36524 4856 36576
rect 7472 36669 7481 36703
rect 7481 36669 7515 36703
rect 7515 36669 7524 36703
rect 7472 36660 7524 36669
rect 8208 36660 8260 36712
rect 10048 36660 10100 36712
rect 10784 36660 10836 36712
rect 8392 36524 8444 36576
rect 8944 36524 8996 36576
rect 10508 36524 10560 36576
rect 17408 36660 17460 36712
rect 17316 36592 17368 36644
rect 12532 36567 12584 36576
rect 12532 36533 12541 36567
rect 12541 36533 12575 36567
rect 12575 36533 12584 36567
rect 12532 36524 12584 36533
rect 17960 36524 18012 36576
rect 18236 36592 18288 36644
rect 19340 36592 19392 36644
rect 19708 36592 19760 36644
rect 20536 36771 20588 36780
rect 20536 36737 20545 36771
rect 20545 36737 20579 36771
rect 20579 36737 20588 36771
rect 20536 36728 20588 36737
rect 23848 36864 23900 36916
rect 24032 36864 24084 36916
rect 23020 36771 23072 36780
rect 23020 36737 23029 36771
rect 23029 36737 23063 36771
rect 23063 36737 23072 36771
rect 23020 36728 23072 36737
rect 24032 36728 24084 36780
rect 22376 36660 22428 36712
rect 25596 36728 25648 36780
rect 20536 36524 20588 36576
rect 24216 36592 24268 36644
rect 22836 36567 22888 36576
rect 22836 36533 22845 36567
rect 22845 36533 22879 36567
rect 22879 36533 22888 36567
rect 22836 36524 22888 36533
rect 24400 36567 24452 36576
rect 24400 36533 24409 36567
rect 24409 36533 24443 36567
rect 24443 36533 24452 36567
rect 24400 36524 24452 36533
rect 3917 36422 3969 36474
rect 3981 36422 4033 36474
rect 4045 36422 4097 36474
rect 4109 36422 4161 36474
rect 4173 36422 4225 36474
rect 9851 36422 9903 36474
rect 9915 36422 9967 36474
rect 9979 36422 10031 36474
rect 10043 36422 10095 36474
rect 10107 36422 10159 36474
rect 15785 36422 15837 36474
rect 15849 36422 15901 36474
rect 15913 36422 15965 36474
rect 15977 36422 16029 36474
rect 16041 36422 16093 36474
rect 21719 36422 21771 36474
rect 21783 36422 21835 36474
rect 21847 36422 21899 36474
rect 21911 36422 21963 36474
rect 21975 36422 22027 36474
rect 1768 36320 1820 36372
rect 2504 36320 2556 36372
rect 3148 36252 3200 36304
rect 3424 36252 3476 36304
rect 3792 36252 3844 36304
rect 4620 36252 4672 36304
rect 4804 36252 4856 36304
rect 1676 36116 1728 36168
rect 2872 36159 2924 36168
rect 2872 36125 2881 36159
rect 2881 36125 2915 36159
rect 2915 36125 2924 36159
rect 2872 36116 2924 36125
rect 2044 35980 2096 36032
rect 2688 35980 2740 36032
rect 3056 35980 3108 36032
rect 4344 36184 4396 36236
rect 4528 36184 4580 36236
rect 4712 36184 4764 36236
rect 3792 36159 3844 36168
rect 3792 36125 3801 36159
rect 3801 36125 3835 36159
rect 3835 36125 3844 36159
rect 3792 36116 3844 36125
rect 4804 36116 4856 36168
rect 5080 36159 5132 36168
rect 5080 36125 5089 36159
rect 5089 36125 5123 36159
rect 5123 36125 5132 36159
rect 5080 36116 5132 36125
rect 5448 36252 5500 36304
rect 6920 36320 6972 36372
rect 7840 36320 7892 36372
rect 8024 36320 8076 36372
rect 22100 36320 22152 36372
rect 22376 36363 22428 36372
rect 22376 36329 22385 36363
rect 22385 36329 22419 36363
rect 22419 36329 22428 36363
rect 22376 36320 22428 36329
rect 22836 36320 22888 36372
rect 23572 36320 23624 36372
rect 5356 36184 5408 36236
rect 6460 36184 6512 36236
rect 6644 36184 6696 36236
rect 4068 36091 4120 36100
rect 4068 36057 4077 36091
rect 4077 36057 4111 36091
rect 4111 36057 4120 36091
rect 4068 36048 4120 36057
rect 3608 35980 3660 36032
rect 4896 35980 4948 36032
rect 5080 35980 5132 36032
rect 6000 36159 6052 36168
rect 6000 36125 6009 36159
rect 6009 36125 6043 36159
rect 6043 36125 6052 36159
rect 6000 36116 6052 36125
rect 7104 36116 7156 36168
rect 11060 36252 11112 36304
rect 7472 36184 7524 36236
rect 8944 36227 8996 36236
rect 8944 36193 8953 36227
rect 8953 36193 8987 36227
rect 8987 36193 8996 36227
rect 8944 36184 8996 36193
rect 9864 36184 9916 36236
rect 10600 36184 10652 36236
rect 12532 36252 12584 36304
rect 7380 36116 7432 36168
rect 8668 36116 8720 36168
rect 9312 36116 9364 36168
rect 9680 36116 9732 36168
rect 5540 35980 5592 36032
rect 7012 35980 7064 36032
rect 7380 35980 7432 36032
rect 7748 35980 7800 36032
rect 9864 35980 9916 36032
rect 9956 36023 10008 36032
rect 9956 35989 9965 36023
rect 9965 35989 9999 36023
rect 9999 35989 10008 36023
rect 9956 35980 10008 35989
rect 10140 36048 10192 36100
rect 11244 36159 11296 36168
rect 11244 36125 11253 36159
rect 11253 36125 11287 36159
rect 11287 36125 11296 36159
rect 11244 36116 11296 36125
rect 11428 36116 11480 36168
rect 17408 36091 17460 36100
rect 17408 36057 17420 36091
rect 17420 36057 17460 36091
rect 17408 36048 17460 36057
rect 19248 36116 19300 36168
rect 20260 36116 20312 36168
rect 14280 35980 14332 36032
rect 19340 35980 19392 36032
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 25136 36048 25188 36100
rect 6884 35878 6936 35930
rect 6948 35878 7000 35930
rect 7012 35878 7064 35930
rect 7076 35878 7128 35930
rect 7140 35878 7192 35930
rect 12818 35878 12870 35930
rect 12882 35878 12934 35930
rect 12946 35878 12998 35930
rect 13010 35878 13062 35930
rect 13074 35878 13126 35930
rect 18752 35878 18804 35930
rect 18816 35878 18868 35930
rect 18880 35878 18932 35930
rect 18944 35878 18996 35930
rect 19008 35878 19060 35930
rect 24686 35878 24738 35930
rect 24750 35878 24802 35930
rect 24814 35878 24866 35930
rect 24878 35878 24930 35930
rect 24942 35878 24994 35930
rect 3332 35819 3384 35828
rect 3332 35785 3341 35819
rect 3341 35785 3375 35819
rect 3375 35785 3384 35819
rect 3332 35776 3384 35785
rect 4528 35776 4580 35828
rect 5264 35776 5316 35828
rect 6644 35776 6696 35828
rect 2688 35683 2740 35692
rect 2688 35649 2697 35683
rect 2697 35649 2731 35683
rect 2731 35649 2740 35683
rect 2688 35640 2740 35649
rect 3424 35683 3476 35692
rect 3424 35649 3433 35683
rect 3433 35649 3467 35683
rect 3467 35649 3476 35683
rect 3424 35640 3476 35649
rect 8208 35751 8260 35760
rect 8208 35717 8217 35751
rect 8217 35717 8251 35751
rect 8251 35717 8260 35751
rect 8208 35708 8260 35717
rect 9956 35776 10008 35828
rect 11704 35819 11756 35828
rect 11704 35785 11713 35819
rect 11713 35785 11747 35819
rect 11747 35785 11756 35819
rect 11704 35776 11756 35785
rect 9220 35708 9272 35760
rect 11244 35708 11296 35760
rect 11428 35708 11480 35760
rect 11980 35751 12032 35760
rect 11980 35717 11989 35751
rect 11989 35717 12023 35751
rect 12023 35717 12032 35751
rect 11980 35708 12032 35717
rect 15200 35776 15252 35828
rect 18236 35776 18288 35828
rect 19340 35776 19392 35828
rect 12348 35708 12400 35760
rect 1216 35572 1268 35624
rect 2136 35547 2188 35556
rect 2136 35513 2145 35547
rect 2145 35513 2179 35547
rect 2179 35513 2188 35547
rect 2136 35504 2188 35513
rect 1952 35436 2004 35488
rect 2504 35615 2556 35624
rect 2504 35581 2538 35615
rect 2538 35581 2556 35615
rect 2504 35572 2556 35581
rect 3056 35572 3108 35624
rect 3608 35615 3660 35624
rect 3608 35581 3617 35615
rect 3617 35581 3651 35615
rect 3651 35581 3660 35615
rect 3608 35572 3660 35581
rect 8760 35640 8812 35692
rect 9588 35640 9640 35692
rect 10416 35640 10468 35692
rect 10968 35640 11020 35692
rect 12624 35708 12676 35760
rect 18420 35708 18472 35760
rect 4620 35572 4672 35624
rect 5264 35615 5316 35624
rect 5264 35581 5273 35615
rect 5273 35581 5307 35615
rect 5307 35581 5316 35615
rect 5264 35572 5316 35581
rect 5356 35615 5408 35624
rect 5356 35581 5390 35615
rect 5390 35581 5408 35615
rect 5356 35572 5408 35581
rect 8392 35572 8444 35624
rect 9312 35572 9364 35624
rect 4896 35504 4948 35556
rect 2504 35436 2556 35488
rect 4528 35436 4580 35488
rect 6368 35504 6420 35556
rect 12808 35572 12860 35624
rect 12900 35572 12952 35624
rect 5448 35436 5500 35488
rect 6000 35436 6052 35488
rect 6460 35436 6512 35488
rect 7840 35436 7892 35488
rect 9772 35436 9824 35488
rect 10600 35436 10652 35488
rect 12992 35479 13044 35488
rect 12992 35445 13001 35479
rect 13001 35445 13035 35479
rect 13035 35445 13044 35479
rect 12992 35436 13044 35445
rect 16764 35640 16816 35692
rect 23020 35776 23072 35828
rect 23572 35776 23624 35828
rect 17592 35615 17644 35624
rect 17592 35581 17601 35615
rect 17601 35581 17635 35615
rect 17635 35581 17644 35615
rect 17592 35572 17644 35581
rect 19064 35615 19116 35624
rect 19064 35581 19073 35615
rect 19073 35581 19107 35615
rect 19107 35581 19116 35615
rect 19064 35572 19116 35581
rect 18880 35504 18932 35556
rect 23204 35640 23256 35692
rect 25136 35708 25188 35760
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 23756 35479 23808 35488
rect 23756 35445 23765 35479
rect 23765 35445 23799 35479
rect 23799 35445 23808 35479
rect 23756 35436 23808 35445
rect 24400 35479 24452 35488
rect 24400 35445 24409 35479
rect 24409 35445 24443 35479
rect 24443 35445 24452 35479
rect 24400 35436 24452 35445
rect 3917 35334 3969 35386
rect 3981 35334 4033 35386
rect 4045 35334 4097 35386
rect 4109 35334 4161 35386
rect 4173 35334 4225 35386
rect 9851 35334 9903 35386
rect 9915 35334 9967 35386
rect 9979 35334 10031 35386
rect 10043 35334 10095 35386
rect 10107 35334 10159 35386
rect 15785 35334 15837 35386
rect 15849 35334 15901 35386
rect 15913 35334 15965 35386
rect 15977 35334 16029 35386
rect 16041 35334 16093 35386
rect 21719 35334 21771 35386
rect 21783 35334 21835 35386
rect 21847 35334 21899 35386
rect 21911 35334 21963 35386
rect 21975 35334 22027 35386
rect 1952 35232 2004 35284
rect 2320 35139 2372 35148
rect 2320 35105 2329 35139
rect 2329 35105 2363 35139
rect 2363 35105 2372 35139
rect 2320 35096 2372 35105
rect 3240 35096 3292 35148
rect 5448 35164 5500 35216
rect 6368 35232 6420 35284
rect 7656 35232 7708 35284
rect 7840 35232 7892 35284
rect 9588 35232 9640 35284
rect 7380 35164 7432 35216
rect 11612 35232 11664 35284
rect 11796 35232 11848 35284
rect 12072 35232 12124 35284
rect 12808 35275 12860 35284
rect 12808 35241 12817 35275
rect 12817 35241 12851 35275
rect 12851 35241 12860 35275
rect 12808 35232 12860 35241
rect 13636 35232 13688 35284
rect 10416 35164 10468 35216
rect 10600 35164 10652 35216
rect 19064 35232 19116 35284
rect 756 35028 808 35080
rect 2044 35028 2096 35080
rect 4252 35071 4304 35080
rect 4252 35037 4261 35071
rect 4261 35037 4295 35071
rect 4295 35037 4304 35071
rect 4252 35028 4304 35037
rect 6644 35096 6696 35148
rect 10140 35096 10192 35148
rect 3516 34892 3568 34944
rect 4344 35003 4396 35012
rect 4344 34969 4353 35003
rect 4353 34969 4387 35003
rect 4387 34969 4396 35003
rect 4344 34960 4396 34969
rect 5448 35071 5500 35080
rect 5448 35037 5457 35071
rect 5457 35037 5491 35071
rect 5491 35037 5500 35071
rect 5448 35028 5500 35037
rect 5632 35028 5684 35080
rect 8576 35028 8628 35080
rect 9680 35028 9732 35080
rect 11244 35096 11296 35148
rect 4712 35003 4764 35012
rect 4712 34969 4721 35003
rect 4721 34969 4755 35003
rect 4755 34969 4764 35003
rect 4712 34960 4764 34969
rect 9956 34960 10008 35012
rect 5080 34935 5132 34944
rect 5080 34901 5089 34935
rect 5089 34901 5123 34935
rect 5123 34901 5132 34935
rect 5080 34892 5132 34901
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 5448 34892 5500 34944
rect 5724 34892 5776 34944
rect 6736 34892 6788 34944
rect 10968 35028 11020 35080
rect 11060 35071 11112 35080
rect 11060 35037 11069 35071
rect 11069 35037 11103 35071
rect 11103 35037 11112 35071
rect 11060 35028 11112 35037
rect 15292 35096 15344 35148
rect 16488 35096 16540 35148
rect 18052 35096 18104 35148
rect 22468 35232 22520 35284
rect 23664 35232 23716 35284
rect 24584 35232 24636 35284
rect 11980 35028 12032 35080
rect 12900 35028 12952 35080
rect 14372 35071 14424 35080
rect 14372 35037 14379 35071
rect 14379 35037 14413 35071
rect 14413 35037 14424 35071
rect 14372 35028 14424 35037
rect 15200 35028 15252 35080
rect 16304 35028 16356 35080
rect 17960 35028 18012 35080
rect 19340 35028 19392 35080
rect 12900 34892 12952 34944
rect 19156 34960 19208 35012
rect 23388 35071 23440 35080
rect 23388 35037 23397 35071
rect 23397 35037 23431 35071
rect 23431 35037 23440 35071
rect 23388 35028 23440 35037
rect 14464 34892 14516 34944
rect 16856 34892 16908 34944
rect 17960 34892 18012 34944
rect 18144 34892 18196 34944
rect 19524 34935 19576 34944
rect 19524 34901 19533 34935
rect 19533 34901 19567 34935
rect 19567 34901 19576 34935
rect 19524 34892 19576 34901
rect 23480 34935 23532 34944
rect 23480 34901 23489 34935
rect 23489 34901 23523 34935
rect 23523 34901 23532 34935
rect 23480 34892 23532 34901
rect 25228 34892 25280 34944
rect 6884 34790 6936 34842
rect 6948 34790 7000 34842
rect 7012 34790 7064 34842
rect 7076 34790 7128 34842
rect 7140 34790 7192 34842
rect 12818 34790 12870 34842
rect 12882 34790 12934 34842
rect 12946 34790 12998 34842
rect 13010 34790 13062 34842
rect 13074 34790 13126 34842
rect 18752 34790 18804 34842
rect 18816 34790 18868 34842
rect 18880 34790 18932 34842
rect 18944 34790 18996 34842
rect 19008 34790 19060 34842
rect 24686 34790 24738 34842
rect 24750 34790 24802 34842
rect 24814 34790 24866 34842
rect 24878 34790 24930 34842
rect 24942 34790 24994 34842
rect 2136 34688 2188 34740
rect 4344 34688 4396 34740
rect 4620 34688 4672 34740
rect 4988 34688 5040 34740
rect 5080 34688 5132 34740
rect 8944 34688 8996 34740
rect 9036 34731 9088 34740
rect 9036 34697 9045 34731
rect 9045 34697 9079 34731
rect 9079 34697 9088 34731
rect 9036 34688 9088 34697
rect 9220 34688 9272 34740
rect 9864 34688 9916 34740
rect 9956 34688 10008 34740
rect 10416 34688 10468 34740
rect 11060 34731 11112 34740
rect 11060 34697 11069 34731
rect 11069 34697 11103 34731
rect 11103 34697 11112 34731
rect 11060 34688 11112 34697
rect 11888 34688 11940 34740
rect 12624 34688 12676 34740
rect 15292 34688 15344 34740
rect 15384 34688 15436 34740
rect 19156 34688 19208 34740
rect 8484 34620 8536 34672
rect 1584 34552 1636 34604
rect 2044 34552 2096 34604
rect 2320 34552 2372 34604
rect 2780 34595 2832 34604
rect 2780 34561 2789 34595
rect 2789 34561 2823 34595
rect 2823 34561 2832 34595
rect 2780 34552 2832 34561
rect 3884 34552 3936 34604
rect 4160 34552 4212 34604
rect 5080 34552 5132 34604
rect 5448 34552 5500 34604
rect 5724 34552 5776 34604
rect 9680 34620 9732 34672
rect 10048 34620 10100 34672
rect 10692 34620 10744 34672
rect 16488 34620 16540 34672
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 4528 34484 4580 34536
rect 6184 34484 6236 34536
rect 2228 34416 2280 34468
rect 3332 34416 3384 34468
rect 4620 34416 4672 34468
rect 4988 34416 5040 34468
rect 1216 34348 1268 34400
rect 2504 34348 2556 34400
rect 3608 34348 3660 34400
rect 3884 34348 3936 34400
rect 5448 34348 5500 34400
rect 7380 34391 7432 34400
rect 7380 34357 7389 34391
rect 7389 34357 7423 34391
rect 7423 34357 7432 34391
rect 7380 34348 7432 34357
rect 7472 34348 7524 34400
rect 7656 34348 7708 34400
rect 8116 34348 8168 34400
rect 9036 34348 9088 34400
rect 9220 34484 9272 34536
rect 9588 34595 9640 34604
rect 9588 34561 9597 34595
rect 9597 34561 9631 34595
rect 9631 34561 9640 34595
rect 9588 34552 9640 34561
rect 10416 34552 10468 34604
rect 13452 34552 13504 34604
rect 13728 34552 13780 34604
rect 16856 34620 16908 34672
rect 9772 34484 9824 34536
rect 10048 34527 10100 34536
rect 10048 34493 10057 34527
rect 10057 34493 10091 34527
rect 10091 34493 10100 34527
rect 10048 34484 10100 34493
rect 14096 34484 14148 34536
rect 17040 34595 17092 34604
rect 17040 34561 17049 34595
rect 17049 34561 17083 34595
rect 17083 34561 17092 34595
rect 17040 34552 17092 34561
rect 17408 34620 17460 34672
rect 19524 34620 19576 34672
rect 20444 34620 20496 34672
rect 17500 34595 17552 34604
rect 17500 34561 17509 34595
rect 17509 34561 17543 34595
rect 17543 34561 17552 34595
rect 17500 34552 17552 34561
rect 9496 34348 9548 34400
rect 9864 34348 9916 34400
rect 10876 34348 10928 34400
rect 19156 34552 19208 34604
rect 19340 34595 19392 34604
rect 19340 34561 19374 34595
rect 19374 34561 19392 34595
rect 19340 34552 19392 34561
rect 22192 34552 22244 34604
rect 23664 34731 23716 34740
rect 23664 34697 23673 34731
rect 23673 34697 23707 34731
rect 23707 34697 23716 34731
rect 23664 34688 23716 34697
rect 23756 34688 23808 34740
rect 23940 34620 23992 34672
rect 23756 34552 23808 34604
rect 21088 34484 21140 34536
rect 24400 34527 24452 34536
rect 24400 34493 24409 34527
rect 24409 34493 24443 34527
rect 24443 34493 24452 34527
rect 24400 34484 24452 34493
rect 19984 34348 20036 34400
rect 20444 34391 20496 34400
rect 20444 34357 20453 34391
rect 20453 34357 20487 34391
rect 20487 34357 20496 34391
rect 20444 34348 20496 34357
rect 21548 34348 21600 34400
rect 23112 34348 23164 34400
rect 3917 34246 3969 34298
rect 3981 34246 4033 34298
rect 4045 34246 4097 34298
rect 4109 34246 4161 34298
rect 4173 34246 4225 34298
rect 9851 34246 9903 34298
rect 9915 34246 9967 34298
rect 9979 34246 10031 34298
rect 10043 34246 10095 34298
rect 10107 34246 10159 34298
rect 15785 34246 15837 34298
rect 15849 34246 15901 34298
rect 15913 34246 15965 34298
rect 15977 34246 16029 34298
rect 16041 34246 16093 34298
rect 21719 34246 21771 34298
rect 21783 34246 21835 34298
rect 21847 34246 21899 34298
rect 21911 34246 21963 34298
rect 21975 34246 22027 34298
rect 2412 34144 2464 34196
rect 3056 34144 3108 34196
rect 2596 34076 2648 34128
rect 3976 34076 4028 34128
rect 848 33940 900 33992
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 2964 34008 3016 34060
rect 5724 34144 5776 34196
rect 4528 34051 4580 34060
rect 4528 34017 4537 34051
rect 4537 34017 4571 34051
rect 4571 34017 4580 34051
rect 4528 34008 4580 34017
rect 2780 33983 2832 33992
rect 2780 33949 2789 33983
rect 2789 33949 2823 33983
rect 2823 33949 2832 33983
rect 2780 33940 2832 33949
rect 1216 33872 1268 33924
rect 3332 33872 3384 33924
rect 7380 34076 7432 34128
rect 6368 34008 6420 34060
rect 6736 33940 6788 33992
rect 8760 34008 8812 34060
rect 6276 33872 6328 33924
rect 2136 33804 2188 33856
rect 5540 33847 5592 33856
rect 5540 33813 5549 33847
rect 5549 33813 5583 33847
rect 5583 33813 5592 33847
rect 5540 33804 5592 33813
rect 8024 33983 8076 33992
rect 8024 33949 8033 33983
rect 8033 33949 8067 33983
rect 8067 33949 8076 33983
rect 8024 33940 8076 33949
rect 8944 33983 8996 33992
rect 8944 33949 8953 33983
rect 8953 33949 8987 33983
rect 8987 33949 8996 33983
rect 8944 33940 8996 33949
rect 9680 34144 9732 34196
rect 14372 34144 14424 34196
rect 10968 34076 11020 34128
rect 13544 34119 13596 34128
rect 13544 34085 13553 34119
rect 13553 34085 13587 34119
rect 13587 34085 13596 34119
rect 13544 34076 13596 34085
rect 17500 34144 17552 34196
rect 17592 34144 17644 34196
rect 9680 34008 9732 34060
rect 14004 34008 14056 34060
rect 15200 34008 15252 34060
rect 10232 33940 10284 33992
rect 11888 33940 11940 33992
rect 13636 33940 13688 33992
rect 14832 33940 14884 33992
rect 15108 33940 15160 33992
rect 16764 33940 16816 33992
rect 17500 33983 17552 33992
rect 17500 33949 17509 33983
rect 17509 33949 17543 33983
rect 17543 33949 17552 33983
rect 17500 33940 17552 33949
rect 7840 33804 7892 33856
rect 8484 33804 8536 33856
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 8944 33804 8996 33856
rect 12440 33804 12492 33856
rect 13176 33804 13228 33856
rect 14372 33804 14424 33856
rect 14924 33804 14976 33856
rect 15384 33872 15436 33924
rect 17408 33872 17460 33924
rect 16948 33847 17000 33856
rect 16948 33813 16957 33847
rect 16957 33813 16991 33847
rect 16991 33813 17000 33847
rect 16948 33804 17000 33813
rect 19892 34144 19944 34196
rect 21088 34187 21140 34196
rect 21088 34153 21097 34187
rect 21097 34153 21131 34187
rect 21131 34153 21140 34187
rect 21088 34144 21140 34153
rect 23388 34144 23440 34196
rect 20260 33940 20312 33992
rect 21548 33983 21600 33992
rect 21548 33949 21557 33983
rect 21557 33949 21591 33983
rect 21591 33949 21600 33983
rect 21548 33940 21600 33949
rect 22560 33983 22612 33992
rect 22560 33949 22569 33983
rect 22569 33949 22603 33983
rect 22603 33949 22612 33983
rect 22560 33940 22612 33949
rect 22836 33983 22888 33992
rect 22836 33949 22845 33983
rect 22845 33949 22879 33983
rect 22879 33949 22888 33983
rect 22836 33940 22888 33949
rect 17776 33804 17828 33856
rect 18236 33847 18288 33856
rect 18236 33813 18245 33847
rect 18245 33813 18279 33847
rect 18279 33813 18288 33847
rect 18236 33804 18288 33813
rect 21640 33804 21692 33856
rect 22652 33847 22704 33856
rect 22652 33813 22661 33847
rect 22661 33813 22695 33847
rect 22695 33813 22704 33847
rect 22652 33804 22704 33813
rect 23480 33940 23532 33992
rect 23480 33804 23532 33856
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 25228 33804 25280 33856
rect 6884 33702 6936 33754
rect 6948 33702 7000 33754
rect 7012 33702 7064 33754
rect 7076 33702 7128 33754
rect 7140 33702 7192 33754
rect 12818 33702 12870 33754
rect 12882 33702 12934 33754
rect 12946 33702 12998 33754
rect 13010 33702 13062 33754
rect 13074 33702 13126 33754
rect 18752 33702 18804 33754
rect 18816 33702 18868 33754
rect 18880 33702 18932 33754
rect 18944 33702 18996 33754
rect 19008 33702 19060 33754
rect 24686 33702 24738 33754
rect 24750 33702 24802 33754
rect 24814 33702 24866 33754
rect 24878 33702 24930 33754
rect 24942 33702 24994 33754
rect 1952 33600 2004 33652
rect 1124 33532 1176 33584
rect 3240 33600 3292 33652
rect 3792 33600 3844 33652
rect 8208 33600 8260 33652
rect 8668 33600 8720 33652
rect 3148 33532 3200 33584
rect 3976 33532 4028 33584
rect 4620 33532 4672 33584
rect 4896 33532 4948 33584
rect 2228 33464 2280 33516
rect 3424 33507 3476 33516
rect 3424 33473 3433 33507
rect 3433 33473 3467 33507
rect 3467 33473 3476 33507
rect 3424 33464 3476 33473
rect 1400 33396 1452 33448
rect 4344 33396 4396 33448
rect 6552 33532 6604 33584
rect 6736 33532 6788 33584
rect 5908 33464 5960 33516
rect 4528 33328 4580 33380
rect 6644 33396 6696 33448
rect 7012 33396 7064 33448
rect 7196 33396 7248 33448
rect 8116 33507 8168 33516
rect 8116 33473 8125 33507
rect 8125 33473 8159 33507
rect 8159 33473 8168 33507
rect 8116 33464 8168 33473
rect 9496 33600 9548 33652
rect 9680 33600 9732 33652
rect 9220 33532 9272 33584
rect 10692 33600 10744 33652
rect 15384 33600 15436 33652
rect 17040 33600 17092 33652
rect 11060 33532 11112 33584
rect 18880 33600 18932 33652
rect 19064 33600 19116 33652
rect 20996 33600 21048 33652
rect 22652 33600 22704 33652
rect 22836 33600 22888 33652
rect 23664 33600 23716 33652
rect 7380 33328 7432 33380
rect 9864 33464 9916 33516
rect 10692 33464 10744 33516
rect 11980 33507 12032 33516
rect 11980 33473 11989 33507
rect 11989 33473 12023 33507
rect 12023 33473 12032 33507
rect 11980 33464 12032 33473
rect 14004 33464 14056 33516
rect 16580 33464 16632 33516
rect 17132 33507 17184 33516
rect 17132 33473 17141 33507
rect 17141 33473 17175 33507
rect 17175 33473 17184 33507
rect 17132 33464 17184 33473
rect 17684 33532 17736 33584
rect 19156 33532 19208 33584
rect 5908 33303 5960 33312
rect 5908 33269 5917 33303
rect 5917 33269 5951 33303
rect 5951 33269 5960 33303
rect 5908 33260 5960 33269
rect 6552 33260 6604 33312
rect 9772 33260 9824 33312
rect 11704 33328 11756 33380
rect 12532 33396 12584 33448
rect 12808 33439 12860 33448
rect 12808 33405 12842 33439
rect 12842 33405 12860 33439
rect 12808 33396 12860 33405
rect 13636 33396 13688 33448
rect 15200 33439 15252 33448
rect 15200 33405 15209 33439
rect 15209 33405 15243 33439
rect 15243 33405 15252 33439
rect 15200 33396 15252 33405
rect 17776 33464 17828 33516
rect 18236 33464 18288 33516
rect 18604 33464 18656 33516
rect 10508 33303 10560 33312
rect 10508 33269 10517 33303
rect 10517 33269 10551 33303
rect 10551 33269 10560 33303
rect 10508 33260 10560 33269
rect 10784 33260 10836 33312
rect 13820 33328 13872 33380
rect 12900 33260 12952 33312
rect 14188 33260 14240 33312
rect 16212 33303 16264 33312
rect 16212 33269 16221 33303
rect 16221 33269 16255 33303
rect 16255 33269 16264 33303
rect 16212 33260 16264 33269
rect 18880 33303 18932 33312
rect 18880 33269 18889 33303
rect 18889 33269 18923 33303
rect 18923 33269 18932 33303
rect 18880 33260 18932 33269
rect 20996 33464 21048 33516
rect 23112 33464 23164 33516
rect 22192 33260 22244 33312
rect 23388 33303 23440 33312
rect 23388 33269 23397 33303
rect 23397 33269 23431 33303
rect 23431 33269 23440 33303
rect 23388 33260 23440 33269
rect 23480 33303 23532 33312
rect 23480 33269 23489 33303
rect 23489 33269 23523 33303
rect 23523 33269 23532 33303
rect 23480 33260 23532 33269
rect 24400 33303 24452 33312
rect 24400 33269 24409 33303
rect 24409 33269 24443 33303
rect 24443 33269 24452 33303
rect 24400 33260 24452 33269
rect 3917 33158 3969 33210
rect 3981 33158 4033 33210
rect 4045 33158 4097 33210
rect 4109 33158 4161 33210
rect 4173 33158 4225 33210
rect 9851 33158 9903 33210
rect 9915 33158 9967 33210
rect 9979 33158 10031 33210
rect 10043 33158 10095 33210
rect 10107 33158 10159 33210
rect 15785 33158 15837 33210
rect 15849 33158 15901 33210
rect 15913 33158 15965 33210
rect 15977 33158 16029 33210
rect 16041 33158 16093 33210
rect 21719 33158 21771 33210
rect 21783 33158 21835 33210
rect 21847 33158 21899 33210
rect 21911 33158 21963 33210
rect 21975 33158 22027 33210
rect 1400 33056 1452 33108
rect 2596 33056 2648 33108
rect 3240 33056 3292 33108
rect 3424 33056 3476 33108
rect 3792 33056 3844 33108
rect 8116 33056 8168 33108
rect 9680 33056 9732 33108
rect 2320 32963 2372 32972
rect 2320 32929 2329 32963
rect 2329 32929 2363 32963
rect 2363 32929 2372 32963
rect 2320 32920 2372 32929
rect 3332 32920 3384 32972
rect 4896 32988 4948 33040
rect 10508 32988 10560 33040
rect 11612 32988 11664 33040
rect 12900 33099 12952 33108
rect 12900 33065 12909 33099
rect 12909 33065 12943 33099
rect 12943 33065 12952 33099
rect 12900 33056 12952 33065
rect 16120 33056 16172 33108
rect 16580 33056 16632 33108
rect 14004 32988 14056 33040
rect 14832 32988 14884 33040
rect 18604 33099 18656 33108
rect 18604 33065 18613 33099
rect 18613 33065 18647 33099
rect 18647 33065 18656 33099
rect 18604 33056 18656 33065
rect 20628 33056 20680 33108
rect 23388 33056 23440 33108
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 1676 32827 1728 32836
rect 1676 32793 1685 32827
rect 1685 32793 1719 32827
rect 1719 32793 1728 32827
rect 1676 32784 1728 32793
rect 3148 32852 3200 32904
rect 5540 32920 5592 32972
rect 6184 32920 6236 32972
rect 9036 32920 9088 32972
rect 10692 32920 10744 32972
rect 11336 32920 11388 32972
rect 3424 32784 3476 32836
rect 1216 32716 1268 32768
rect 5908 32852 5960 32904
rect 6920 32852 6972 32904
rect 4344 32784 4396 32836
rect 4712 32716 4764 32768
rect 5356 32716 5408 32768
rect 7012 32784 7064 32836
rect 8024 32852 8076 32904
rect 8760 32852 8812 32904
rect 9220 32852 9272 32904
rect 5908 32716 5960 32768
rect 6092 32759 6144 32768
rect 6092 32725 6101 32759
rect 6101 32725 6135 32759
rect 6135 32725 6144 32759
rect 6092 32716 6144 32725
rect 6276 32759 6328 32768
rect 6276 32725 6285 32759
rect 6285 32725 6319 32759
rect 6319 32725 6328 32759
rect 6276 32716 6328 32725
rect 7748 32716 7800 32768
rect 10876 32895 10928 32904
rect 10876 32861 10885 32895
rect 10885 32861 10919 32895
rect 10919 32861 10928 32895
rect 10876 32852 10928 32861
rect 11152 32895 11204 32904
rect 11152 32861 11161 32895
rect 11161 32861 11195 32895
rect 11195 32861 11204 32895
rect 11152 32852 11204 32861
rect 11888 32963 11940 32972
rect 11888 32929 11897 32963
rect 11897 32929 11931 32963
rect 11931 32929 11940 32963
rect 11888 32920 11940 32929
rect 13912 32920 13964 32972
rect 17592 32963 17644 32972
rect 17592 32929 17601 32963
rect 17601 32929 17635 32963
rect 17635 32929 17644 32963
rect 17592 32920 17644 32929
rect 21272 32920 21324 32972
rect 22652 32920 22704 32972
rect 12164 32895 12216 32904
rect 12164 32861 12173 32895
rect 12173 32861 12216 32895
rect 12164 32852 12216 32861
rect 12532 32852 12584 32904
rect 14188 32784 14240 32836
rect 10416 32716 10468 32768
rect 12808 32716 12860 32768
rect 15016 32895 15068 32904
rect 15016 32861 15025 32895
rect 15025 32861 15059 32895
rect 15059 32861 15068 32895
rect 15016 32852 15068 32861
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 16028 32852 16080 32904
rect 16120 32852 16172 32904
rect 17408 32852 17460 32904
rect 17776 32852 17828 32904
rect 22100 32895 22152 32904
rect 22100 32861 22101 32895
rect 22101 32861 22135 32895
rect 22135 32861 22152 32895
rect 22100 32852 22152 32861
rect 22192 32897 22244 32904
rect 22192 32863 22201 32897
rect 22201 32863 22235 32897
rect 22235 32863 22244 32897
rect 22192 32852 22244 32863
rect 25688 32920 25740 32972
rect 23756 32852 23808 32904
rect 15200 32716 15252 32768
rect 15384 32716 15436 32768
rect 23296 32784 23348 32836
rect 23940 32895 23992 32904
rect 23940 32861 23949 32895
rect 23949 32861 23983 32895
rect 23983 32861 23992 32895
rect 23940 32852 23992 32861
rect 25044 32784 25096 32836
rect 25228 32716 25280 32768
rect 6884 32614 6936 32666
rect 6948 32614 7000 32666
rect 7012 32614 7064 32666
rect 7076 32614 7128 32666
rect 7140 32614 7192 32666
rect 12818 32614 12870 32666
rect 12882 32614 12934 32666
rect 12946 32614 12998 32666
rect 13010 32614 13062 32666
rect 13074 32614 13126 32666
rect 18752 32614 18804 32666
rect 18816 32614 18868 32666
rect 18880 32614 18932 32666
rect 18944 32614 18996 32666
rect 19008 32614 19060 32666
rect 24686 32614 24738 32666
rect 24750 32614 24802 32666
rect 24814 32614 24866 32666
rect 24878 32614 24930 32666
rect 24942 32614 24994 32666
rect 1124 32512 1176 32564
rect 4620 32512 4672 32564
rect 4988 32512 5040 32564
rect 6092 32512 6144 32564
rect 6276 32512 6328 32564
rect 7564 32512 7616 32564
rect 7748 32512 7800 32564
rect 5724 32444 5776 32496
rect 10140 32444 10192 32496
rect 11152 32512 11204 32564
rect 13912 32512 13964 32564
rect 15200 32555 15252 32564
rect 15200 32521 15209 32555
rect 15209 32521 15243 32555
rect 15243 32521 15252 32555
rect 15200 32512 15252 32521
rect 15384 32555 15436 32564
rect 15384 32521 15393 32555
rect 15393 32521 15427 32555
rect 15427 32521 15436 32555
rect 15384 32512 15436 32521
rect 16764 32512 16816 32564
rect 2412 32419 2464 32428
rect 2412 32385 2446 32419
rect 2446 32385 2464 32419
rect 2412 32376 2464 32385
rect 1492 32308 1544 32360
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 2136 32308 2188 32360
rect 2320 32351 2372 32360
rect 2320 32317 2329 32351
rect 2329 32317 2363 32351
rect 2363 32317 2372 32351
rect 2320 32308 2372 32317
rect 2596 32351 2648 32360
rect 2596 32317 2605 32351
rect 2605 32317 2639 32351
rect 2639 32317 2648 32351
rect 2596 32308 2648 32317
rect 2964 32308 3016 32360
rect 1216 32172 1268 32224
rect 6092 32376 6144 32428
rect 3424 32308 3476 32360
rect 3792 32308 3844 32360
rect 4252 32308 4304 32360
rect 4620 32351 4672 32360
rect 4620 32317 4629 32351
rect 4629 32317 4663 32351
rect 4663 32317 4672 32351
rect 4620 32308 4672 32317
rect 8760 32376 8812 32428
rect 9772 32376 9824 32428
rect 10600 32444 10652 32496
rect 13728 32444 13780 32496
rect 5632 32240 5684 32292
rect 5356 32172 5408 32224
rect 6736 32172 6788 32224
rect 9312 32308 9364 32360
rect 8392 32172 8444 32224
rect 9036 32215 9088 32224
rect 9036 32181 9045 32215
rect 9045 32181 9079 32215
rect 9079 32181 9088 32215
rect 9036 32172 9088 32181
rect 10876 32376 10928 32428
rect 11980 32376 12032 32428
rect 14188 32444 14240 32496
rect 14464 32487 14516 32496
rect 14464 32453 14473 32487
rect 14473 32453 14507 32487
rect 14507 32453 14516 32487
rect 14464 32444 14516 32453
rect 16580 32444 16632 32496
rect 19524 32444 19576 32496
rect 19248 32376 19300 32428
rect 23940 32512 23992 32564
rect 11336 32308 11388 32360
rect 11520 32308 11572 32360
rect 15108 32308 15160 32360
rect 15200 32308 15252 32360
rect 15476 32308 15528 32360
rect 11152 32172 11204 32224
rect 15568 32172 15620 32224
rect 16304 32172 16356 32224
rect 19156 32172 19208 32224
rect 20536 32215 20588 32224
rect 20536 32181 20545 32215
rect 20545 32181 20579 32215
rect 20579 32181 20588 32215
rect 20536 32172 20588 32181
rect 24124 32419 24176 32428
rect 24124 32385 24133 32419
rect 24133 32385 24167 32419
rect 24167 32385 24176 32419
rect 24124 32376 24176 32385
rect 24032 32172 24084 32224
rect 24400 32215 24452 32224
rect 24400 32181 24409 32215
rect 24409 32181 24443 32215
rect 24443 32181 24452 32215
rect 24400 32172 24452 32181
rect 3917 32070 3969 32122
rect 3981 32070 4033 32122
rect 4045 32070 4097 32122
rect 4109 32070 4161 32122
rect 4173 32070 4225 32122
rect 9851 32070 9903 32122
rect 9915 32070 9967 32122
rect 9979 32070 10031 32122
rect 10043 32070 10095 32122
rect 10107 32070 10159 32122
rect 15785 32070 15837 32122
rect 15849 32070 15901 32122
rect 15913 32070 15965 32122
rect 15977 32070 16029 32122
rect 16041 32070 16093 32122
rect 21719 32070 21771 32122
rect 21783 32070 21835 32122
rect 21847 32070 21899 32122
rect 21911 32070 21963 32122
rect 21975 32070 22027 32122
rect 2596 31968 2648 32020
rect 5172 31968 5224 32020
rect 9588 31968 9640 32020
rect 848 31832 900 31884
rect 2412 31832 2464 31884
rect 2964 31832 3016 31884
rect 6736 31900 6788 31952
rect 2688 31764 2740 31816
rect 2780 31807 2832 31816
rect 2780 31773 2789 31807
rect 2789 31773 2823 31807
rect 2823 31773 2832 31807
rect 2780 31764 2832 31773
rect 7656 31832 7708 31884
rect 8116 31832 8168 31884
rect 8392 31832 8444 31884
rect 9128 31832 9180 31884
rect 11888 31968 11940 32020
rect 14464 31968 14516 32020
rect 15108 32011 15160 32020
rect 15108 31977 15117 32011
rect 15117 31977 15151 32011
rect 15151 31977 15160 32011
rect 15108 31968 15160 31977
rect 15292 31968 15344 32020
rect 15568 31968 15620 32020
rect 16212 31943 16264 31952
rect 16212 31909 16221 31943
rect 16221 31909 16255 31943
rect 16255 31909 16264 31943
rect 16212 31900 16264 31909
rect 2228 31696 2280 31748
rect 2412 31696 2464 31748
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 4896 31807 4948 31816
rect 4896 31773 4905 31807
rect 4905 31773 4939 31807
rect 4939 31773 4948 31807
rect 4896 31764 4948 31773
rect 5540 31764 5592 31816
rect 6092 31807 6144 31816
rect 6092 31773 6099 31807
rect 6099 31773 6133 31807
rect 6133 31773 6144 31807
rect 6092 31764 6144 31773
rect 6184 31764 6236 31816
rect 6460 31764 6512 31816
rect 8484 31764 8536 31816
rect 10876 31764 10928 31816
rect 1308 31628 1360 31680
rect 2964 31628 3016 31680
rect 6276 31696 6328 31748
rect 7472 31696 7524 31748
rect 12348 31764 12400 31816
rect 12532 31764 12584 31816
rect 13820 31832 13872 31884
rect 15476 31832 15528 31884
rect 16764 31968 16816 32020
rect 17132 31968 17184 32020
rect 18420 31968 18472 32020
rect 16580 31875 16632 31884
rect 16580 31841 16614 31875
rect 16614 31841 16632 31875
rect 16580 31832 16632 31841
rect 16948 31832 17000 31884
rect 18052 31832 18104 31884
rect 18420 31832 18472 31884
rect 20536 31900 20588 31952
rect 20720 31900 20772 31952
rect 5816 31628 5868 31680
rect 6368 31628 6420 31680
rect 6736 31628 6788 31680
rect 9036 31628 9088 31680
rect 9220 31628 9272 31680
rect 11244 31628 11296 31680
rect 12072 31671 12124 31680
rect 12072 31637 12081 31671
rect 12081 31637 12115 31671
rect 12115 31637 12124 31671
rect 12072 31628 12124 31637
rect 13544 31628 13596 31680
rect 14280 31764 14332 31816
rect 15292 31764 15344 31816
rect 15568 31807 15620 31816
rect 15568 31773 15577 31807
rect 15577 31773 15611 31807
rect 15611 31773 15620 31807
rect 15568 31764 15620 31773
rect 19524 31696 19576 31748
rect 16120 31628 16172 31680
rect 16580 31628 16632 31680
rect 24124 31968 24176 32020
rect 21732 31832 21784 31884
rect 23756 31900 23808 31952
rect 23480 31764 23532 31816
rect 25136 31764 25188 31816
rect 25504 31764 25556 31816
rect 20536 31628 20588 31680
rect 20628 31628 20680 31680
rect 21180 31628 21232 31680
rect 24308 31628 24360 31680
rect 6884 31526 6936 31578
rect 6948 31526 7000 31578
rect 7012 31526 7064 31578
rect 7076 31526 7128 31578
rect 7140 31526 7192 31578
rect 12818 31526 12870 31578
rect 12882 31526 12934 31578
rect 12946 31526 12998 31578
rect 13010 31526 13062 31578
rect 13074 31526 13126 31578
rect 18752 31526 18804 31578
rect 18816 31526 18868 31578
rect 18880 31526 18932 31578
rect 18944 31526 18996 31578
rect 19008 31526 19060 31578
rect 24686 31526 24738 31578
rect 24750 31526 24802 31578
rect 24814 31526 24866 31578
rect 24878 31526 24930 31578
rect 24942 31526 24994 31578
rect 1768 31424 1820 31476
rect 1952 31424 2004 31476
rect 3700 31424 3752 31476
rect 4344 31356 4396 31408
rect 4436 31399 4488 31408
rect 4436 31365 4445 31399
rect 4445 31365 4479 31399
rect 4479 31365 4488 31399
rect 4436 31356 4488 31365
rect 4528 31399 4580 31408
rect 4528 31365 4537 31399
rect 4537 31365 4571 31399
rect 4571 31365 4580 31399
rect 4528 31356 4580 31365
rect 5448 31356 5500 31408
rect 5540 31288 5592 31340
rect 6368 31356 6420 31408
rect 6460 31356 6512 31408
rect 7196 31424 7248 31476
rect 7564 31424 7616 31476
rect 7840 31424 7892 31476
rect 7288 31331 7340 31340
rect 7288 31297 7297 31331
rect 7297 31297 7331 31331
rect 7331 31297 7340 31331
rect 7288 31288 7340 31297
rect 7472 31356 7524 31408
rect 8944 31399 8996 31408
rect 8944 31365 8953 31399
rect 8953 31365 8987 31399
rect 8987 31365 8996 31399
rect 8944 31356 8996 31365
rect 9036 31399 9088 31408
rect 9036 31365 9045 31399
rect 9045 31365 9079 31399
rect 9079 31365 9088 31399
rect 9036 31356 9088 31365
rect 9404 31331 9456 31340
rect 9404 31297 9413 31331
rect 9413 31297 9447 31331
rect 9447 31297 9456 31331
rect 9404 31288 9456 31297
rect 9772 31399 9824 31408
rect 9772 31365 9781 31399
rect 9781 31365 9815 31399
rect 9815 31365 9824 31399
rect 9772 31356 9824 31365
rect 12164 31356 12216 31408
rect 13636 31424 13688 31476
rect 22192 31424 22244 31476
rect 14648 31356 14700 31408
rect 15108 31356 15160 31408
rect 10600 31288 10652 31340
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 3332 31220 3384 31272
rect 6736 31220 6788 31272
rect 9220 31220 9272 31272
rect 1308 31084 1360 31136
rect 5448 31195 5500 31204
rect 5448 31161 5457 31195
rect 5457 31161 5491 31195
rect 5491 31161 5500 31195
rect 5448 31152 5500 31161
rect 6184 31152 6236 31204
rect 7840 31195 7892 31204
rect 7840 31161 7849 31195
rect 7849 31161 7883 31195
rect 7883 31161 7892 31195
rect 7840 31152 7892 31161
rect 10876 31152 10928 31204
rect 2228 31084 2280 31136
rect 6552 31084 6604 31136
rect 11704 31127 11756 31136
rect 11704 31093 11713 31127
rect 11713 31093 11747 31127
rect 11747 31093 11756 31127
rect 11704 31084 11756 31093
rect 13912 31331 13964 31340
rect 12348 31220 12400 31272
rect 12440 31195 12492 31204
rect 12440 31161 12449 31195
rect 12449 31161 12483 31195
rect 12483 31161 12492 31195
rect 12440 31152 12492 31161
rect 13912 31297 13921 31331
rect 13921 31297 13955 31331
rect 13955 31297 13964 31331
rect 13912 31288 13964 31297
rect 16304 31288 16356 31340
rect 17316 31356 17368 31408
rect 14648 31220 14700 31272
rect 16856 31288 16908 31340
rect 23296 31356 23348 31408
rect 17960 31288 18012 31340
rect 19800 31331 19852 31340
rect 19800 31297 19807 31331
rect 19807 31297 19841 31331
rect 19841 31297 19852 31331
rect 19800 31288 19852 31297
rect 20168 31288 20220 31340
rect 20720 31288 20772 31340
rect 21456 31331 21508 31340
rect 21456 31297 21465 31331
rect 21465 31297 21499 31331
rect 21499 31297 21508 31331
rect 21456 31288 21508 31297
rect 22192 31288 22244 31340
rect 12164 31084 12216 31136
rect 14924 31152 14976 31204
rect 14004 31127 14056 31136
rect 14004 31093 14013 31127
rect 14013 31093 14047 31127
rect 14047 31093 14056 31127
rect 14004 31084 14056 31093
rect 14464 31084 14516 31136
rect 16120 31127 16172 31136
rect 16120 31093 16129 31127
rect 16129 31093 16163 31127
rect 16163 31093 16172 31127
rect 16120 31084 16172 31093
rect 17408 31084 17460 31136
rect 18604 31127 18656 31136
rect 18604 31093 18613 31127
rect 18613 31093 18647 31127
rect 18647 31093 18656 31127
rect 18604 31084 18656 31093
rect 20628 31152 20680 31204
rect 23848 31288 23900 31340
rect 21364 31127 21416 31136
rect 21364 31093 21373 31127
rect 21373 31093 21407 31127
rect 21407 31093 21416 31127
rect 21364 31084 21416 31093
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 24400 31127 24452 31136
rect 24400 31093 24409 31127
rect 24409 31093 24443 31127
rect 24443 31093 24452 31127
rect 24400 31084 24452 31093
rect 3917 30982 3969 31034
rect 3981 30982 4033 31034
rect 4045 30982 4097 31034
rect 4109 30982 4161 31034
rect 4173 30982 4225 31034
rect 9851 30982 9903 31034
rect 9915 30982 9967 31034
rect 9979 30982 10031 31034
rect 10043 30982 10095 31034
rect 10107 30982 10159 31034
rect 15785 30982 15837 31034
rect 15849 30982 15901 31034
rect 15913 30982 15965 31034
rect 15977 30982 16029 31034
rect 16041 30982 16093 31034
rect 21719 30982 21771 31034
rect 21783 30982 21835 31034
rect 21847 30982 21899 31034
rect 21911 30982 21963 31034
rect 21975 30982 22027 31034
rect 1584 30880 1636 30932
rect 2320 30880 2372 30932
rect 3332 30923 3384 30932
rect 3332 30889 3341 30923
rect 3341 30889 3375 30923
rect 3375 30889 3384 30923
rect 3332 30880 3384 30889
rect 4528 30880 4580 30932
rect 6000 30880 6052 30932
rect 7196 30880 7248 30932
rect 9036 30880 9088 30932
rect 10140 30880 10192 30932
rect 12348 30880 12400 30932
rect 12532 30923 12584 30932
rect 12532 30889 12541 30923
rect 12541 30889 12575 30923
rect 12575 30889 12584 30923
rect 12532 30880 12584 30889
rect 8392 30812 8444 30864
rect 11060 30812 11112 30864
rect 6276 30744 6328 30796
rect 8300 30744 8352 30796
rect 8944 30787 8996 30796
rect 8944 30753 8953 30787
rect 8953 30753 8987 30787
rect 8987 30753 8996 30787
rect 8944 30744 8996 30753
rect 10416 30744 10468 30796
rect 10784 30744 10836 30796
rect 11152 30787 11204 30796
rect 11152 30753 11161 30787
rect 11161 30753 11195 30787
rect 11195 30753 11204 30787
rect 11152 30744 11204 30753
rect 11428 30787 11480 30796
rect 11428 30753 11437 30787
rect 11437 30753 11471 30787
rect 11471 30753 11480 30787
rect 11428 30744 11480 30753
rect 11520 30787 11572 30796
rect 11520 30753 11554 30787
rect 11554 30753 11572 30787
rect 11520 30744 11572 30753
rect 11888 30744 11940 30796
rect 12072 30744 12124 30796
rect 14648 30880 14700 30932
rect 16120 30880 16172 30932
rect 17408 30880 17460 30932
rect 12532 30744 12584 30796
rect 13912 30744 13964 30796
rect 14004 30744 14056 30796
rect 2136 30676 2188 30728
rect 2596 30719 2648 30728
rect 1492 30651 1544 30660
rect 1492 30617 1501 30651
rect 1501 30617 1535 30651
rect 1535 30617 1544 30651
rect 1492 30608 1544 30617
rect 1676 30651 1728 30660
rect 1676 30617 1685 30651
rect 1685 30617 1719 30651
rect 1719 30617 1728 30651
rect 1676 30608 1728 30617
rect 2596 30685 2603 30719
rect 2603 30685 2637 30719
rect 2637 30685 2648 30719
rect 2596 30676 2648 30685
rect 3792 30719 3844 30728
rect 3792 30685 3801 30719
rect 3801 30685 3835 30719
rect 3835 30685 3844 30719
rect 3792 30676 3844 30685
rect 4160 30676 4212 30728
rect 4436 30676 4488 30728
rect 5356 30676 5408 30728
rect 9128 30676 9180 30728
rect 10600 30676 10652 30728
rect 15108 30787 15160 30796
rect 15108 30753 15117 30787
rect 15117 30753 15151 30787
rect 15151 30753 15160 30787
rect 15108 30744 15160 30753
rect 15568 30744 15620 30796
rect 4344 30608 4396 30660
rect 6828 30608 6880 30660
rect 10324 30608 10376 30660
rect 10508 30608 10560 30660
rect 940 30540 992 30592
rect 1216 30540 1268 30592
rect 4252 30540 4304 30592
rect 12164 30540 12216 30592
rect 12348 30540 12400 30592
rect 13544 30608 13596 30660
rect 15292 30676 15344 30728
rect 16764 30787 16816 30796
rect 16764 30753 16798 30787
rect 16798 30753 16816 30787
rect 16764 30744 16816 30753
rect 16120 30676 16172 30728
rect 16672 30719 16724 30728
rect 16672 30685 16681 30719
rect 16681 30685 16715 30719
rect 16715 30685 16724 30719
rect 16672 30676 16724 30685
rect 17960 30880 18012 30932
rect 18604 30880 18656 30932
rect 17684 30787 17736 30796
rect 17684 30753 17693 30787
rect 17693 30753 17727 30787
rect 17727 30753 17736 30787
rect 17684 30744 17736 30753
rect 20628 30880 20680 30932
rect 21456 30880 21508 30932
rect 20812 30719 20864 30728
rect 20812 30685 20821 30719
rect 20821 30685 20855 30719
rect 20855 30685 20864 30719
rect 20812 30676 20864 30685
rect 22284 30719 22336 30728
rect 22284 30685 22293 30719
rect 22293 30685 22327 30719
rect 22327 30685 22336 30719
rect 22284 30676 22336 30685
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 24584 30676 24636 30728
rect 25872 30676 25924 30728
rect 13452 30540 13504 30592
rect 14464 30540 14516 30592
rect 16304 30540 16356 30592
rect 18604 30540 18656 30592
rect 19248 30540 19300 30592
rect 22560 30540 22612 30592
rect 25136 30608 25188 30660
rect 23296 30540 23348 30592
rect 23572 30540 23624 30592
rect 24584 30540 24636 30592
rect 6884 30438 6936 30490
rect 6948 30438 7000 30490
rect 7012 30438 7064 30490
rect 7076 30438 7128 30490
rect 7140 30438 7192 30490
rect 12818 30438 12870 30490
rect 12882 30438 12934 30490
rect 12946 30438 12998 30490
rect 13010 30438 13062 30490
rect 13074 30438 13126 30490
rect 18752 30438 18804 30490
rect 18816 30438 18868 30490
rect 18880 30438 18932 30490
rect 18944 30438 18996 30490
rect 19008 30438 19060 30490
rect 24686 30438 24738 30490
rect 24750 30438 24802 30490
rect 24814 30438 24866 30490
rect 24878 30438 24930 30490
rect 24942 30438 24994 30490
rect 1308 30268 1360 30320
rect 3976 30336 4028 30388
rect 4436 30336 4488 30388
rect 4712 30336 4764 30388
rect 6460 30268 6512 30320
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 3424 30243 3476 30252
rect 3424 30209 3433 30243
rect 3433 30209 3467 30243
rect 3467 30209 3476 30243
rect 3424 30200 3476 30209
rect 3700 30243 3752 30252
rect 3700 30209 3709 30243
rect 3709 30209 3743 30243
rect 3743 30209 3752 30243
rect 3700 30200 3752 30209
rect 3884 30200 3936 30252
rect 4528 30200 4580 30252
rect 9404 30268 9456 30320
rect 11152 30336 11204 30388
rect 11520 30336 11572 30388
rect 11704 30336 11756 30388
rect 23572 30336 23624 30388
rect 23848 30336 23900 30388
rect 23940 30336 23992 30388
rect 7196 30200 7248 30252
rect 8116 30200 8168 30252
rect 10140 30200 10192 30252
rect 18236 30273 18288 30320
rect 12532 30200 12584 30252
rect 13820 30200 13872 30252
rect 14096 30200 14148 30252
rect 1584 30132 1636 30184
rect 1676 30175 1728 30184
rect 1676 30141 1685 30175
rect 1685 30141 1719 30175
rect 1719 30141 1728 30175
rect 1676 30132 1728 30141
rect 2228 30132 2280 30184
rect 3792 30132 3844 30184
rect 4160 30175 4212 30184
rect 4160 30141 4169 30175
rect 4169 30141 4203 30175
rect 4203 30141 4212 30175
rect 4160 30132 4212 30141
rect 6460 30132 6512 30184
rect 7656 30132 7708 30184
rect 7932 30132 7984 30184
rect 10692 30132 10744 30184
rect 10968 30132 11020 30184
rect 12164 30132 12216 30184
rect 17592 30200 17644 30252
rect 17868 30200 17920 30252
rect 18236 30268 18261 30273
rect 18261 30268 18288 30273
rect 18420 30268 18472 30320
rect 19340 30268 19392 30320
rect 18604 30200 18656 30252
rect 20536 30243 20588 30252
rect 20536 30209 20559 30243
rect 20559 30209 20588 30243
rect 20536 30200 20588 30209
rect 22192 30200 22244 30252
rect 22744 30200 22796 30252
rect 3056 29996 3108 30048
rect 4896 29996 4948 30048
rect 5172 30039 5224 30048
rect 5172 30005 5181 30039
rect 5181 30005 5215 30039
rect 5215 30005 5224 30039
rect 5172 29996 5224 30005
rect 6276 29996 6328 30048
rect 8760 30064 8812 30116
rect 7840 30039 7892 30048
rect 7840 30005 7849 30039
rect 7849 30005 7883 30039
rect 7883 30005 7892 30039
rect 7840 29996 7892 30005
rect 7932 29996 7984 30048
rect 11244 30064 11296 30116
rect 12624 30064 12676 30116
rect 19432 30132 19484 30184
rect 19248 30064 19300 30116
rect 14740 29996 14792 30048
rect 14924 30039 14976 30048
rect 14924 30005 14933 30039
rect 14933 30005 14967 30039
rect 14967 30005 14976 30039
rect 14924 29996 14976 30005
rect 17592 29996 17644 30048
rect 19984 29996 20036 30048
rect 22284 29996 22336 30048
rect 22836 30039 22888 30048
rect 22836 30005 22845 30039
rect 22845 30005 22879 30039
rect 22879 30005 22888 30039
rect 22836 29996 22888 30005
rect 23204 30039 23256 30048
rect 23204 30005 23213 30039
rect 23213 30005 23247 30039
rect 23247 30005 23256 30039
rect 23204 29996 23256 30005
rect 24400 30039 24452 30048
rect 24400 30005 24409 30039
rect 24409 30005 24443 30039
rect 24443 30005 24452 30039
rect 24400 29996 24452 30005
rect 3917 29894 3969 29946
rect 3981 29894 4033 29946
rect 4045 29894 4097 29946
rect 4109 29894 4161 29946
rect 4173 29894 4225 29946
rect 9851 29894 9903 29946
rect 9915 29894 9967 29946
rect 9979 29894 10031 29946
rect 10043 29894 10095 29946
rect 10107 29894 10159 29946
rect 15785 29894 15837 29946
rect 15849 29894 15901 29946
rect 15913 29894 15965 29946
rect 15977 29894 16029 29946
rect 16041 29894 16093 29946
rect 21719 29894 21771 29946
rect 21783 29894 21835 29946
rect 21847 29894 21899 29946
rect 21911 29894 21963 29946
rect 21975 29894 22027 29946
rect 1584 29792 1636 29844
rect 2688 29835 2740 29844
rect 2688 29801 2697 29835
rect 2697 29801 2731 29835
rect 2731 29801 2740 29835
rect 2688 29792 2740 29801
rect 2780 29792 2832 29844
rect 3240 29835 3292 29844
rect 3240 29801 3249 29835
rect 3249 29801 3283 29835
rect 3283 29801 3292 29835
rect 3240 29792 3292 29801
rect 3608 29835 3660 29844
rect 3608 29801 3617 29835
rect 3617 29801 3651 29835
rect 3651 29801 3660 29835
rect 3608 29792 3660 29801
rect 4712 29792 4764 29844
rect 2964 29724 3016 29776
rect 3700 29724 3752 29776
rect 3792 29724 3844 29776
rect 2412 29656 2464 29708
rect 1584 29588 1636 29640
rect 2044 29588 2096 29640
rect 2596 29588 2648 29640
rect 1308 29520 1360 29572
rect 7840 29792 7892 29844
rect 8116 29792 8168 29844
rect 8852 29792 8904 29844
rect 9036 29792 9088 29844
rect 10876 29792 10928 29844
rect 11152 29767 11204 29776
rect 11152 29733 11161 29767
rect 11161 29733 11195 29767
rect 11195 29733 11204 29767
rect 11152 29724 11204 29733
rect 5172 29656 5224 29708
rect 3148 29563 3200 29572
rect 3148 29529 3157 29563
rect 3157 29529 3191 29563
rect 3191 29529 3200 29563
rect 3148 29520 3200 29529
rect 7656 29656 7708 29708
rect 7840 29699 7892 29708
rect 7840 29665 7849 29699
rect 7849 29665 7883 29699
rect 7883 29665 7892 29699
rect 7840 29656 7892 29665
rect 8300 29656 8352 29708
rect 9404 29656 9456 29708
rect 10692 29699 10744 29708
rect 10692 29665 10701 29699
rect 10701 29665 10735 29699
rect 10735 29665 10744 29699
rect 10692 29656 10744 29665
rect 11060 29656 11112 29708
rect 11612 29656 11664 29708
rect 11888 29656 11940 29708
rect 12348 29835 12400 29844
rect 12348 29801 12357 29835
rect 12357 29801 12391 29835
rect 12391 29801 12400 29835
rect 12348 29792 12400 29801
rect 17500 29792 17552 29844
rect 17592 29792 17644 29844
rect 20720 29792 20772 29844
rect 13636 29724 13688 29776
rect 16212 29767 16264 29776
rect 16212 29733 16221 29767
rect 16221 29733 16255 29767
rect 16255 29733 16264 29767
rect 16212 29724 16264 29733
rect 1676 29452 1728 29504
rect 2228 29452 2280 29504
rect 2412 29452 2464 29504
rect 2688 29452 2740 29504
rect 3240 29452 3292 29504
rect 4988 29495 5040 29504
rect 4988 29461 4997 29495
rect 4997 29461 5031 29495
rect 5031 29461 5040 29495
rect 4988 29452 5040 29461
rect 5632 29520 5684 29572
rect 5724 29563 5776 29572
rect 5724 29529 5733 29563
rect 5733 29529 5767 29563
rect 5767 29529 5776 29563
rect 5724 29520 5776 29529
rect 5816 29520 5868 29572
rect 7104 29631 7156 29640
rect 7104 29597 7113 29631
rect 7113 29597 7147 29631
rect 7147 29597 7156 29631
rect 7104 29588 7156 29597
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 10508 29631 10560 29640
rect 10508 29597 10517 29631
rect 10517 29597 10551 29631
rect 10551 29597 10560 29631
rect 10508 29588 10560 29597
rect 7932 29452 7984 29504
rect 8392 29452 8444 29504
rect 9772 29520 9824 29572
rect 8760 29452 8812 29504
rect 12164 29452 12216 29504
rect 13820 29656 13872 29708
rect 12348 29588 12400 29640
rect 12716 29631 12768 29640
rect 12716 29597 12723 29631
rect 12723 29597 12757 29631
rect 12757 29597 12768 29631
rect 12716 29588 12768 29597
rect 15752 29699 15804 29708
rect 15752 29665 15761 29699
rect 15761 29665 15795 29699
rect 15795 29665 15804 29699
rect 15752 29656 15804 29665
rect 16948 29656 17000 29708
rect 12624 29520 12676 29572
rect 13544 29520 13596 29572
rect 14188 29520 14240 29572
rect 14740 29520 14792 29572
rect 15108 29452 15160 29504
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 16580 29631 16632 29640
rect 16580 29597 16614 29631
rect 16614 29597 16632 29631
rect 16580 29588 16632 29597
rect 19248 29520 19300 29572
rect 20536 29520 20588 29572
rect 22836 29792 22888 29844
rect 23204 29792 23256 29844
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 16672 29452 16724 29504
rect 17040 29452 17092 29504
rect 17868 29452 17920 29504
rect 19984 29452 20036 29504
rect 24216 29520 24268 29572
rect 25136 29452 25188 29504
rect 204 29384 256 29436
rect 572 29384 624 29436
rect 6884 29350 6936 29402
rect 6948 29350 7000 29402
rect 7012 29350 7064 29402
rect 7076 29350 7128 29402
rect 7140 29350 7192 29402
rect 12818 29350 12870 29402
rect 12882 29350 12934 29402
rect 12946 29350 12998 29402
rect 13010 29350 13062 29402
rect 13074 29350 13126 29402
rect 18752 29350 18804 29402
rect 18816 29350 18868 29402
rect 18880 29350 18932 29402
rect 18944 29350 18996 29402
rect 19008 29350 19060 29402
rect 24686 29350 24738 29402
rect 24750 29350 24802 29402
rect 24814 29350 24866 29402
rect 24878 29350 24930 29402
rect 24942 29350 24994 29402
rect 664 29248 716 29300
rect 4528 29248 4580 29300
rect 940 29180 992 29232
rect 1952 29180 2004 29232
rect 1492 29155 1544 29164
rect 1492 29121 1501 29155
rect 1501 29121 1535 29155
rect 1535 29121 1544 29155
rect 1492 29112 1544 29121
rect 2872 29112 2924 29164
rect 3608 29155 3660 29164
rect 3608 29121 3617 29155
rect 3617 29121 3651 29155
rect 3651 29121 3660 29155
rect 3608 29112 3660 29121
rect 4988 29180 5040 29232
rect 5632 29248 5684 29300
rect 8116 29248 8168 29300
rect 8576 29248 8628 29300
rect 8852 29248 8904 29300
rect 10692 29248 10744 29300
rect 11244 29248 11296 29300
rect 13728 29248 13780 29300
rect 5172 29155 5224 29164
rect 5172 29121 5179 29155
rect 5179 29121 5213 29155
rect 5213 29121 5224 29155
rect 13360 29180 13412 29232
rect 5172 29112 5224 29121
rect 2136 29044 2188 29096
rect 4896 29087 4948 29096
rect 4896 29053 4905 29087
rect 4905 29053 4939 29087
rect 4939 29053 4948 29087
rect 4896 29044 4948 29053
rect 6460 29112 6512 29164
rect 7196 29112 7248 29164
rect 7656 29155 7708 29164
rect 7656 29121 7663 29155
rect 7663 29121 7697 29155
rect 7697 29121 7708 29155
rect 7656 29112 7708 29121
rect 8760 29112 8812 29164
rect 9404 29112 9456 29164
rect 1952 28976 2004 29028
rect 3240 29019 3292 29028
rect 3240 28985 3249 29019
rect 3249 28985 3283 29019
rect 3283 28985 3292 29019
rect 3240 28976 3292 28985
rect 7104 28976 7156 29028
rect 8576 29044 8628 29096
rect 11336 29112 11388 29164
rect 12072 29112 12124 29164
rect 15200 29180 15252 29232
rect 14740 29112 14792 29164
rect 15108 29112 15160 29164
rect 16580 29180 16632 29232
rect 17592 29180 17644 29232
rect 19156 29185 19208 29232
rect 15568 29112 15620 29164
rect 16948 29155 17000 29164
rect 16948 29121 16955 29155
rect 16955 29121 16989 29155
rect 16989 29121 17000 29155
rect 16948 29112 17000 29121
rect 17868 29112 17920 29164
rect 19156 29180 19181 29185
rect 19181 29180 19208 29185
rect 19524 29180 19576 29232
rect 11152 28976 11204 29028
rect 12532 29087 12584 29096
rect 12532 29053 12541 29087
rect 12541 29053 12575 29087
rect 12575 29053 12584 29087
rect 12532 29044 12584 29053
rect 13452 29044 13504 29096
rect 13636 29044 13688 29096
rect 14924 29044 14976 29096
rect 16672 29087 16724 29096
rect 16672 29053 16681 29087
rect 16681 29053 16715 29087
rect 16715 29053 16724 29087
rect 16672 29044 16724 29053
rect 8116 28908 8168 28960
rect 11060 28908 11112 28960
rect 11428 28908 11480 28960
rect 15476 28976 15528 29028
rect 13728 28908 13780 28960
rect 14096 28908 14148 28960
rect 17132 28908 17184 28960
rect 17868 28908 17920 28960
rect 19800 28976 19852 29028
rect 19616 28908 19668 28960
rect 20260 28908 20312 28960
rect 20352 28951 20404 28960
rect 20352 28917 20361 28951
rect 20361 28917 20395 28951
rect 20395 28917 20404 28951
rect 20352 28908 20404 28917
rect 22744 28908 22796 28960
rect 24400 28951 24452 28960
rect 24400 28917 24409 28951
rect 24409 28917 24443 28951
rect 24443 28917 24452 28951
rect 24400 28908 24452 28917
rect 3917 28806 3969 28858
rect 3981 28806 4033 28858
rect 4045 28806 4097 28858
rect 4109 28806 4161 28858
rect 4173 28806 4225 28858
rect 9851 28806 9903 28858
rect 9915 28806 9967 28858
rect 9979 28806 10031 28858
rect 10043 28806 10095 28858
rect 10107 28806 10159 28858
rect 15785 28806 15837 28858
rect 15849 28806 15901 28858
rect 15913 28806 15965 28858
rect 15977 28806 16029 28858
rect 16041 28806 16093 28858
rect 21719 28806 21771 28858
rect 21783 28806 21835 28858
rect 21847 28806 21899 28858
rect 21911 28806 21963 28858
rect 21975 28806 22027 28858
rect 1584 28704 1636 28756
rect 1860 28704 1912 28756
rect 11152 28747 11204 28756
rect 11152 28713 11161 28747
rect 11161 28713 11195 28747
rect 11195 28713 11204 28747
rect 11152 28704 11204 28713
rect 11428 28747 11480 28756
rect 11428 28713 11437 28747
rect 11437 28713 11471 28747
rect 11471 28713 11480 28747
rect 11428 28704 11480 28713
rect 11612 28704 11664 28756
rect 2136 28568 2188 28620
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 2044 28543 2096 28552
rect 2044 28509 2053 28543
rect 2053 28509 2087 28543
rect 2087 28509 2096 28543
rect 2044 28500 2096 28509
rect 2596 28543 2648 28552
rect 2596 28509 2603 28543
rect 2603 28509 2637 28543
rect 2637 28509 2648 28543
rect 2596 28500 2648 28509
rect 3792 28500 3844 28552
rect 4160 28543 4212 28552
rect 4160 28509 4167 28543
rect 4167 28509 4201 28543
rect 4201 28509 4212 28543
rect 4160 28500 4212 28509
rect 756 28432 808 28484
rect 1676 28432 1728 28484
rect 8116 28568 8168 28620
rect 7196 28500 7248 28552
rect 7748 28500 7800 28552
rect 9220 28543 9272 28552
rect 9220 28509 9227 28543
rect 9227 28509 9261 28543
rect 9261 28509 9272 28543
rect 9220 28500 9272 28509
rect 9588 28500 9640 28552
rect 5264 28432 5316 28484
rect 10416 28432 10468 28484
rect 19524 28704 19576 28756
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 11336 28500 11388 28509
rect 11704 28543 11756 28552
rect 11704 28509 11713 28543
rect 11713 28509 11747 28543
rect 11747 28509 11756 28543
rect 11704 28500 11756 28509
rect 11888 28500 11940 28552
rect 13820 28500 13872 28552
rect 14096 28543 14148 28552
rect 14096 28509 14105 28543
rect 14105 28509 14139 28543
rect 14139 28509 14148 28543
rect 14096 28500 14148 28509
rect 14372 28543 14424 28552
rect 14372 28509 14379 28543
rect 14379 28509 14413 28543
rect 14413 28509 14424 28543
rect 16672 28611 16724 28620
rect 16672 28577 16681 28611
rect 16681 28577 16715 28611
rect 16715 28577 16724 28611
rect 16672 28568 16724 28577
rect 16948 28611 17000 28620
rect 16948 28577 16957 28611
rect 16957 28577 16991 28611
rect 16991 28577 17000 28611
rect 16948 28568 17000 28577
rect 17224 28611 17276 28620
rect 17224 28577 17233 28611
rect 17233 28577 17267 28611
rect 17267 28577 17276 28611
rect 17224 28568 17276 28577
rect 19432 28636 19484 28688
rect 14372 28500 14424 28509
rect 15292 28500 15344 28552
rect 16120 28500 16172 28552
rect 17040 28543 17092 28552
rect 17040 28509 17074 28543
rect 17074 28509 17092 28543
rect 17040 28500 17092 28509
rect 17960 28500 18012 28552
rect 18696 28500 18748 28552
rect 20352 28704 20404 28756
rect 19616 28543 19668 28552
rect 19616 28509 19625 28543
rect 19625 28509 19659 28543
rect 19659 28509 19668 28543
rect 19616 28500 19668 28509
rect 19984 28543 20036 28552
rect 19984 28509 19993 28543
rect 19993 28509 20027 28543
rect 20027 28509 20036 28543
rect 19984 28500 20036 28509
rect 20352 28500 20404 28552
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 1952 28407 2004 28416
rect 1952 28373 1961 28407
rect 1961 28373 1995 28407
rect 1995 28373 2004 28407
rect 1952 28364 2004 28373
rect 3332 28407 3384 28416
rect 3332 28373 3341 28407
rect 3341 28373 3375 28407
rect 3375 28373 3384 28407
rect 3332 28364 3384 28373
rect 4988 28364 5040 28416
rect 5172 28364 5224 28416
rect 5448 28364 5500 28416
rect 6552 28364 6604 28416
rect 7288 28364 7340 28416
rect 9036 28364 9088 28416
rect 9220 28364 9272 28416
rect 9680 28364 9732 28416
rect 10048 28364 10100 28416
rect 11888 28364 11940 28416
rect 13176 28364 13228 28416
rect 13912 28364 13964 28416
rect 14004 28364 14056 28416
rect 14280 28364 14332 28416
rect 20536 28364 20588 28416
rect 20996 28407 21048 28416
rect 20996 28373 21005 28407
rect 21005 28373 21039 28407
rect 21039 28373 21048 28407
rect 20996 28364 21048 28373
rect 25136 28364 25188 28416
rect 6884 28262 6936 28314
rect 6948 28262 7000 28314
rect 7012 28262 7064 28314
rect 7076 28262 7128 28314
rect 7140 28262 7192 28314
rect 12818 28262 12870 28314
rect 12882 28262 12934 28314
rect 12946 28262 12998 28314
rect 13010 28262 13062 28314
rect 13074 28262 13126 28314
rect 18752 28262 18804 28314
rect 18816 28262 18868 28314
rect 18880 28262 18932 28314
rect 18944 28262 18996 28314
rect 19008 28262 19060 28314
rect 24686 28262 24738 28314
rect 24750 28262 24802 28314
rect 24814 28262 24866 28314
rect 24878 28262 24930 28314
rect 24942 28262 24994 28314
rect 1676 28160 1728 28212
rect 3976 28160 4028 28212
rect 2780 28135 2832 28144
rect 2780 28101 2789 28135
rect 2789 28101 2823 28135
rect 2823 28101 2832 28135
rect 2780 28092 2832 28101
rect 3332 28092 3384 28144
rect 4160 28092 4212 28144
rect 4252 28092 4304 28144
rect 4528 28135 4580 28144
rect 4528 28101 4537 28135
rect 4537 28101 4571 28135
rect 4571 28101 4580 28135
rect 4528 28092 4580 28101
rect 756 28024 808 28076
rect 1676 28024 1728 28076
rect 2320 28067 2372 28076
rect 2320 28033 2329 28067
rect 2329 28033 2363 28067
rect 2363 28033 2372 28067
rect 2320 28024 2372 28033
rect 2964 28024 3016 28076
rect 3516 28067 3568 28076
rect 3516 28033 3525 28067
rect 3525 28033 3559 28067
rect 3559 28033 3568 28067
rect 5356 28092 5408 28144
rect 9956 28160 10008 28212
rect 3516 28024 3568 28033
rect 4804 28067 4856 28076
rect 4804 28033 4813 28067
rect 4813 28033 4847 28067
rect 4847 28033 4856 28067
rect 4804 28024 4856 28033
rect 5448 28024 5500 28076
rect 7656 28024 7708 28076
rect 9588 28024 9640 28076
rect 3240 27956 3292 28008
rect 4988 27956 5040 28008
rect 5632 27956 5684 28008
rect 6276 27956 6328 28008
rect 7196 27956 7248 28008
rect 9864 27956 9916 28008
rect 14924 28160 14976 28212
rect 16672 28160 16724 28212
rect 11152 28092 11204 28144
rect 11704 28092 11756 28144
rect 14740 28092 14792 28144
rect 19616 28160 19668 28212
rect 17316 28092 17368 28144
rect 17776 28092 17828 28144
rect 10416 28024 10468 28076
rect 11060 28024 11112 28076
rect 11336 28024 11388 28076
rect 13176 28024 13228 28076
rect 14004 28067 14056 28076
rect 14004 28033 14013 28067
rect 14013 28033 14047 28067
rect 14047 28033 14056 28067
rect 14004 28024 14056 28033
rect 7288 27888 7340 27940
rect 6828 27820 6880 27872
rect 12624 27956 12676 28008
rect 12992 27999 13044 28008
rect 12992 27965 13001 27999
rect 13001 27965 13035 27999
rect 13035 27965 13044 27999
rect 12992 27956 13044 27965
rect 11704 27888 11756 27940
rect 13820 27999 13872 28008
rect 13820 27965 13854 27999
rect 13854 27965 13872 27999
rect 13820 27956 13872 27965
rect 14372 27956 14424 28008
rect 14648 27956 14700 28008
rect 17684 28024 17736 28076
rect 19340 28092 19392 28144
rect 19432 28092 19484 28144
rect 20996 28160 21048 28212
rect 21088 28160 21140 28212
rect 17960 28024 18012 28076
rect 18604 28024 18656 28076
rect 15200 27999 15252 28008
rect 15200 27965 15209 27999
rect 15209 27965 15243 27999
rect 15243 27965 15252 27999
rect 15200 27956 15252 27965
rect 22192 28092 22244 28144
rect 22928 28092 22980 28144
rect 19432 27999 19484 28008
rect 19432 27965 19441 27999
rect 19441 27965 19475 27999
rect 19475 27965 19484 27999
rect 19432 27956 19484 27965
rect 20720 27956 20772 28008
rect 22100 28024 22152 28076
rect 22836 28067 22888 28076
rect 22836 28033 22845 28067
rect 22845 28033 22879 28067
rect 22879 28033 22888 28067
rect 22836 28024 22888 28033
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 11060 27863 11112 27872
rect 11060 27829 11069 27863
rect 11069 27829 11103 27863
rect 11103 27829 11112 27863
rect 11060 27820 11112 27829
rect 11428 27820 11480 27872
rect 11980 27820 12032 27872
rect 12992 27820 13044 27872
rect 13728 27820 13780 27872
rect 13912 27820 13964 27872
rect 14648 27863 14700 27872
rect 14648 27829 14657 27863
rect 14657 27829 14691 27863
rect 14691 27829 14700 27863
rect 14648 27820 14700 27829
rect 14740 27820 14792 27872
rect 14924 27820 14976 27872
rect 19616 27820 19668 27872
rect 20812 27863 20864 27872
rect 20812 27829 20821 27863
rect 20821 27829 20855 27863
rect 20855 27829 20864 27863
rect 20812 27820 20864 27829
rect 22560 27888 22612 27940
rect 22468 27820 22520 27872
rect 23020 27820 23072 27872
rect 23756 27863 23808 27872
rect 23756 27829 23765 27863
rect 23765 27829 23799 27863
rect 23799 27829 23808 27863
rect 23756 27820 23808 27829
rect 24400 27863 24452 27872
rect 24400 27829 24409 27863
rect 24409 27829 24443 27863
rect 24443 27829 24452 27863
rect 24400 27820 24452 27829
rect 3917 27718 3969 27770
rect 3981 27718 4033 27770
rect 4045 27718 4097 27770
rect 4109 27718 4161 27770
rect 4173 27718 4225 27770
rect 9851 27718 9903 27770
rect 9915 27718 9967 27770
rect 9979 27718 10031 27770
rect 10043 27718 10095 27770
rect 10107 27718 10159 27770
rect 15785 27718 15837 27770
rect 15849 27718 15901 27770
rect 15913 27718 15965 27770
rect 15977 27718 16029 27770
rect 16041 27718 16093 27770
rect 21719 27718 21771 27770
rect 21783 27718 21835 27770
rect 21847 27718 21899 27770
rect 21911 27718 21963 27770
rect 21975 27718 22027 27770
rect 480 27616 532 27668
rect 3332 27616 3384 27668
rect 4528 27616 4580 27668
rect 6368 27616 6420 27668
rect 10324 27616 10376 27668
rect 1400 27523 1452 27532
rect 1400 27489 1409 27523
rect 1409 27489 1443 27523
rect 1443 27489 1452 27523
rect 1400 27480 1452 27489
rect 7840 27548 7892 27600
rect 8024 27548 8076 27600
rect 10416 27591 10468 27600
rect 10416 27557 10425 27591
rect 10425 27557 10459 27591
rect 10459 27557 10468 27591
rect 10416 27548 10468 27557
rect 8760 27480 8812 27532
rect 1584 27412 1636 27464
rect 1216 27344 1268 27396
rect 4436 27412 4488 27464
rect 4988 27412 5040 27464
rect 6552 27412 6604 27464
rect 6828 27412 6880 27464
rect 7104 27455 7156 27464
rect 7104 27421 7113 27455
rect 7113 27421 7147 27455
rect 7147 27421 7156 27455
rect 7104 27412 7156 27421
rect 7840 27412 7892 27464
rect 9680 27412 9732 27464
rect 2044 27276 2096 27328
rect 2964 27319 3016 27328
rect 2964 27285 2973 27319
rect 2973 27285 3007 27319
rect 3007 27285 3016 27319
rect 2964 27276 3016 27285
rect 4988 27276 5040 27328
rect 6276 27276 6328 27328
rect 6368 27319 6420 27328
rect 6368 27285 6377 27319
rect 6377 27285 6411 27319
rect 6411 27285 6420 27319
rect 6368 27276 6420 27285
rect 6460 27276 6512 27328
rect 6828 27276 6880 27328
rect 7472 27319 7524 27328
rect 7472 27285 7481 27319
rect 7481 27285 7515 27319
rect 7515 27285 7524 27319
rect 7472 27276 7524 27285
rect 7656 27319 7708 27328
rect 7656 27285 7665 27319
rect 7665 27285 7699 27319
rect 7699 27285 7708 27319
rect 7656 27276 7708 27285
rect 9220 27276 9272 27328
rect 9404 27387 9456 27396
rect 9404 27353 9413 27387
rect 9413 27353 9447 27387
rect 9447 27353 9456 27387
rect 9404 27344 9456 27353
rect 9588 27344 9640 27396
rect 9864 27387 9916 27396
rect 9864 27353 9873 27387
rect 9873 27353 9907 27387
rect 9907 27353 9916 27387
rect 9864 27344 9916 27353
rect 11428 27412 11480 27464
rect 11520 27455 11572 27464
rect 11520 27421 11529 27455
rect 11529 27421 11563 27455
rect 11563 27421 11572 27455
rect 11520 27412 11572 27421
rect 11796 27391 11821 27396
rect 11821 27391 11848 27396
rect 11796 27344 11848 27391
rect 12072 27344 12124 27396
rect 15292 27548 15344 27600
rect 12348 27480 12400 27532
rect 12532 27480 12584 27532
rect 15844 27480 15896 27532
rect 22468 27616 22520 27668
rect 22836 27616 22888 27668
rect 23020 27616 23072 27668
rect 20720 27548 20772 27600
rect 20812 27548 20864 27600
rect 21088 27548 21140 27600
rect 14004 27412 14056 27464
rect 14648 27412 14700 27464
rect 15292 27412 15344 27464
rect 15568 27412 15620 27464
rect 16488 27455 16540 27464
rect 16488 27421 16513 27455
rect 16513 27421 16540 27455
rect 12256 27276 12308 27328
rect 13820 27344 13872 27396
rect 16488 27412 16540 27421
rect 12716 27276 12768 27328
rect 13636 27276 13688 27328
rect 14924 27276 14976 27328
rect 15016 27319 15068 27328
rect 15016 27285 15025 27319
rect 15025 27285 15059 27319
rect 15059 27285 15068 27319
rect 15016 27276 15068 27285
rect 15200 27276 15252 27328
rect 19616 27412 19668 27464
rect 23940 27616 23992 27668
rect 21180 27455 21232 27464
rect 21180 27421 21189 27455
rect 21189 27421 21223 27455
rect 21223 27421 21232 27455
rect 21180 27412 21232 27421
rect 23572 27480 23624 27532
rect 22008 27344 22060 27396
rect 22836 27344 22888 27396
rect 16580 27276 16632 27328
rect 17224 27319 17276 27328
rect 17224 27285 17233 27319
rect 17233 27285 17267 27319
rect 17267 27285 17276 27319
rect 17224 27276 17276 27285
rect 17408 27276 17460 27328
rect 17868 27276 17920 27328
rect 19340 27276 19392 27328
rect 21180 27276 21232 27328
rect 22928 27319 22980 27328
rect 22928 27285 22937 27319
rect 22937 27285 22971 27319
rect 22971 27285 22980 27319
rect 22928 27276 22980 27285
rect 23020 27276 23072 27328
rect 25136 27276 25188 27328
rect 6884 27174 6936 27226
rect 6948 27174 7000 27226
rect 7012 27174 7064 27226
rect 7076 27174 7128 27226
rect 7140 27174 7192 27226
rect 12818 27174 12870 27226
rect 12882 27174 12934 27226
rect 12946 27174 12998 27226
rect 13010 27174 13062 27226
rect 13074 27174 13126 27226
rect 18752 27174 18804 27226
rect 18816 27174 18868 27226
rect 18880 27174 18932 27226
rect 18944 27174 18996 27226
rect 19008 27174 19060 27226
rect 24686 27174 24738 27226
rect 24750 27174 24802 27226
rect 24814 27174 24866 27226
rect 24878 27174 24930 27226
rect 24942 27174 24994 27226
rect 1676 27072 1728 27124
rect 2780 27072 2832 27124
rect 2964 27072 3016 27124
rect 3332 27115 3384 27124
rect 3332 27081 3341 27115
rect 3341 27081 3375 27115
rect 3375 27081 3384 27115
rect 3332 27072 3384 27081
rect 2596 27004 2648 27056
rect 2412 26979 2464 26988
rect 2412 26945 2421 26979
rect 2421 26945 2455 26979
rect 2455 26945 2464 26979
rect 2412 26936 2464 26945
rect 4528 27004 4580 27056
rect 2044 26868 2096 26920
rect 3792 26936 3844 26988
rect 4988 27004 5040 27056
rect 5448 27072 5500 27124
rect 8116 27072 8168 27124
rect 8484 27072 8536 27124
rect 8760 27115 8812 27124
rect 8760 27081 8769 27115
rect 8769 27081 8803 27115
rect 8803 27081 8812 27115
rect 8760 27072 8812 27081
rect 9404 27072 9456 27124
rect 10508 27072 10560 27124
rect 11612 27072 11664 27124
rect 12532 27072 12584 27124
rect 12624 27004 12676 27056
rect 13636 27072 13688 27124
rect 14004 27072 14056 27124
rect 8116 26936 8168 26988
rect 19340 27072 19392 27124
rect 13820 26979 13872 26988
rect 13820 26945 13854 26979
rect 13854 26945 13872 26979
rect 15200 27004 15252 27056
rect 15844 27004 15896 27056
rect 19800 27004 19852 27056
rect 21088 27004 21140 27056
rect 21640 27004 21692 27056
rect 22836 27115 22888 27124
rect 22836 27081 22845 27115
rect 22845 27081 22879 27115
rect 22879 27081 22888 27115
rect 22836 27072 22888 27081
rect 23020 27072 23072 27124
rect 23572 27072 23624 27124
rect 23756 27072 23808 27124
rect 13820 26936 13872 26945
rect 14924 26936 14976 26988
rect 3608 26868 3660 26920
rect 4528 26911 4580 26920
rect 4528 26877 4537 26911
rect 4537 26877 4571 26911
rect 4571 26877 4580 26911
rect 4528 26868 4580 26877
rect 7748 26911 7800 26920
rect 7748 26877 7757 26911
rect 7757 26877 7791 26911
rect 7791 26877 7800 26911
rect 7748 26868 7800 26877
rect 9220 26868 9272 26920
rect 9772 26868 9824 26920
rect 9864 26868 9916 26920
rect 12256 26868 12308 26920
rect 13360 26868 13412 26920
rect 13452 26911 13504 26920
rect 13452 26877 13461 26911
rect 13461 26877 13495 26911
rect 13495 26877 13504 26911
rect 13452 26868 13504 26877
rect 12900 26800 12952 26852
rect 16764 26936 16816 26988
rect 17868 26979 17920 26988
rect 17868 26945 17877 26979
rect 17877 26945 17911 26979
rect 17911 26945 17920 26979
rect 17868 26936 17920 26945
rect 20076 26936 20128 26988
rect 23020 26936 23072 26988
rect 23756 26979 23808 26988
rect 23756 26945 23765 26979
rect 23765 26945 23799 26979
rect 23799 26945 23808 26979
rect 23756 26936 23808 26945
rect 16580 26868 16632 26920
rect 16948 26868 17000 26920
rect 17224 26868 17276 26920
rect 3240 26732 3292 26784
rect 8024 26732 8076 26784
rect 9312 26732 9364 26784
rect 17132 26800 17184 26852
rect 17776 26868 17828 26920
rect 21088 26868 21140 26920
rect 21548 26868 21600 26920
rect 24860 26936 24912 26988
rect 25596 26936 25648 26988
rect 19432 26732 19484 26784
rect 22928 26732 22980 26784
rect 24124 26732 24176 26784
rect 24400 26775 24452 26784
rect 24400 26741 24409 26775
rect 24409 26741 24443 26775
rect 24443 26741 24452 26775
rect 24400 26732 24452 26741
rect 3917 26630 3969 26682
rect 3981 26630 4033 26682
rect 4045 26630 4097 26682
rect 4109 26630 4161 26682
rect 4173 26630 4225 26682
rect 9851 26630 9903 26682
rect 9915 26630 9967 26682
rect 9979 26630 10031 26682
rect 10043 26630 10095 26682
rect 10107 26630 10159 26682
rect 15785 26630 15837 26682
rect 15849 26630 15901 26682
rect 15913 26630 15965 26682
rect 15977 26630 16029 26682
rect 16041 26630 16093 26682
rect 21719 26630 21771 26682
rect 21783 26630 21835 26682
rect 21847 26630 21899 26682
rect 21911 26630 21963 26682
rect 21975 26630 22027 26682
rect 2412 26528 2464 26580
rect 3516 26528 3568 26580
rect 8668 26528 8720 26580
rect 1400 26392 1452 26444
rect 2872 26324 2924 26376
rect 3516 26392 3568 26444
rect 4252 26392 4304 26444
rect 4528 26392 4580 26444
rect 6552 26435 6604 26444
rect 6552 26401 6561 26435
rect 6561 26401 6595 26435
rect 6595 26401 6604 26435
rect 6552 26392 6604 26401
rect 9680 26460 9732 26512
rect 9956 26392 10008 26444
rect 10968 26528 11020 26580
rect 3240 26256 3292 26308
rect 3424 26367 3476 26376
rect 3424 26333 3433 26367
rect 3433 26333 3467 26367
rect 3467 26333 3476 26367
rect 3424 26324 3476 26333
rect 3792 26367 3844 26376
rect 3792 26333 3801 26367
rect 3801 26333 3835 26367
rect 3835 26333 3844 26367
rect 3792 26324 3844 26333
rect 6736 26324 6788 26376
rect 7472 26324 7524 26376
rect 8208 26324 8260 26376
rect 9312 26324 9364 26376
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 10416 26367 10468 26376
rect 10416 26333 10425 26367
rect 10425 26333 10459 26367
rect 10459 26333 10468 26367
rect 10416 26324 10468 26333
rect 11060 26392 11112 26444
rect 11796 26367 11848 26376
rect 11796 26333 11805 26367
rect 11805 26333 11839 26367
rect 11839 26333 11848 26367
rect 11796 26324 11848 26333
rect 11888 26367 11940 26376
rect 11888 26333 11897 26367
rect 11897 26333 11931 26367
rect 11931 26333 11940 26367
rect 11888 26324 11940 26333
rect 13912 26324 13964 26376
rect 14096 26324 14148 26376
rect 15200 26367 15252 26376
rect 15200 26333 15207 26367
rect 15207 26333 15241 26367
rect 15241 26333 15252 26367
rect 16304 26528 16356 26580
rect 19708 26528 19760 26580
rect 23756 26528 23808 26580
rect 15936 26503 15988 26512
rect 15936 26469 15945 26503
rect 15945 26469 15979 26503
rect 15979 26469 15988 26503
rect 15936 26460 15988 26469
rect 19524 26460 19576 26512
rect 20444 26460 20496 26512
rect 17684 26435 17736 26444
rect 17684 26401 17693 26435
rect 17693 26401 17727 26435
rect 17727 26401 17736 26435
rect 17684 26392 17736 26401
rect 23572 26460 23624 26512
rect 24492 26460 24544 26512
rect 24860 26460 24912 26512
rect 15200 26324 15252 26333
rect 15660 26324 15712 26376
rect 5356 26188 5408 26240
rect 5816 26188 5868 26240
rect 7656 26188 7708 26240
rect 7748 26188 7800 26240
rect 8300 26188 8352 26240
rect 12164 26256 12216 26308
rect 10968 26188 11020 26240
rect 11428 26188 11480 26240
rect 12624 26231 12676 26240
rect 12624 26197 12633 26231
rect 12633 26197 12667 26231
rect 12667 26197 12676 26231
rect 12624 26188 12676 26197
rect 16856 26299 16908 26308
rect 16856 26265 16865 26299
rect 16865 26265 16899 26299
rect 16899 26265 16908 26299
rect 16856 26256 16908 26265
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 20536 26324 20588 26376
rect 20720 26324 20772 26376
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 23572 26324 23624 26376
rect 19616 26256 19668 26308
rect 25136 26256 25188 26308
rect 12900 26188 12952 26240
rect 13268 26188 13320 26240
rect 14832 26188 14884 26240
rect 16120 26188 16172 26240
rect 19248 26231 19300 26240
rect 19248 26197 19257 26231
rect 19257 26197 19291 26231
rect 19291 26197 19300 26231
rect 19248 26188 19300 26197
rect 23664 26231 23716 26240
rect 23664 26197 23673 26231
rect 23673 26197 23707 26231
rect 23707 26197 23716 26231
rect 23664 26188 23716 26197
rect 6884 26086 6936 26138
rect 6948 26086 7000 26138
rect 7012 26086 7064 26138
rect 7076 26086 7128 26138
rect 7140 26086 7192 26138
rect 12818 26086 12870 26138
rect 12882 26086 12934 26138
rect 12946 26086 12998 26138
rect 13010 26086 13062 26138
rect 13074 26086 13126 26138
rect 18752 26086 18804 26138
rect 18816 26086 18868 26138
rect 18880 26086 18932 26138
rect 18944 26086 18996 26138
rect 19008 26086 19060 26138
rect 24686 26086 24738 26138
rect 24750 26086 24802 26138
rect 24814 26086 24866 26138
rect 24878 26086 24930 26138
rect 24942 26086 24994 26138
rect 2412 25984 2464 26036
rect 1308 25916 1360 25968
rect 1400 25848 1452 25900
rect 2780 25848 2832 25900
rect 6000 25916 6052 25968
rect 4252 25848 4304 25900
rect 6276 25848 6328 25900
rect 7288 25916 7340 25968
rect 7656 25916 7708 25968
rect 7840 25959 7892 25968
rect 7840 25925 7849 25959
rect 7849 25925 7883 25959
rect 7883 25925 7892 25959
rect 7840 25916 7892 25925
rect 8208 25959 8260 25968
rect 8208 25925 8217 25959
rect 8217 25925 8251 25959
rect 8251 25925 8260 25959
rect 8208 25916 8260 25925
rect 7748 25848 7800 25900
rect 1216 25644 1268 25696
rect 2228 25644 2280 25696
rect 2596 25644 2648 25696
rect 2780 25644 2832 25696
rect 3148 25644 3200 25696
rect 3700 25644 3752 25696
rect 4436 25687 4488 25696
rect 4436 25653 4445 25687
rect 4445 25653 4479 25687
rect 4479 25653 4488 25687
rect 4436 25644 4488 25653
rect 7564 25780 7616 25832
rect 5264 25644 5316 25696
rect 5816 25687 5868 25696
rect 5816 25653 5825 25687
rect 5825 25653 5859 25687
rect 5859 25653 5868 25687
rect 5816 25644 5868 25653
rect 8392 25687 8444 25696
rect 8392 25653 8401 25687
rect 8401 25653 8435 25687
rect 8435 25653 8444 25687
rect 8392 25644 8444 25653
rect 8760 25780 8812 25832
rect 11612 25984 11664 26036
rect 11796 25984 11848 26036
rect 11888 25984 11940 26036
rect 14832 25984 14884 26036
rect 15016 25984 15068 26036
rect 15660 26027 15712 26036
rect 15660 25993 15669 26027
rect 15669 25993 15703 26027
rect 15703 25993 15712 26027
rect 15660 25984 15712 25993
rect 15936 25984 15988 26036
rect 16856 25984 16908 26036
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 12256 25848 12308 25900
rect 9588 25780 9640 25832
rect 9772 25780 9824 25832
rect 10048 25823 10100 25832
rect 10048 25789 10082 25823
rect 10082 25789 10100 25823
rect 10048 25780 10100 25789
rect 10416 25780 10468 25832
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 14004 25891 14056 25900
rect 14004 25857 14013 25891
rect 14013 25857 14047 25891
rect 14047 25857 14056 25891
rect 14004 25848 14056 25857
rect 14280 25891 14332 25900
rect 14280 25857 14289 25891
rect 14289 25857 14323 25891
rect 14323 25857 14332 25891
rect 14280 25848 14332 25857
rect 17132 25916 17184 25968
rect 20720 25916 20772 25968
rect 23572 25984 23624 26036
rect 24308 25984 24360 26036
rect 9680 25755 9732 25764
rect 9680 25721 9689 25755
rect 9689 25721 9723 25755
rect 9723 25721 9732 25755
rect 9680 25712 9732 25721
rect 10692 25712 10744 25764
rect 12992 25712 13044 25764
rect 13728 25823 13780 25832
rect 13728 25789 13737 25823
rect 13737 25789 13771 25823
rect 13771 25789 13780 25823
rect 13728 25780 13780 25789
rect 17960 25848 18012 25900
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 13268 25644 13320 25696
rect 13452 25644 13504 25696
rect 16120 25780 16172 25832
rect 16488 25780 16540 25832
rect 15660 25712 15712 25764
rect 16672 25712 16724 25764
rect 14832 25644 14884 25696
rect 17408 25644 17460 25696
rect 20352 25712 20404 25764
rect 21364 25891 21416 25900
rect 21364 25857 21373 25891
rect 21373 25857 21407 25891
rect 21407 25857 21416 25891
rect 21364 25848 21416 25857
rect 21548 25891 21600 25900
rect 21548 25857 21557 25891
rect 21557 25857 21591 25891
rect 21591 25857 21600 25891
rect 21548 25848 21600 25857
rect 22100 25848 22152 25900
rect 23848 25916 23900 25968
rect 23572 25848 23624 25900
rect 23388 25780 23440 25832
rect 19432 25644 19484 25696
rect 19984 25644 20036 25696
rect 20076 25687 20128 25696
rect 20076 25653 20085 25687
rect 20085 25653 20119 25687
rect 20119 25653 20128 25687
rect 20076 25644 20128 25653
rect 21088 25644 21140 25696
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 23112 25687 23164 25696
rect 23112 25653 23121 25687
rect 23121 25653 23155 25687
rect 23155 25653 23164 25687
rect 23112 25644 23164 25653
rect 24400 25687 24452 25696
rect 24400 25653 24409 25687
rect 24409 25653 24443 25687
rect 24443 25653 24452 25687
rect 24400 25644 24452 25653
rect 3917 25542 3969 25594
rect 3981 25542 4033 25594
rect 4045 25542 4097 25594
rect 4109 25542 4161 25594
rect 4173 25542 4225 25594
rect 9851 25542 9903 25594
rect 9915 25542 9967 25594
rect 9979 25542 10031 25594
rect 10043 25542 10095 25594
rect 10107 25542 10159 25594
rect 15785 25542 15837 25594
rect 15849 25542 15901 25594
rect 15913 25542 15965 25594
rect 15977 25542 16029 25594
rect 16041 25542 16093 25594
rect 21719 25542 21771 25594
rect 21783 25542 21835 25594
rect 21847 25542 21899 25594
rect 21911 25542 21963 25594
rect 21975 25542 22027 25594
rect 2228 25440 2280 25492
rect 7748 25440 7800 25492
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 1676 25279 1728 25288
rect 1676 25245 1685 25279
rect 1685 25245 1719 25279
rect 1719 25245 1728 25279
rect 1676 25236 1728 25245
rect 2044 25236 2096 25288
rect 2136 25279 2188 25288
rect 2136 25245 2145 25279
rect 2145 25245 2179 25279
rect 2179 25245 2188 25279
rect 2136 25236 2188 25245
rect 3700 25372 3752 25424
rect 10416 25440 10468 25492
rect 11152 25440 11204 25492
rect 12992 25440 13044 25492
rect 16580 25440 16632 25492
rect 16856 25440 16908 25492
rect 5264 25304 5316 25356
rect 2320 25168 2372 25220
rect 3516 25236 3568 25288
rect 5080 25236 5132 25288
rect 1860 25143 1912 25152
rect 1860 25109 1869 25143
rect 1869 25109 1903 25143
rect 1903 25109 1912 25143
rect 1860 25100 1912 25109
rect 3700 25100 3752 25152
rect 3884 25100 3936 25152
rect 4068 25100 4120 25152
rect 4436 25168 4488 25220
rect 6184 25304 6236 25356
rect 6552 25304 6604 25356
rect 7012 25236 7064 25288
rect 8024 25236 8076 25288
rect 12532 25304 12584 25356
rect 15384 25372 15436 25424
rect 16488 25372 16540 25424
rect 16764 25304 16816 25356
rect 17316 25347 17368 25356
rect 17316 25313 17325 25347
rect 17325 25313 17359 25347
rect 17359 25313 17368 25347
rect 17316 25304 17368 25313
rect 20076 25440 20128 25492
rect 20352 25440 20404 25492
rect 21364 25483 21416 25492
rect 21364 25449 21373 25483
rect 21373 25449 21407 25483
rect 21407 25449 21416 25483
rect 21364 25440 21416 25449
rect 23112 25440 23164 25492
rect 23572 25440 23624 25492
rect 23664 25440 23716 25492
rect 19524 25372 19576 25424
rect 8484 25236 8536 25288
rect 10324 25236 10376 25288
rect 11060 25236 11112 25288
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 12716 25236 12768 25288
rect 17592 25279 17644 25288
rect 17592 25245 17601 25279
rect 17601 25245 17635 25279
rect 17635 25245 17644 25279
rect 17592 25236 17644 25245
rect 17868 25279 17920 25288
rect 17868 25245 17877 25279
rect 17877 25245 17911 25279
rect 17911 25245 17920 25279
rect 17868 25236 17920 25245
rect 19248 25279 19300 25288
rect 19248 25245 19257 25279
rect 19257 25245 19291 25279
rect 19291 25245 19300 25279
rect 19248 25236 19300 25245
rect 19984 25304 20036 25356
rect 23480 25304 23532 25356
rect 20076 25236 20128 25288
rect 5264 25143 5316 25152
rect 5264 25109 5273 25143
rect 5273 25109 5307 25143
rect 5307 25109 5316 25143
rect 5264 25100 5316 25109
rect 6368 25100 6420 25152
rect 8760 25168 8812 25220
rect 7288 25100 7340 25152
rect 9772 25100 9824 25152
rect 11060 25100 11112 25152
rect 11336 25100 11388 25152
rect 11612 25168 11664 25220
rect 11888 25100 11940 25152
rect 12164 25211 12216 25220
rect 12164 25177 12173 25211
rect 12173 25177 12207 25211
rect 12207 25177 12216 25211
rect 12164 25168 12216 25177
rect 12624 25100 12676 25152
rect 19156 25168 19208 25220
rect 21180 25236 21232 25288
rect 22560 25236 22612 25288
rect 21732 25168 21784 25220
rect 22100 25211 22152 25220
rect 22100 25177 22134 25211
rect 22134 25177 22152 25211
rect 22100 25168 22152 25177
rect 25136 25168 25188 25220
rect 19432 25100 19484 25152
rect 19708 25100 19760 25152
rect 22560 25100 22612 25152
rect 23756 25100 23808 25152
rect 6884 24998 6936 25050
rect 6948 24998 7000 25050
rect 7012 24998 7064 25050
rect 7076 24998 7128 25050
rect 7140 24998 7192 25050
rect 12818 24998 12870 25050
rect 12882 24998 12934 25050
rect 12946 24998 12998 25050
rect 13010 24998 13062 25050
rect 13074 24998 13126 25050
rect 18752 24998 18804 25050
rect 18816 24998 18868 25050
rect 18880 24998 18932 25050
rect 18944 24998 18996 25050
rect 19008 24998 19060 25050
rect 24686 24998 24738 25050
rect 24750 24998 24802 25050
rect 24814 24998 24866 25050
rect 24878 24998 24930 25050
rect 24942 24998 24994 25050
rect 1124 24896 1176 24948
rect 1308 24896 1360 24948
rect 1584 24939 1636 24948
rect 1584 24905 1593 24939
rect 1593 24905 1627 24939
rect 1627 24905 1636 24939
rect 1584 24896 1636 24905
rect 1952 24896 2004 24948
rect 1032 24828 1084 24880
rect 3700 24896 3752 24948
rect 4712 24896 4764 24948
rect 4988 24896 5040 24948
rect 5264 24896 5316 24948
rect 756 24760 808 24812
rect 1584 24760 1636 24812
rect 1124 24692 1176 24744
rect 3056 24760 3108 24812
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3283 24803
rect 3283 24769 3292 24803
rect 3240 24760 3292 24769
rect 3884 24828 3936 24880
rect 6276 24828 6328 24880
rect 3424 24760 3476 24812
rect 6920 24760 6972 24812
rect 8392 24828 8444 24880
rect 17132 24828 17184 24880
rect 17316 24896 17368 24948
rect 19708 24896 19760 24948
rect 19984 24896 20036 24948
rect 17960 24828 18012 24880
rect 8668 24760 8720 24812
rect 8852 24760 8904 24812
rect 11520 24760 11572 24812
rect 11612 24760 11664 24812
rect 13636 24760 13688 24812
rect 13912 24760 13964 24812
rect 15476 24760 15528 24812
rect 17408 24760 17460 24812
rect 17500 24760 17552 24812
rect 19432 24828 19484 24880
rect 21548 24896 21600 24948
rect 23480 24939 23532 24948
rect 23480 24905 23489 24939
rect 23489 24905 23523 24939
rect 23523 24905 23532 24939
rect 23480 24896 23532 24905
rect 20168 24803 20220 24812
rect 20168 24769 20191 24803
rect 20191 24769 20220 24803
rect 20168 24760 20220 24769
rect 21364 24803 21416 24812
rect 21364 24769 21373 24803
rect 21373 24769 21407 24803
rect 21407 24769 21416 24803
rect 21364 24760 21416 24769
rect 3516 24692 3568 24744
rect 4712 24692 4764 24744
rect 5080 24692 5132 24744
rect 5264 24735 5316 24744
rect 5264 24701 5273 24735
rect 5273 24701 5307 24735
rect 5307 24701 5316 24735
rect 5264 24692 5316 24701
rect 5448 24692 5500 24744
rect 6368 24692 6420 24744
rect 8208 24692 8260 24744
rect 8484 24735 8536 24744
rect 8484 24701 8493 24735
rect 8493 24701 8527 24735
rect 8527 24701 8536 24735
rect 8484 24692 8536 24701
rect 11152 24692 11204 24744
rect 12164 24735 12216 24744
rect 12164 24701 12173 24735
rect 12173 24701 12207 24735
rect 12207 24701 12216 24735
rect 12164 24692 12216 24701
rect 14280 24692 14332 24744
rect 16672 24735 16724 24744
rect 16672 24701 16681 24735
rect 16681 24701 16715 24735
rect 16715 24701 16724 24735
rect 16672 24692 16724 24701
rect 2320 24624 2372 24676
rect 4068 24624 4120 24676
rect 4620 24624 4672 24676
rect 1768 24556 1820 24608
rect 2780 24556 2832 24608
rect 4896 24556 4948 24608
rect 6552 24624 6604 24676
rect 7932 24624 7984 24676
rect 9680 24624 9732 24676
rect 10324 24624 10376 24676
rect 11888 24624 11940 24676
rect 5724 24556 5776 24608
rect 6276 24556 6328 24608
rect 17868 24624 17920 24676
rect 13176 24599 13228 24608
rect 13176 24565 13185 24599
rect 13185 24565 13219 24599
rect 13219 24565 13228 24599
rect 13176 24556 13228 24565
rect 14464 24556 14516 24608
rect 15384 24556 15436 24608
rect 16120 24556 16172 24608
rect 16580 24556 16632 24608
rect 17776 24556 17828 24608
rect 21548 24692 21600 24744
rect 22376 24760 22428 24812
rect 24216 24760 24268 24812
rect 22192 24692 22244 24744
rect 20628 24556 20680 24608
rect 21180 24556 21232 24608
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 24308 24624 24360 24676
rect 24400 24599 24452 24608
rect 24400 24565 24409 24599
rect 24409 24565 24443 24599
rect 24443 24565 24452 24599
rect 24400 24556 24452 24565
rect 3917 24454 3969 24506
rect 3981 24454 4033 24506
rect 4045 24454 4097 24506
rect 4109 24454 4161 24506
rect 4173 24454 4225 24506
rect 9851 24454 9903 24506
rect 9915 24454 9967 24506
rect 9979 24454 10031 24506
rect 10043 24454 10095 24506
rect 10107 24454 10159 24506
rect 15785 24454 15837 24506
rect 15849 24454 15901 24506
rect 15913 24454 15965 24506
rect 15977 24454 16029 24506
rect 16041 24454 16093 24506
rect 21719 24454 21771 24506
rect 21783 24454 21835 24506
rect 21847 24454 21899 24506
rect 21911 24454 21963 24506
rect 21975 24454 22027 24506
rect 2780 24352 2832 24404
rect 2872 24395 2924 24404
rect 2872 24361 2881 24395
rect 2881 24361 2915 24395
rect 2915 24361 2924 24395
rect 2872 24352 2924 24361
rect 3056 24352 3108 24404
rect 6920 24352 6972 24404
rect 2412 24216 2464 24268
rect 5448 24284 5500 24336
rect 5816 24327 5868 24336
rect 5816 24293 5825 24327
rect 5825 24293 5859 24327
rect 5859 24293 5868 24327
rect 5816 24284 5868 24293
rect 4160 24216 4212 24268
rect 4528 24216 4580 24268
rect 4804 24216 4856 24268
rect 5264 24216 5316 24268
rect 6368 24259 6420 24268
rect 6368 24225 6377 24259
rect 6377 24225 6411 24259
rect 6411 24225 6420 24259
rect 6368 24216 6420 24225
rect 2504 24148 2556 24200
rect 1492 24080 1544 24132
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 3424 24148 3476 24200
rect 3700 24148 3752 24200
rect 4988 24148 5040 24200
rect 6092 24191 6144 24200
rect 6092 24157 6101 24191
rect 6101 24157 6135 24191
rect 6135 24157 6144 24191
rect 6092 24148 6144 24157
rect 9036 24352 9088 24404
rect 10324 24352 10376 24404
rect 8392 24284 8444 24336
rect 9772 24216 9824 24268
rect 10232 24216 10284 24268
rect 10968 24352 11020 24404
rect 11520 24352 11572 24404
rect 16580 24352 16632 24404
rect 14096 24284 14148 24336
rect 12164 24216 12216 24268
rect 13544 24216 13596 24268
rect 14924 24216 14976 24268
rect 15108 24216 15160 24268
rect 15292 24216 15344 24268
rect 15660 24259 15712 24268
rect 15660 24225 15669 24259
rect 15669 24225 15703 24259
rect 15703 24225 15712 24259
rect 15660 24216 15712 24225
rect 16764 24216 16816 24268
rect 8300 24148 8352 24200
rect 9588 24148 9640 24200
rect 10876 24191 10928 24200
rect 10876 24157 10883 24191
rect 10883 24157 10917 24191
rect 10917 24157 10928 24191
rect 10876 24148 10928 24157
rect 11888 24148 11940 24200
rect 4436 24080 4488 24132
rect 4620 24080 4672 24132
rect 5264 24080 5316 24132
rect 2596 24012 2648 24064
rect 4160 24012 4212 24064
rect 10324 24080 10376 24132
rect 12256 24080 12308 24132
rect 14464 24080 14516 24132
rect 15936 24191 15988 24200
rect 15936 24157 15945 24191
rect 15945 24157 15979 24191
rect 15979 24157 15988 24191
rect 15936 24148 15988 24157
rect 16028 24191 16080 24200
rect 16028 24157 16062 24191
rect 16062 24157 16080 24191
rect 16028 24148 16080 24157
rect 7564 24055 7616 24064
rect 7564 24021 7573 24055
rect 7573 24021 7607 24055
rect 7607 24021 7616 24055
rect 7564 24012 7616 24021
rect 7748 24055 7800 24064
rect 7748 24021 7757 24055
rect 7757 24021 7791 24055
rect 7791 24021 7800 24055
rect 7748 24012 7800 24021
rect 9680 24012 9732 24064
rect 11244 24012 11296 24064
rect 13820 24012 13872 24064
rect 14556 24012 14608 24064
rect 14924 24012 14976 24064
rect 17500 24080 17552 24132
rect 19248 24148 19300 24200
rect 17408 24012 17460 24064
rect 19616 24012 19668 24064
rect 21456 24352 21508 24404
rect 22376 24352 22428 24404
rect 22652 24352 22704 24404
rect 23388 24395 23440 24404
rect 23388 24361 23397 24395
rect 23397 24361 23431 24395
rect 23431 24361 23440 24395
rect 23388 24352 23440 24361
rect 21088 24216 21140 24268
rect 20168 24148 20220 24200
rect 22468 24148 22520 24200
rect 23296 24148 23348 24200
rect 23572 24191 23624 24200
rect 23572 24157 23581 24191
rect 23581 24157 23615 24191
rect 23615 24157 23624 24191
rect 23572 24148 23624 24157
rect 23664 24191 23716 24200
rect 23664 24157 23673 24191
rect 23673 24157 23707 24191
rect 23707 24157 23716 24191
rect 23664 24148 23716 24157
rect 19892 24055 19944 24064
rect 19892 24021 19901 24055
rect 19901 24021 19935 24055
rect 19935 24021 19944 24055
rect 19892 24012 19944 24021
rect 20904 24012 20956 24064
rect 21180 24012 21232 24064
rect 25136 24012 25188 24064
rect 6884 23910 6936 23962
rect 6948 23910 7000 23962
rect 7012 23910 7064 23962
rect 7076 23910 7128 23962
rect 7140 23910 7192 23962
rect 12818 23910 12870 23962
rect 12882 23910 12934 23962
rect 12946 23910 12998 23962
rect 13010 23910 13062 23962
rect 13074 23910 13126 23962
rect 18752 23910 18804 23962
rect 18816 23910 18868 23962
rect 18880 23910 18932 23962
rect 18944 23910 18996 23962
rect 19008 23910 19060 23962
rect 24686 23910 24738 23962
rect 24750 23910 24802 23962
rect 24814 23910 24866 23962
rect 24878 23910 24930 23962
rect 24942 23910 24994 23962
rect 1860 23808 1912 23860
rect 3516 23851 3568 23860
rect 3516 23817 3525 23851
rect 3525 23817 3559 23851
rect 3559 23817 3568 23851
rect 3516 23808 3568 23817
rect 4068 23851 4120 23860
rect 4068 23817 4077 23851
rect 4077 23817 4111 23851
rect 4111 23817 4120 23851
rect 4068 23808 4120 23817
rect 4896 23808 4948 23860
rect 9772 23808 9824 23860
rect 9864 23808 9916 23860
rect 10324 23808 10376 23860
rect 3608 23740 3660 23792
rect 6092 23740 6144 23792
rect 6368 23740 6420 23792
rect 2780 23715 2832 23724
rect 2780 23681 2787 23715
rect 2787 23681 2821 23715
rect 2821 23681 2832 23715
rect 2780 23672 2832 23681
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 2228 23604 2280 23656
rect 5448 23672 5500 23724
rect 7288 23740 7340 23792
rect 7748 23740 7800 23792
rect 8116 23672 8168 23724
rect 8852 23783 8904 23792
rect 8852 23749 8861 23783
rect 8861 23749 8895 23783
rect 8895 23749 8904 23783
rect 8852 23740 8904 23749
rect 9220 23783 9272 23792
rect 9220 23749 9229 23783
rect 9229 23749 9263 23783
rect 9263 23749 9272 23783
rect 9220 23740 9272 23749
rect 10140 23740 10192 23792
rect 11796 23740 11848 23792
rect 12256 23740 12308 23792
rect 9588 23715 9640 23724
rect 9588 23681 9597 23715
rect 9597 23681 9631 23715
rect 9631 23681 9640 23715
rect 9588 23672 9640 23681
rect 9772 23672 9824 23724
rect 11612 23672 11664 23724
rect 13360 23808 13412 23860
rect 15660 23851 15712 23860
rect 15660 23817 15669 23851
rect 15669 23817 15703 23851
rect 15703 23817 15712 23851
rect 15660 23808 15712 23817
rect 15936 23808 15988 23860
rect 19248 23851 19300 23860
rect 19248 23817 19257 23851
rect 19257 23817 19291 23851
rect 19291 23817 19300 23851
rect 19248 23808 19300 23817
rect 13728 23672 13780 23724
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 14464 23672 14516 23724
rect 16580 23740 16632 23792
rect 19708 23808 19760 23860
rect 22560 23808 22612 23860
rect 19984 23740 20036 23792
rect 17684 23672 17736 23724
rect 8392 23604 8444 23656
rect 9680 23604 9732 23656
rect 11980 23604 12032 23656
rect 13176 23604 13228 23656
rect 13360 23604 13412 23656
rect 3516 23536 3568 23588
rect 10140 23579 10192 23588
rect 10140 23545 10149 23579
rect 10149 23545 10183 23579
rect 10183 23545 10192 23579
rect 10140 23536 10192 23545
rect 12624 23536 12676 23588
rect 6552 23468 6604 23520
rect 7932 23511 7984 23520
rect 7932 23477 7941 23511
rect 7941 23477 7975 23511
rect 7975 23477 7984 23511
rect 7932 23468 7984 23477
rect 8116 23468 8168 23520
rect 8392 23511 8444 23520
rect 8392 23477 8401 23511
rect 8401 23477 8435 23511
rect 8435 23477 8444 23511
rect 8392 23468 8444 23477
rect 11520 23468 11572 23520
rect 13820 23468 13872 23520
rect 14280 23468 14332 23520
rect 18420 23672 18472 23724
rect 23296 23808 23348 23860
rect 22652 23672 22704 23724
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 16028 23536 16080 23588
rect 16212 23536 16264 23588
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 19432 23468 19484 23520
rect 19616 23468 19668 23520
rect 23296 23511 23348 23520
rect 23296 23477 23305 23511
rect 23305 23477 23339 23511
rect 23339 23477 23348 23511
rect 23296 23468 23348 23477
rect 23572 23511 23624 23520
rect 23572 23477 23581 23511
rect 23581 23477 23615 23511
rect 23615 23477 23624 23511
rect 23572 23468 23624 23477
rect 24400 23511 24452 23520
rect 24400 23477 24409 23511
rect 24409 23477 24443 23511
rect 24443 23477 24452 23511
rect 24400 23468 24452 23477
rect 572 23400 624 23452
rect 3917 23366 3969 23418
rect 3981 23366 4033 23418
rect 4045 23366 4097 23418
rect 4109 23366 4161 23418
rect 4173 23366 4225 23418
rect 9851 23366 9903 23418
rect 9915 23366 9967 23418
rect 9979 23366 10031 23418
rect 10043 23366 10095 23418
rect 10107 23366 10159 23418
rect 15785 23366 15837 23418
rect 15849 23366 15901 23418
rect 15913 23366 15965 23418
rect 15977 23366 16029 23418
rect 16041 23366 16093 23418
rect 21719 23366 21771 23418
rect 21783 23366 21835 23418
rect 21847 23366 21899 23418
rect 21911 23366 21963 23418
rect 21975 23366 22027 23418
rect 572 23196 624 23248
rect 664 23196 716 23248
rect 2412 23307 2464 23316
rect 2412 23273 2421 23307
rect 2421 23273 2455 23307
rect 2455 23273 2464 23307
rect 2412 23264 2464 23273
rect 2872 23264 2924 23316
rect 3424 23264 3476 23316
rect 5724 23264 5776 23316
rect 19892 23264 19944 23316
rect 23940 23264 23992 23316
rect 24400 23264 24452 23316
rect 25412 23264 25464 23316
rect 3516 23196 3568 23248
rect 3976 23196 4028 23248
rect 5632 23196 5684 23248
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2872 23128 2924 23180
rect 4620 23128 4672 23180
rect 1308 22992 1360 23044
rect 2872 22992 2924 23044
rect 5264 23060 5316 23112
rect 5448 23060 5500 23112
rect 7472 23060 7524 23112
rect 7564 23060 7616 23112
rect 7932 23171 7984 23180
rect 7932 23137 7941 23171
rect 7941 23137 7975 23171
rect 7975 23137 7984 23171
rect 7932 23128 7984 23137
rect 11060 23128 11112 23180
rect 12164 23128 12216 23180
rect 13268 23128 13320 23180
rect 13820 23128 13872 23180
rect 8392 23060 8444 23112
rect 10692 23060 10744 23112
rect 11244 23060 11296 23112
rect 11796 23060 11848 23112
rect 14372 23103 14424 23112
rect 14372 23069 14379 23103
rect 14379 23069 14413 23103
rect 14413 23069 14424 23103
rect 14372 23060 14424 23069
rect 14832 23060 14884 23112
rect 18420 23060 18472 23112
rect 19616 23103 19668 23112
rect 19616 23069 19625 23103
rect 19625 23069 19659 23103
rect 19659 23069 19668 23103
rect 19616 23060 19668 23069
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 1676 22924 1728 22976
rect 8116 23035 8168 23044
rect 8116 23001 8125 23035
rect 8125 23001 8159 23035
rect 8159 23001 8168 23035
rect 8116 22992 8168 23001
rect 10140 23035 10192 23044
rect 10140 23001 10149 23035
rect 10149 23001 10183 23035
rect 10183 23001 10192 23035
rect 10140 22992 10192 23001
rect 14280 22992 14332 23044
rect 18052 22992 18104 23044
rect 19340 22992 19392 23044
rect 20536 22992 20588 23044
rect 21732 23060 21784 23112
rect 22376 23103 22428 23112
rect 22376 23069 22385 23103
rect 22385 23069 22419 23103
rect 22419 23069 22428 23103
rect 22376 23060 22428 23069
rect 22652 23103 22704 23112
rect 22652 23069 22686 23103
rect 22686 23069 22704 23103
rect 22652 23060 22704 23069
rect 23756 23060 23808 23112
rect 6644 22924 6696 22976
rect 7472 22924 7524 22976
rect 9404 22924 9456 22976
rect 10416 22924 10468 22976
rect 11612 22924 11664 22976
rect 14464 22924 14516 22976
rect 15292 22924 15344 22976
rect 21272 22924 21324 22976
rect 22100 22924 22152 22976
rect 22192 22967 22244 22976
rect 22192 22933 22201 22967
rect 22201 22933 22235 22967
rect 22235 22933 22244 22967
rect 22192 22924 22244 22933
rect 23480 22924 23532 22976
rect 24032 22924 24084 22976
rect 25136 22924 25188 22976
rect 6884 22822 6936 22874
rect 6948 22822 7000 22874
rect 7012 22822 7064 22874
rect 7076 22822 7128 22874
rect 7140 22822 7192 22874
rect 12818 22822 12870 22874
rect 12882 22822 12934 22874
rect 12946 22822 12998 22874
rect 13010 22822 13062 22874
rect 13074 22822 13126 22874
rect 18752 22822 18804 22874
rect 18816 22822 18868 22874
rect 18880 22822 18932 22874
rect 18944 22822 18996 22874
rect 19008 22822 19060 22874
rect 24686 22822 24738 22874
rect 24750 22822 24802 22874
rect 24814 22822 24866 22874
rect 24878 22822 24930 22874
rect 24942 22822 24994 22874
rect 204 22720 256 22772
rect 3056 22720 3108 22772
rect 3148 22720 3200 22772
rect 3240 22720 3292 22772
rect 4344 22720 4396 22772
rect 4436 22720 4488 22772
rect 5632 22720 5684 22772
rect 6552 22720 6604 22772
rect 7564 22720 7616 22772
rect 9220 22720 9272 22772
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 14004 22720 14056 22772
rect 16028 22720 16080 22772
rect 16856 22720 16908 22772
rect 19524 22720 19576 22772
rect 20076 22720 20128 22772
rect 20536 22720 20588 22772
rect 21732 22720 21784 22772
rect 1952 22652 2004 22704
rect 2228 22584 2280 22636
rect 4252 22652 4304 22704
rect 4620 22652 4672 22704
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 2412 22423 2464 22432
rect 2412 22389 2421 22423
rect 2421 22389 2455 22423
rect 2455 22389 2464 22423
rect 2412 22380 2464 22389
rect 2780 22380 2832 22432
rect 4896 22584 4948 22636
rect 6184 22584 6236 22636
rect 12072 22652 12124 22704
rect 10324 22627 10376 22636
rect 10324 22593 10331 22627
rect 10331 22593 10365 22627
rect 10365 22593 10376 22627
rect 10324 22584 10376 22593
rect 8300 22516 8352 22568
rect 7288 22448 7340 22500
rect 8116 22448 8168 22500
rect 4620 22380 4672 22432
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 6736 22380 6788 22432
rect 10968 22516 11020 22568
rect 11060 22516 11112 22568
rect 11336 22516 11388 22568
rect 11704 22516 11756 22568
rect 12164 22516 12216 22568
rect 12348 22516 12400 22568
rect 15476 22516 15528 22568
rect 14188 22448 14240 22500
rect 14372 22448 14424 22500
rect 11612 22380 11664 22432
rect 14832 22423 14884 22432
rect 14832 22389 14841 22423
rect 14841 22389 14875 22423
rect 14875 22389 14884 22423
rect 14832 22380 14884 22389
rect 15660 22516 15712 22568
rect 16580 22584 16632 22636
rect 16856 22627 16908 22636
rect 16856 22593 16865 22627
rect 16865 22593 16899 22627
rect 16899 22593 16908 22627
rect 16856 22584 16908 22593
rect 17776 22584 17828 22636
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 21732 22584 21784 22636
rect 22008 22584 22060 22636
rect 22284 22652 22336 22704
rect 23204 22720 23256 22772
rect 23848 22652 23900 22704
rect 24492 22652 24544 22704
rect 22560 22584 22612 22636
rect 23480 22627 23532 22636
rect 23480 22593 23487 22627
rect 23487 22593 23521 22627
rect 23521 22593 23532 22627
rect 23480 22584 23532 22593
rect 17868 22559 17920 22568
rect 17868 22525 17877 22559
rect 17877 22525 17911 22559
rect 17911 22525 17920 22559
rect 17868 22516 17920 22525
rect 17316 22491 17368 22500
rect 17316 22457 17325 22491
rect 17325 22457 17359 22491
rect 17359 22457 17368 22491
rect 17316 22448 17368 22457
rect 16672 22380 16724 22432
rect 17224 22380 17276 22432
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 22284 22380 22336 22432
rect 22836 22423 22888 22432
rect 22836 22389 22845 22423
rect 22845 22389 22879 22423
rect 22879 22389 22888 22423
rect 22836 22380 22888 22389
rect 3917 22278 3969 22330
rect 3981 22278 4033 22330
rect 4045 22278 4097 22330
rect 4109 22278 4161 22330
rect 4173 22278 4225 22330
rect 9851 22278 9903 22330
rect 9915 22278 9967 22330
rect 9979 22278 10031 22330
rect 10043 22278 10095 22330
rect 10107 22278 10159 22330
rect 15785 22278 15837 22330
rect 15849 22278 15901 22330
rect 15913 22278 15965 22330
rect 15977 22278 16029 22330
rect 16041 22278 16093 22330
rect 21719 22278 21771 22330
rect 21783 22278 21835 22330
rect 21847 22278 21899 22330
rect 21911 22278 21963 22330
rect 21975 22278 22027 22330
rect 3056 22219 3108 22228
rect 3056 22185 3065 22219
rect 3065 22185 3099 22219
rect 3099 22185 3108 22219
rect 3056 22176 3108 22185
rect 3240 22176 3292 22228
rect 3516 22176 3568 22228
rect 3608 22176 3660 22228
rect 3792 22176 3844 22228
rect 9036 22176 9088 22228
rect 9128 22176 9180 22228
rect 9496 22176 9548 22228
rect 9956 22176 10008 22228
rect 10876 22176 10928 22228
rect 2320 22040 2372 22092
rect 2412 21972 2464 22024
rect 3608 21972 3660 22024
rect 1768 21947 1820 21956
rect 1768 21913 1777 21947
rect 1777 21913 1811 21947
rect 1811 21913 1820 21947
rect 1768 21904 1820 21913
rect 2044 21947 2096 21956
rect 2044 21913 2053 21947
rect 2053 21913 2087 21947
rect 2087 21913 2096 21947
rect 2044 21904 2096 21913
rect 6184 22108 6236 22160
rect 6552 22151 6604 22160
rect 6552 22117 6561 22151
rect 6561 22117 6595 22151
rect 6595 22117 6604 22151
rect 6552 22108 6604 22117
rect 7656 22108 7708 22160
rect 5172 22040 5224 22092
rect 19156 22176 19208 22228
rect 17316 22151 17368 22160
rect 17316 22117 17325 22151
rect 17325 22117 17359 22151
rect 17359 22117 17368 22151
rect 17316 22108 17368 22117
rect 18512 22108 18564 22160
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 14832 22040 14884 22092
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 5264 21972 5316 22024
rect 1216 21836 1268 21888
rect 3976 21904 4028 21956
rect 5172 21904 5224 21956
rect 5632 21904 5684 21956
rect 6552 21972 6604 22024
rect 7656 21972 7708 22024
rect 8024 21972 8076 22024
rect 9588 21972 9640 22024
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 10416 21972 10468 22024
rect 13360 21972 13412 22024
rect 3056 21836 3108 21888
rect 4068 21836 4120 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 6000 21836 6052 21888
rect 7380 21836 7432 21888
rect 10600 21836 10652 21888
rect 11244 21836 11296 21888
rect 11888 21947 11940 21956
rect 11888 21913 11897 21947
rect 11897 21913 11931 21947
rect 11931 21913 11940 21947
rect 11888 21904 11940 21913
rect 11980 21947 12032 21956
rect 11980 21913 11989 21947
rect 11989 21913 12023 21947
rect 12023 21913 12032 21947
rect 11980 21904 12032 21913
rect 12164 21904 12216 21956
rect 15108 22015 15160 22024
rect 15108 21981 15142 22015
rect 15142 21981 15160 22015
rect 15108 21972 15160 21981
rect 16120 21972 16172 22024
rect 16580 22015 16632 22024
rect 16580 21981 16587 22015
rect 16587 21981 16621 22015
rect 16621 21981 16632 22015
rect 16580 21972 16632 21981
rect 14832 21836 14884 21888
rect 17224 21904 17276 21956
rect 17500 21904 17552 21956
rect 20628 22176 20680 22228
rect 20720 22176 20772 22228
rect 22008 22176 22060 22228
rect 22192 22176 22244 22228
rect 21456 22108 21508 22160
rect 22836 22176 22888 22228
rect 23572 22176 23624 22228
rect 20260 22040 20312 22092
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 19800 21972 19852 22024
rect 20076 21972 20128 22024
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 19892 21904 19944 21956
rect 20352 21904 20404 21956
rect 20720 21904 20772 21956
rect 22468 22108 22520 22160
rect 22284 22083 22336 22092
rect 22284 22049 22293 22083
rect 22293 22049 22327 22083
rect 22327 22049 22336 22083
rect 22284 22040 22336 22049
rect 23388 22083 23440 22092
rect 23388 22049 23397 22083
rect 23397 22049 23431 22083
rect 23431 22049 23440 22083
rect 23388 22040 23440 22049
rect 22100 21972 22152 22024
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 24032 22040 24084 22092
rect 23756 21972 23808 22024
rect 24216 22015 24268 22024
rect 24216 21981 24225 22015
rect 24225 21981 24259 22015
rect 24259 21981 24268 22015
rect 24216 21972 24268 21981
rect 23480 21904 23532 21956
rect 17776 21836 17828 21888
rect 18604 21836 18656 21888
rect 20904 21836 20956 21888
rect 20996 21879 21048 21888
rect 20996 21845 21005 21879
rect 21005 21845 21039 21879
rect 21039 21845 21048 21879
rect 20996 21836 21048 21845
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23388 21879 23440 21888
rect 23388 21845 23397 21879
rect 23397 21845 23431 21879
rect 23431 21845 23440 21879
rect 23388 21836 23440 21845
rect 25136 21904 25188 21956
rect 6884 21734 6936 21786
rect 6948 21734 7000 21786
rect 7012 21734 7064 21786
rect 7076 21734 7128 21786
rect 7140 21734 7192 21786
rect 12818 21734 12870 21786
rect 12882 21734 12934 21786
rect 12946 21734 12998 21786
rect 13010 21734 13062 21786
rect 13074 21734 13126 21786
rect 18752 21734 18804 21786
rect 18816 21734 18868 21786
rect 18880 21734 18932 21786
rect 18944 21734 18996 21786
rect 19008 21734 19060 21786
rect 24686 21734 24738 21786
rect 24750 21734 24802 21786
rect 24814 21734 24866 21786
rect 24878 21734 24930 21786
rect 24942 21734 24994 21786
rect 1308 21632 1360 21684
rect 1676 21569 1728 21616
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 1676 21564 1701 21569
rect 1701 21564 1728 21569
rect 2320 21632 2372 21684
rect 2596 21632 2648 21684
rect 4068 21632 4120 21684
rect 4620 21632 4672 21684
rect 5080 21632 5132 21684
rect 6092 21632 6144 21684
rect 6368 21564 6420 21616
rect 6644 21564 6696 21616
rect 7380 21564 7432 21616
rect 7472 21564 7524 21616
rect 8944 21632 8996 21684
rect 9128 21632 9180 21684
rect 9680 21632 9732 21684
rect 10692 21632 10744 21684
rect 10968 21632 11020 21684
rect 11980 21632 12032 21684
rect 14740 21632 14792 21684
rect 8392 21564 8444 21616
rect 11060 21564 11112 21616
rect 12164 21564 12216 21616
rect 20260 21632 20312 21684
rect 20812 21632 20864 21684
rect 7196 21496 7248 21548
rect 8760 21539 8812 21548
rect 8760 21505 8769 21539
rect 8769 21505 8803 21539
rect 8803 21505 8812 21539
rect 8760 21496 8812 21505
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 8944 21496 8996 21548
rect 15200 21564 15252 21616
rect 13544 21539 13596 21548
rect 13544 21505 13551 21539
rect 13551 21505 13585 21539
rect 13585 21505 13596 21539
rect 16304 21564 16356 21616
rect 16764 21564 16816 21616
rect 18604 21564 18656 21616
rect 13544 21496 13596 21505
rect 6736 21428 6788 21480
rect 8484 21428 8536 21480
rect 9588 21428 9640 21480
rect 9864 21428 9916 21480
rect 10600 21428 10652 21480
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 1308 21292 1360 21344
rect 4620 21360 4672 21412
rect 5632 21360 5684 21412
rect 5908 21360 5960 21412
rect 7840 21403 7892 21412
rect 7840 21369 7849 21403
rect 7849 21369 7883 21403
rect 7883 21369 7892 21403
rect 7840 21360 7892 21369
rect 10048 21360 10100 21412
rect 10416 21360 10468 21412
rect 4804 21292 4856 21344
rect 6000 21292 6052 21344
rect 10324 21292 10376 21344
rect 10692 21292 10744 21344
rect 14372 21292 14424 21344
rect 16120 21428 16172 21480
rect 16488 21428 16540 21480
rect 17592 21539 17644 21548
rect 17592 21505 17601 21539
rect 17601 21505 17635 21539
rect 17635 21505 17644 21539
rect 17592 21496 17644 21505
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 16764 21428 16816 21480
rect 17040 21428 17092 21480
rect 17684 21471 17736 21480
rect 17684 21437 17718 21471
rect 17718 21437 17736 21471
rect 17684 21428 17736 21437
rect 18052 21428 18104 21480
rect 19524 21496 19576 21548
rect 19800 21539 19852 21548
rect 19800 21505 19809 21539
rect 19809 21505 19843 21539
rect 19843 21505 19852 21539
rect 19800 21496 19852 21505
rect 20996 21632 21048 21684
rect 21548 21632 21600 21684
rect 22284 21632 22336 21684
rect 24492 21632 24544 21684
rect 21456 21496 21508 21548
rect 23480 21496 23532 21548
rect 23112 21428 23164 21480
rect 23664 21539 23716 21548
rect 23664 21505 23673 21539
rect 23673 21505 23707 21539
rect 23707 21505 23716 21539
rect 23664 21496 23716 21505
rect 15016 21335 15068 21344
rect 15016 21301 15025 21335
rect 15025 21301 15059 21335
rect 15059 21301 15068 21335
rect 15016 21292 15068 21301
rect 15108 21292 15160 21344
rect 16120 21335 16172 21344
rect 16120 21301 16129 21335
rect 16129 21301 16163 21335
rect 16163 21301 16172 21335
rect 16120 21292 16172 21301
rect 17132 21360 17184 21412
rect 17224 21360 17276 21412
rect 19340 21360 19392 21412
rect 23664 21360 23716 21412
rect 17592 21292 17644 21344
rect 18788 21292 18840 21344
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 21364 21335 21416 21344
rect 21364 21301 21373 21335
rect 21373 21301 21407 21335
rect 21407 21301 21416 21335
rect 21364 21292 21416 21301
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 23848 21335 23900 21344
rect 23848 21301 23857 21335
rect 23857 21301 23891 21335
rect 23891 21301 23900 21335
rect 23848 21292 23900 21301
rect 3917 21190 3969 21242
rect 3981 21190 4033 21242
rect 4045 21190 4097 21242
rect 4109 21190 4161 21242
rect 4173 21190 4225 21242
rect 9851 21190 9903 21242
rect 9915 21190 9967 21242
rect 9979 21190 10031 21242
rect 10043 21190 10095 21242
rect 10107 21190 10159 21242
rect 15785 21190 15837 21242
rect 15849 21190 15901 21242
rect 15913 21190 15965 21242
rect 15977 21190 16029 21242
rect 16041 21190 16093 21242
rect 21719 21190 21771 21242
rect 21783 21190 21835 21242
rect 21847 21190 21899 21242
rect 21911 21190 21963 21242
rect 21975 21190 22027 21242
rect 1400 21088 1452 21140
rect 8392 21088 8444 21140
rect 8484 21131 8536 21140
rect 8484 21097 8493 21131
rect 8493 21097 8527 21131
rect 8527 21097 8536 21131
rect 8484 21088 8536 21097
rect 8852 21088 8904 21140
rect 1216 20952 1268 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 2136 20884 2188 20936
rect 1308 20816 1360 20868
rect 2872 21020 2924 21072
rect 4712 21020 4764 21072
rect 8208 21020 8260 21072
rect 5908 20952 5960 21004
rect 8484 20952 8536 21004
rect 8668 20952 8720 21004
rect 8852 20952 8904 21004
rect 2780 20884 2832 20936
rect 4160 20884 4212 20936
rect 4436 20884 4488 20936
rect 5264 20884 5316 20936
rect 7840 20884 7892 20936
rect 8300 20816 8352 20868
rect 9588 20884 9640 20936
rect 14832 21088 14884 21140
rect 15016 21088 15068 21140
rect 15384 21088 15436 21140
rect 17868 21088 17920 21140
rect 19616 21088 19668 21140
rect 21364 21088 21416 21140
rect 10324 20995 10376 21004
rect 10324 20961 10333 20995
rect 10333 20961 10367 20995
rect 10367 20961 10376 20995
rect 10324 20952 10376 20961
rect 13360 20952 13412 21004
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 16120 20952 16172 21004
rect 16304 20952 16356 21004
rect 16488 20952 16540 21004
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10652 20927
rect 10600 20884 10652 20893
rect 11704 20884 11756 20936
rect 11796 20884 11848 20936
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 1952 20748 2004 20800
rect 2964 20748 3016 20800
rect 4068 20748 4120 20800
rect 5080 20748 5132 20800
rect 7656 20748 7708 20800
rect 8116 20748 8168 20800
rect 9404 20816 9456 20868
rect 12348 20884 12400 20936
rect 13268 20884 13320 20936
rect 15752 20927 15804 20936
rect 18788 20952 18840 21004
rect 15752 20893 15786 20927
rect 15786 20893 15804 20927
rect 15752 20884 15804 20893
rect 16672 20816 16724 20868
rect 19340 20952 19392 21004
rect 19156 20884 19208 20936
rect 20720 21063 20772 21072
rect 20720 21029 20729 21063
rect 20729 21029 20763 21063
rect 20763 21029 20772 21063
rect 20720 21020 20772 21029
rect 20260 20952 20312 21004
rect 24216 21088 24268 21140
rect 22376 20952 22428 21004
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 22100 20884 22152 20936
rect 24032 20927 24084 20936
rect 24032 20893 24041 20927
rect 24041 20893 24075 20927
rect 24075 20893 24084 20927
rect 24032 20884 24084 20893
rect 8668 20748 8720 20800
rect 10968 20748 11020 20800
rect 12716 20748 12768 20800
rect 14464 20748 14516 20800
rect 15752 20748 15804 20800
rect 16580 20791 16632 20800
rect 16580 20757 16589 20791
rect 16589 20757 16623 20791
rect 16623 20757 16632 20791
rect 16580 20748 16632 20757
rect 22652 20816 22704 20868
rect 19708 20748 19760 20800
rect 23296 20748 23348 20800
rect 24216 20748 24268 20800
rect 6884 20646 6936 20698
rect 6948 20646 7000 20698
rect 7012 20646 7064 20698
rect 7076 20646 7128 20698
rect 7140 20646 7192 20698
rect 12818 20646 12870 20698
rect 12882 20646 12934 20698
rect 12946 20646 12998 20698
rect 13010 20646 13062 20698
rect 13074 20646 13126 20698
rect 18752 20646 18804 20698
rect 18816 20646 18868 20698
rect 18880 20646 18932 20698
rect 18944 20646 18996 20698
rect 19008 20646 19060 20698
rect 24686 20646 24738 20698
rect 24750 20646 24802 20698
rect 24814 20646 24866 20698
rect 24878 20646 24930 20698
rect 24942 20646 24994 20698
rect 3792 20544 3844 20596
rect 7840 20544 7892 20596
rect 8852 20544 8904 20596
rect 9220 20544 9272 20596
rect 2596 20408 2648 20460
rect 3884 20451 3936 20460
rect 3884 20417 3918 20451
rect 3918 20417 3936 20451
rect 3884 20408 3936 20417
rect 4068 20451 4120 20460
rect 4068 20417 4077 20451
rect 4077 20417 4111 20451
rect 4111 20417 4120 20451
rect 4068 20408 4120 20417
rect 5264 20476 5316 20528
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 2964 20340 3016 20392
rect 4252 20340 4304 20392
rect 6552 20408 6604 20460
rect 10416 20544 10468 20596
rect 10508 20476 10560 20528
rect 11244 20544 11296 20596
rect 11336 20476 11388 20528
rect 10600 20408 10652 20460
rect 11428 20408 11480 20460
rect 8668 20340 8720 20392
rect 10968 20340 11020 20392
rect 1860 20204 1912 20256
rect 3516 20315 3568 20324
rect 3516 20281 3525 20315
rect 3525 20281 3559 20315
rect 3559 20281 3568 20315
rect 3516 20272 3568 20281
rect 11704 20408 11756 20460
rect 13268 20544 13320 20596
rect 15384 20587 15436 20596
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 15476 20544 15528 20596
rect 16212 20544 16264 20596
rect 18052 20544 18104 20596
rect 19156 20544 19208 20596
rect 22100 20544 22152 20596
rect 23572 20544 23624 20596
rect 14740 20476 14792 20528
rect 19616 20476 19668 20528
rect 13360 20451 13412 20460
rect 13360 20417 13394 20451
rect 13394 20417 13412 20451
rect 13360 20408 13412 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 14372 20451 14424 20460
rect 14372 20417 14381 20451
rect 14381 20417 14415 20451
rect 14415 20417 14424 20451
rect 14372 20408 14424 20417
rect 14648 20451 14700 20460
rect 14648 20417 14657 20451
rect 14657 20417 14700 20451
rect 14648 20408 14700 20417
rect 16304 20408 16356 20460
rect 17960 20408 18012 20460
rect 18512 20408 18564 20460
rect 19156 20408 19208 20460
rect 22100 20408 22152 20460
rect 22560 20408 22612 20460
rect 22836 20476 22888 20528
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 12624 20340 12676 20392
rect 12716 20340 12768 20392
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 4712 20247 4764 20256
rect 4712 20213 4721 20247
rect 4721 20213 4755 20247
rect 4755 20213 4764 20247
rect 4712 20204 4764 20213
rect 5816 20247 5868 20256
rect 5816 20213 5825 20247
rect 5825 20213 5859 20247
rect 5859 20213 5868 20247
rect 5816 20204 5868 20213
rect 6644 20204 6696 20256
rect 9404 20204 9456 20256
rect 11244 20247 11296 20256
rect 11244 20213 11253 20247
rect 11253 20213 11287 20247
rect 11287 20213 11296 20247
rect 11244 20204 11296 20213
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 15384 20340 15436 20392
rect 15752 20340 15804 20392
rect 23480 20340 23532 20392
rect 16948 20272 17000 20324
rect 17684 20272 17736 20324
rect 22652 20272 22704 20324
rect 16120 20204 16172 20256
rect 16672 20204 16724 20256
rect 24032 20272 24084 20324
rect 24216 20204 24268 20256
rect 3917 20102 3969 20154
rect 3981 20102 4033 20154
rect 4045 20102 4097 20154
rect 4109 20102 4161 20154
rect 4173 20102 4225 20154
rect 9851 20102 9903 20154
rect 9915 20102 9967 20154
rect 9979 20102 10031 20154
rect 10043 20102 10095 20154
rect 10107 20102 10159 20154
rect 15785 20102 15837 20154
rect 15849 20102 15901 20154
rect 15913 20102 15965 20154
rect 15977 20102 16029 20154
rect 16041 20102 16093 20154
rect 21719 20102 21771 20154
rect 21783 20102 21835 20154
rect 21847 20102 21899 20154
rect 21911 20102 21963 20154
rect 21975 20102 22027 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 2228 19864 2280 19916
rect 2780 20000 2832 20052
rect 3516 20000 3568 20052
rect 5172 20000 5224 20052
rect 10600 20000 10652 20052
rect 11980 20000 12032 20052
rect 5816 19864 5868 19916
rect 6552 19864 6604 19916
rect 7656 19864 7708 19916
rect 13360 20000 13412 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 14004 20000 14056 20052
rect 16304 20000 16356 20052
rect 16580 20000 16632 20052
rect 17776 19932 17828 19984
rect 14188 19864 14240 19916
rect 16304 19907 16356 19916
rect 16304 19873 16313 19907
rect 16313 19873 16347 19907
rect 16347 19873 16356 19907
rect 16304 19864 16356 19873
rect 16396 19864 16448 19916
rect 756 19796 808 19848
rect 2596 19839 2648 19848
rect 2596 19805 2603 19839
rect 2603 19805 2637 19839
rect 2637 19805 2648 19839
rect 2596 19796 2648 19805
rect 1308 19728 1360 19780
rect 4436 19728 4488 19780
rect 5356 19796 5408 19848
rect 5540 19771 5592 19780
rect 5540 19737 5549 19771
rect 5549 19737 5583 19771
rect 5583 19737 5592 19771
rect 5540 19728 5592 19737
rect 5908 19839 5960 19848
rect 5908 19805 5917 19839
rect 5917 19805 5951 19839
rect 5951 19805 5960 19839
rect 5908 19796 5960 19805
rect 8300 19796 8352 19848
rect 8392 19796 8444 19848
rect 10048 19796 10100 19848
rect 10324 19796 10376 19848
rect 10876 19796 10928 19848
rect 11244 19796 11296 19848
rect 11612 19796 11664 19848
rect 12716 19796 12768 19848
rect 13268 19796 13320 19848
rect 13452 19796 13504 19848
rect 14648 19796 14700 19848
rect 17040 19864 17092 19916
rect 7564 19728 7616 19780
rect 8944 19728 8996 19780
rect 15108 19728 15160 19780
rect 16856 19839 16908 19848
rect 16856 19805 16865 19839
rect 16865 19805 16899 19839
rect 16899 19805 16908 19839
rect 16856 19796 16908 19805
rect 22100 20043 22152 20052
rect 22100 20009 22109 20043
rect 22109 20009 22143 20043
rect 22143 20009 22152 20043
rect 22100 20000 22152 20009
rect 22560 20000 22612 20052
rect 24032 20000 24084 20052
rect 19248 19839 19300 19848
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 21272 19796 21324 19848
rect 21548 19796 21600 19848
rect 23664 19839 23716 19848
rect 23664 19805 23673 19839
rect 23673 19805 23707 19839
rect 23707 19805 23716 19839
rect 23664 19796 23716 19805
rect 6736 19660 6788 19712
rect 6828 19660 6880 19712
rect 11704 19660 11756 19712
rect 11980 19660 12032 19712
rect 14280 19660 14332 19712
rect 16580 19660 16632 19712
rect 17316 19660 17368 19712
rect 17960 19660 18012 19712
rect 18604 19660 18656 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 20812 19660 20864 19712
rect 23848 19728 23900 19780
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 6884 19558 6936 19610
rect 6948 19558 7000 19610
rect 7012 19558 7064 19610
rect 7076 19558 7128 19610
rect 7140 19558 7192 19610
rect 12818 19558 12870 19610
rect 12882 19558 12934 19610
rect 12946 19558 12998 19610
rect 13010 19558 13062 19610
rect 13074 19558 13126 19610
rect 18752 19558 18804 19610
rect 18816 19558 18868 19610
rect 18880 19558 18932 19610
rect 18944 19558 18996 19610
rect 19008 19558 19060 19610
rect 24686 19558 24738 19610
rect 24750 19558 24802 19610
rect 24814 19558 24866 19610
rect 24878 19558 24930 19610
rect 24942 19558 24994 19610
rect 1584 19499 1636 19508
rect 1584 19465 1593 19499
rect 1593 19465 1627 19499
rect 1627 19465 1636 19499
rect 1584 19456 1636 19465
rect 2044 19456 2096 19508
rect 4620 19456 4672 19508
rect 4712 19456 4764 19508
rect 5264 19456 5316 19508
rect 5540 19456 5592 19508
rect 6644 19456 6696 19508
rect 7472 19456 7524 19508
rect 7932 19456 7984 19508
rect 848 19320 900 19372
rect 2596 19320 2648 19372
rect 3332 19363 3384 19372
rect 3332 19329 3341 19363
rect 3341 19329 3375 19363
rect 3375 19329 3384 19363
rect 3332 19320 3384 19329
rect 8300 19456 8352 19508
rect 9128 19456 9180 19508
rect 14188 19456 14240 19508
rect 14280 19456 14332 19508
rect 8208 19431 8260 19440
rect 8208 19397 8217 19431
rect 8217 19397 8251 19431
rect 8251 19397 8260 19431
rect 8208 19388 8260 19397
rect 8576 19388 8628 19440
rect 9772 19388 9824 19440
rect 10048 19388 10100 19440
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 8300 19320 8352 19372
rect 8392 19320 8444 19372
rect 10324 19320 10376 19372
rect 11704 19320 11756 19372
rect 12256 19320 12308 19372
rect 14004 19388 14056 19440
rect 16120 19388 16172 19440
rect 16580 19388 16632 19440
rect 16856 19456 16908 19508
rect 13728 19363 13780 19372
rect 13728 19329 13735 19363
rect 13735 19329 13769 19363
rect 13769 19329 13780 19363
rect 13728 19320 13780 19329
rect 14464 19320 14516 19372
rect 16396 19320 16448 19372
rect 17316 19388 17368 19440
rect 19524 19388 19576 19440
rect 19616 19388 19668 19440
rect 19800 19320 19852 19372
rect 20812 19499 20864 19508
rect 20812 19465 20821 19499
rect 20821 19465 20855 19499
rect 20855 19465 20864 19499
rect 20812 19456 20864 19465
rect 22836 19456 22888 19508
rect 23204 19456 23256 19508
rect 23296 19456 23348 19508
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 21272 19320 21324 19372
rect 1676 19295 1728 19304
rect 1676 19261 1685 19295
rect 1685 19261 1719 19295
rect 1719 19261 1728 19295
rect 1676 19252 1728 19261
rect 4252 19252 4304 19304
rect 204 19116 256 19168
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 4252 19116 4304 19168
rect 7656 19252 7708 19304
rect 11244 19252 11296 19304
rect 22652 19363 22704 19372
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 23112 19320 23164 19372
rect 23940 19388 23992 19440
rect 24124 19431 24176 19440
rect 24124 19397 24133 19431
rect 24133 19397 24167 19431
rect 24167 19397 24176 19431
rect 24124 19388 24176 19397
rect 5356 19116 5408 19168
rect 9680 19116 9732 19168
rect 9956 19116 10008 19168
rect 10324 19116 10376 19168
rect 12716 19116 12768 19168
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14464 19116 14516 19125
rect 14740 19116 14792 19168
rect 15568 19116 15620 19168
rect 20536 19184 20588 19236
rect 21180 19184 21232 19236
rect 23112 19184 23164 19236
rect 25136 19252 25188 19304
rect 20260 19116 20312 19168
rect 23848 19159 23900 19168
rect 23848 19125 23857 19159
rect 23857 19125 23891 19159
rect 23891 19125 23900 19159
rect 23848 19116 23900 19125
rect 3917 19014 3969 19066
rect 3981 19014 4033 19066
rect 4045 19014 4097 19066
rect 4109 19014 4161 19066
rect 4173 19014 4225 19066
rect 9851 19014 9903 19066
rect 9915 19014 9967 19066
rect 9979 19014 10031 19066
rect 10043 19014 10095 19066
rect 10107 19014 10159 19066
rect 15785 19014 15837 19066
rect 15849 19014 15901 19066
rect 15913 19014 15965 19066
rect 15977 19014 16029 19066
rect 16041 19014 16093 19066
rect 21719 19014 21771 19066
rect 21783 19014 21835 19066
rect 21847 19014 21899 19066
rect 21911 19014 21963 19066
rect 21975 19014 22027 19066
rect 1400 18912 1452 18964
rect 4620 18912 4672 18964
rect 7472 18912 7524 18964
rect 10508 18912 10560 18964
rect 13820 18912 13872 18964
rect 16120 18912 16172 18964
rect 16304 18912 16356 18964
rect 18604 18912 18656 18964
rect 20260 18912 20312 18964
rect 21088 18912 21140 18964
rect 4712 18844 4764 18896
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 6644 18776 6696 18828
rect 8944 18776 8996 18828
rect 2320 18708 2372 18760
rect 1308 18640 1360 18692
rect 4068 18741 4120 18760
rect 4068 18708 4093 18741
rect 4093 18708 4120 18741
rect 5816 18708 5868 18760
rect 8024 18708 8076 18760
rect 12072 18776 12124 18828
rect 14188 18776 14240 18828
rect 14464 18844 14516 18896
rect 15016 18819 15068 18828
rect 15016 18785 15025 18819
rect 15025 18785 15059 18819
rect 15059 18785 15068 18819
rect 15016 18776 15068 18785
rect 15108 18819 15160 18828
rect 15108 18785 15142 18819
rect 15142 18785 15160 18819
rect 15108 18776 15160 18785
rect 8300 18640 8352 18692
rect 9496 18683 9548 18692
rect 9496 18649 9505 18683
rect 9505 18649 9539 18683
rect 9539 18649 9548 18683
rect 9496 18640 9548 18649
rect 9864 18683 9916 18692
rect 9864 18649 9873 18683
rect 9873 18649 9907 18683
rect 9907 18649 9916 18683
rect 9864 18640 9916 18649
rect 10048 18640 10100 18692
rect 10876 18640 10928 18692
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 11612 18708 11664 18760
rect 14280 18751 14332 18760
rect 14280 18717 14289 18751
rect 14289 18717 14323 18751
rect 14323 18717 14332 18751
rect 14280 18708 14332 18717
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 17132 18708 17184 18760
rect 16304 18687 16329 18692
rect 16329 18687 16356 18692
rect 940 18572 992 18624
rect 1216 18572 1268 18624
rect 2872 18572 2924 18624
rect 3884 18572 3936 18624
rect 3976 18572 4028 18624
rect 8668 18572 8720 18624
rect 9588 18572 9640 18624
rect 10600 18572 10652 18624
rect 12072 18572 12124 18624
rect 12256 18615 12308 18624
rect 12256 18581 12265 18615
rect 12265 18581 12299 18615
rect 12299 18581 12308 18615
rect 12256 18572 12308 18581
rect 16304 18640 16356 18687
rect 20628 18708 20680 18760
rect 23480 18844 23532 18896
rect 25136 18844 25188 18896
rect 23664 18776 23716 18828
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 14832 18572 14884 18624
rect 15936 18615 15988 18624
rect 15936 18581 15945 18615
rect 15945 18581 15979 18615
rect 15979 18581 15988 18615
rect 15936 18572 15988 18581
rect 18328 18572 18380 18624
rect 23388 18751 23440 18760
rect 23388 18717 23397 18751
rect 23397 18717 23431 18751
rect 23431 18717 23440 18751
rect 23388 18708 23440 18717
rect 24308 18776 24360 18828
rect 25504 18708 25556 18760
rect 20904 18572 20956 18624
rect 23020 18615 23072 18624
rect 23020 18581 23029 18615
rect 23029 18581 23063 18615
rect 23063 18581 23072 18615
rect 23020 18572 23072 18581
rect 23112 18572 23164 18624
rect 6884 18470 6936 18522
rect 6948 18470 7000 18522
rect 7012 18470 7064 18522
rect 7076 18470 7128 18522
rect 7140 18470 7192 18522
rect 12818 18470 12870 18522
rect 12882 18470 12934 18522
rect 12946 18470 12998 18522
rect 13010 18470 13062 18522
rect 13074 18470 13126 18522
rect 18752 18470 18804 18522
rect 18816 18470 18868 18522
rect 18880 18470 18932 18522
rect 18944 18470 18996 18522
rect 19008 18470 19060 18522
rect 24686 18470 24738 18522
rect 24750 18470 24802 18522
rect 24814 18470 24866 18522
rect 24878 18470 24930 18522
rect 24942 18470 24994 18522
rect 1952 18368 2004 18420
rect 2136 18368 2188 18420
rect 3976 18368 4028 18420
rect 4252 18368 4304 18420
rect 1216 18300 1268 18352
rect 1676 18232 1728 18284
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 2320 18275 2372 18284
rect 2320 18241 2327 18275
rect 2327 18241 2361 18275
rect 2361 18241 2372 18275
rect 2320 18232 2372 18241
rect 4252 18275 4304 18284
rect 5816 18300 5868 18352
rect 4252 18241 4259 18275
rect 4259 18241 4293 18275
rect 4293 18241 4304 18275
rect 4252 18232 4304 18241
rect 5172 18232 5224 18284
rect 8300 18368 8352 18420
rect 8944 18368 8996 18420
rect 9496 18368 9548 18420
rect 8116 18300 8168 18352
rect 8484 18275 8536 18284
rect 8484 18241 8491 18275
rect 8491 18241 8525 18275
rect 8525 18241 8536 18275
rect 8484 18232 8536 18241
rect 8760 18300 8812 18352
rect 9588 18300 9640 18352
rect 10692 18300 10744 18352
rect 11796 18300 11848 18352
rect 12256 18300 12308 18352
rect 12624 18300 12676 18352
rect 12164 18232 12216 18284
rect 3976 18207 4028 18216
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 12716 18164 12768 18216
rect 13820 18300 13872 18352
rect 15292 18368 15344 18420
rect 21364 18368 21416 18420
rect 23112 18300 23164 18352
rect 14004 18232 14056 18284
rect 14464 18275 14516 18284
rect 14464 18241 14471 18275
rect 14471 18241 14505 18275
rect 14505 18241 14516 18275
rect 14464 18232 14516 18241
rect 17224 18232 17276 18284
rect 2964 18028 3016 18080
rect 4988 18071 5040 18080
rect 4988 18037 4997 18071
rect 4997 18037 5031 18071
rect 5031 18037 5040 18071
rect 4988 18028 5040 18037
rect 5356 18028 5408 18080
rect 7288 18028 7340 18080
rect 11336 18096 11388 18148
rect 13084 18096 13136 18148
rect 17500 18232 17552 18284
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 20996 18232 21048 18284
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 18052 18164 18104 18173
rect 10508 18028 10560 18080
rect 14280 18028 14332 18080
rect 17868 18096 17920 18148
rect 16120 18028 16172 18080
rect 21272 18164 21324 18216
rect 22376 18164 22428 18216
rect 19432 18028 19484 18080
rect 23572 18028 23624 18080
rect 24400 18071 24452 18080
rect 24400 18037 24409 18071
rect 24409 18037 24443 18071
rect 24443 18037 24452 18071
rect 24400 18028 24452 18037
rect 3917 17926 3969 17978
rect 3981 17926 4033 17978
rect 4045 17926 4097 17978
rect 4109 17926 4161 17978
rect 4173 17926 4225 17978
rect 9851 17926 9903 17978
rect 9915 17926 9967 17978
rect 9979 17926 10031 17978
rect 10043 17926 10095 17978
rect 10107 17926 10159 17978
rect 15785 17926 15837 17978
rect 15849 17926 15901 17978
rect 15913 17926 15965 17978
rect 15977 17926 16029 17978
rect 16041 17926 16093 17978
rect 21719 17926 21771 17978
rect 21783 17926 21835 17978
rect 21847 17926 21899 17978
rect 21911 17926 21963 17978
rect 21975 17926 22027 17978
rect 2688 17824 2740 17876
rect 2780 17824 2832 17876
rect 3700 17824 3752 17876
rect 3608 17756 3660 17808
rect 4712 17824 4764 17876
rect 3516 17688 3568 17740
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2688 17663 2740 17672
rect 2688 17629 2697 17663
rect 2697 17629 2731 17663
rect 2731 17629 2740 17663
rect 2688 17620 2740 17629
rect 2780 17663 2832 17672
rect 2780 17629 2814 17663
rect 2814 17629 2832 17663
rect 2780 17620 2832 17629
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3976 17663 4028 17672
rect 3976 17629 3985 17663
rect 3985 17629 4019 17663
rect 4019 17629 4028 17663
rect 3976 17620 4028 17629
rect 5356 17688 5408 17740
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 1952 17552 2004 17604
rect 14280 17824 14332 17876
rect 17868 17824 17920 17876
rect 22560 17824 22612 17876
rect 6000 17799 6052 17808
rect 6000 17765 6009 17799
rect 6009 17765 6043 17799
rect 6043 17765 6052 17799
rect 6000 17756 6052 17765
rect 10508 17756 10560 17808
rect 18052 17756 18104 17808
rect 3608 17527 3660 17536
rect 3608 17493 3617 17527
rect 3617 17493 3651 17527
rect 3651 17493 3660 17527
rect 3608 17484 3660 17493
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 9864 17688 9916 17740
rect 11336 17688 11388 17740
rect 12716 17731 12768 17740
rect 12716 17697 12725 17731
rect 12725 17697 12759 17731
rect 12759 17697 12768 17731
rect 12716 17688 12768 17697
rect 5816 17620 5868 17672
rect 6736 17620 6788 17672
rect 7288 17620 7340 17672
rect 10140 17620 10192 17672
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 10968 17663 11020 17672
rect 10968 17629 10977 17663
rect 10977 17629 11011 17663
rect 11011 17629 11020 17663
rect 10968 17620 11020 17629
rect 5908 17552 5960 17604
rect 5816 17484 5868 17536
rect 7472 17484 7524 17536
rect 9312 17484 9364 17536
rect 9864 17484 9916 17536
rect 10508 17484 10560 17536
rect 10876 17484 10928 17536
rect 11888 17620 11940 17672
rect 12164 17620 12216 17672
rect 13084 17663 13136 17672
rect 13084 17629 13118 17663
rect 13118 17629 13136 17663
rect 13084 17620 13136 17629
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 17132 17663 17184 17672
rect 11888 17527 11940 17536
rect 11888 17493 11897 17527
rect 11897 17493 11931 17527
rect 11931 17493 11940 17527
rect 11888 17484 11940 17493
rect 12440 17484 12492 17536
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 15476 17552 15528 17604
rect 17500 17620 17552 17672
rect 18512 17484 18564 17536
rect 19432 17552 19484 17604
rect 21272 17620 21324 17672
rect 22192 17663 22244 17672
rect 22192 17629 22201 17663
rect 22201 17629 22235 17663
rect 22235 17629 22244 17663
rect 22192 17620 22244 17629
rect 23480 17824 23532 17876
rect 19616 17484 19668 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 20720 17484 20772 17536
rect 21640 17484 21692 17536
rect 24308 17620 24360 17672
rect 24584 17620 24636 17672
rect 22468 17527 22520 17536
rect 22468 17493 22477 17527
rect 22477 17493 22511 17527
rect 22511 17493 22520 17527
rect 22468 17484 22520 17493
rect 23204 17484 23256 17536
rect 6884 17382 6936 17434
rect 6948 17382 7000 17434
rect 7012 17382 7064 17434
rect 7076 17382 7128 17434
rect 7140 17382 7192 17434
rect 12818 17382 12870 17434
rect 12882 17382 12934 17434
rect 12946 17382 12998 17434
rect 13010 17382 13062 17434
rect 13074 17382 13126 17434
rect 18752 17382 18804 17434
rect 18816 17382 18868 17434
rect 18880 17382 18932 17434
rect 18944 17382 18996 17434
rect 19008 17382 19060 17434
rect 24686 17382 24738 17434
rect 24750 17382 24802 17434
rect 24814 17382 24866 17434
rect 24878 17382 24930 17434
rect 24942 17382 24994 17434
rect 3608 17280 3660 17332
rect 4252 17280 4304 17332
rect 6368 17280 6420 17332
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 4804 17144 4856 17196
rect 5356 17212 5408 17264
rect 6460 17212 6512 17264
rect 6552 17255 6604 17264
rect 6552 17221 6561 17255
rect 6561 17221 6595 17255
rect 6595 17221 6604 17255
rect 6552 17212 6604 17221
rect 7472 17212 7524 17264
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 10508 17280 10560 17332
rect 5908 17144 5960 17196
rect 7656 17144 7708 17196
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 1952 17076 2004 17128
rect 2412 17076 2464 17128
rect 2596 17119 2648 17128
rect 2596 17085 2605 17119
rect 2605 17085 2639 17119
rect 2639 17085 2648 17119
rect 2596 17076 2648 17085
rect 4436 17076 4488 17128
rect 1584 16940 1636 16992
rect 3516 16983 3568 16992
rect 3516 16949 3525 16983
rect 3525 16949 3559 16983
rect 3559 16949 3568 16983
rect 3516 16940 3568 16949
rect 3792 16940 3844 16992
rect 9588 17212 9640 17264
rect 10968 17280 11020 17332
rect 13268 17280 13320 17332
rect 19432 17280 19484 17332
rect 8668 17144 8720 17196
rect 10232 17144 10284 17196
rect 10416 17144 10468 17196
rect 11244 17212 11296 17264
rect 12164 17212 12216 17264
rect 12256 17187 12308 17196
rect 12256 17153 12265 17187
rect 12265 17153 12299 17187
rect 12299 17153 12308 17187
rect 12256 17144 12308 17153
rect 12440 17144 12492 17196
rect 13544 17212 13596 17264
rect 14556 17212 14608 17264
rect 13728 17144 13780 17196
rect 16580 17144 16632 17196
rect 17040 17144 17092 17196
rect 20628 17280 20680 17332
rect 22192 17280 22244 17332
rect 22468 17280 22520 17332
rect 23020 17280 23072 17332
rect 25136 17280 25188 17332
rect 21088 17212 21140 17264
rect 7840 17051 7892 17060
rect 7840 17017 7849 17051
rect 7849 17017 7883 17051
rect 7883 17017 7892 17051
rect 7840 17008 7892 17017
rect 11888 17008 11940 17060
rect 10508 16940 10560 16992
rect 12440 16983 12492 16992
rect 12440 16949 12449 16983
rect 12449 16949 12483 16983
rect 12483 16949 12492 16983
rect 12440 16940 12492 16949
rect 14464 16983 14516 16992
rect 14464 16949 14473 16983
rect 14473 16949 14507 16983
rect 14507 16949 14516 16983
rect 14464 16940 14516 16949
rect 16488 17076 16540 17128
rect 19892 17076 19944 17128
rect 20444 17076 20496 17128
rect 20536 17076 20588 17128
rect 22836 17144 22888 17196
rect 23848 17187 23900 17196
rect 23848 17153 23857 17187
rect 23857 17153 23891 17187
rect 23891 17153 23900 17187
rect 23848 17144 23900 17153
rect 21824 17119 21876 17128
rect 21824 17085 21833 17119
rect 21833 17085 21867 17119
rect 21867 17085 21876 17119
rect 21824 17076 21876 17085
rect 21456 17008 21508 17060
rect 16212 16983 16264 16992
rect 16212 16949 16221 16983
rect 16221 16949 16255 16983
rect 16255 16949 16264 16983
rect 16212 16940 16264 16949
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20720 16940 20772 16992
rect 21548 16983 21600 16992
rect 21548 16949 21557 16983
rect 21557 16949 21591 16983
rect 21591 16949 21600 16983
rect 21548 16940 21600 16949
rect 24124 16983 24176 16992
rect 24124 16949 24133 16983
rect 24133 16949 24167 16983
rect 24167 16949 24176 16983
rect 24124 16940 24176 16949
rect 24400 16983 24452 16992
rect 24400 16949 24409 16983
rect 24409 16949 24443 16983
rect 24443 16949 24452 16983
rect 24400 16940 24452 16949
rect 3917 16838 3969 16890
rect 3981 16838 4033 16890
rect 4045 16838 4097 16890
rect 4109 16838 4161 16890
rect 4173 16838 4225 16890
rect 9851 16838 9903 16890
rect 9915 16838 9967 16890
rect 9979 16838 10031 16890
rect 10043 16838 10095 16890
rect 10107 16838 10159 16890
rect 15785 16838 15837 16890
rect 15849 16838 15901 16890
rect 15913 16838 15965 16890
rect 15977 16838 16029 16890
rect 16041 16838 16093 16890
rect 21719 16838 21771 16890
rect 21783 16838 21835 16890
rect 21847 16838 21899 16890
rect 21911 16838 21963 16890
rect 21975 16838 22027 16890
rect 1032 16736 1084 16788
rect 3332 16736 3384 16788
rect 4804 16736 4856 16788
rect 6000 16668 6052 16720
rect 480 16600 532 16652
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 7472 16600 7524 16652
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 9772 16668 9824 16720
rect 11060 16668 11112 16720
rect 8484 16600 8536 16652
rect 11244 16600 11296 16652
rect 16120 16736 16172 16788
rect 16212 16736 16264 16788
rect 17684 16736 17736 16788
rect 19892 16736 19944 16788
rect 20168 16736 20220 16788
rect 21456 16736 21508 16788
rect 21548 16736 21600 16788
rect 15568 16600 15620 16652
rect 15936 16643 15988 16652
rect 15936 16609 15945 16643
rect 15945 16609 15979 16643
rect 15979 16609 15988 16643
rect 15936 16600 15988 16609
rect 16028 16600 16080 16652
rect 16764 16643 16816 16652
rect 16764 16609 16798 16643
rect 16798 16609 16816 16643
rect 16764 16600 16816 16609
rect 20536 16600 20588 16652
rect 21272 16600 21324 16652
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 2136 16464 2188 16516
rect 2964 16507 3016 16516
rect 2964 16473 2973 16507
rect 2973 16473 3007 16507
rect 3007 16473 3016 16507
rect 2964 16464 3016 16473
rect 3332 16532 3384 16584
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 3792 16464 3844 16516
rect 2688 16439 2740 16448
rect 2688 16405 2697 16439
rect 2697 16405 2731 16439
rect 2731 16405 2740 16439
rect 2688 16396 2740 16405
rect 3056 16439 3108 16448
rect 3056 16405 3065 16439
rect 3065 16405 3099 16439
rect 3099 16405 3108 16439
rect 3056 16396 3108 16405
rect 3332 16396 3384 16448
rect 4252 16396 4304 16448
rect 5540 16396 5592 16448
rect 7288 16532 7340 16584
rect 7840 16575 7892 16584
rect 7840 16541 7849 16575
rect 7849 16541 7883 16575
rect 7883 16541 7892 16575
rect 7840 16532 7892 16541
rect 12532 16532 12584 16584
rect 13268 16532 13320 16584
rect 14464 16532 14516 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 17868 16532 17920 16584
rect 18604 16532 18656 16584
rect 21640 16668 21692 16720
rect 12256 16464 12308 16516
rect 14096 16396 14148 16448
rect 14648 16507 14700 16516
rect 14648 16473 14657 16507
rect 14657 16473 14691 16507
rect 14691 16473 14700 16507
rect 14648 16464 14700 16473
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 15936 16464 15988 16516
rect 20996 16396 21048 16448
rect 22928 16532 22980 16584
rect 23572 16532 23624 16584
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 21640 16396 21692 16448
rect 22100 16396 22152 16448
rect 22560 16396 22612 16448
rect 6884 16294 6936 16346
rect 6948 16294 7000 16346
rect 7012 16294 7064 16346
rect 7076 16294 7128 16346
rect 7140 16294 7192 16346
rect 12818 16294 12870 16346
rect 12882 16294 12934 16346
rect 12946 16294 12998 16346
rect 13010 16294 13062 16346
rect 13074 16294 13126 16346
rect 18752 16294 18804 16346
rect 18816 16294 18868 16346
rect 18880 16294 18932 16346
rect 18944 16294 18996 16346
rect 19008 16294 19060 16346
rect 24686 16294 24738 16346
rect 24750 16294 24802 16346
rect 24814 16294 24866 16346
rect 24878 16294 24930 16346
rect 24942 16294 24994 16346
rect 1768 16235 1820 16244
rect 1768 16201 1777 16235
rect 1777 16201 1811 16235
rect 1811 16201 1820 16235
rect 1768 16192 1820 16201
rect 2136 16192 2188 16244
rect 2964 16192 3016 16244
rect 3608 16192 3660 16244
rect 2044 16124 2096 16176
rect 2228 16124 2280 16176
rect 3332 16124 3384 16176
rect 2780 16056 2832 16108
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4528 16099 4580 16108
rect 4528 16065 4562 16099
rect 4562 16065 4580 16099
rect 4528 16056 4580 16065
rect 2964 15988 3016 16040
rect 3700 16031 3752 16040
rect 3700 15997 3709 16031
rect 3709 15997 3743 16031
rect 3743 15997 3752 16031
rect 3700 15988 3752 15997
rect 4712 16031 4764 16040
rect 4712 15997 4721 16031
rect 4721 15997 4755 16031
rect 4755 15997 4764 16031
rect 4712 15988 4764 15997
rect 4896 15988 4948 16040
rect 7012 15988 7064 16040
rect 7840 16056 7892 16108
rect 8392 16192 8444 16244
rect 8484 16235 8536 16244
rect 8484 16201 8493 16235
rect 8493 16201 8527 16235
rect 8527 16201 8536 16235
rect 8484 16192 8536 16201
rect 9036 16124 9088 16176
rect 8668 16056 8720 16108
rect 9772 16056 9824 16108
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 5448 15920 5500 15972
rect 6644 15920 6696 15972
rect 6828 15920 6880 15972
rect 3700 15852 3752 15904
rect 4620 15852 4672 15904
rect 9680 15852 9732 15904
rect 12164 16124 12216 16176
rect 12716 16192 12768 16244
rect 14648 16192 14700 16244
rect 15936 16192 15988 16244
rect 17224 16192 17276 16244
rect 10784 16056 10836 16108
rect 11244 16056 11296 16108
rect 16028 16124 16080 16176
rect 16304 16124 16356 16176
rect 17960 16124 18012 16176
rect 20720 16192 20772 16244
rect 21456 16192 21508 16244
rect 23480 16192 23532 16244
rect 23848 16192 23900 16244
rect 12716 16056 12768 16108
rect 13820 16056 13872 16108
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14700 16099
rect 14648 16056 14700 16065
rect 18880 16056 18932 16108
rect 13268 15988 13320 16040
rect 17224 15988 17276 16040
rect 17868 16031 17920 16040
rect 17868 15997 17877 16031
rect 17877 15997 17911 16031
rect 17911 15997 17920 16031
rect 17868 15988 17920 15997
rect 20996 16056 21048 16108
rect 19800 15920 19852 15972
rect 20996 15920 21048 15972
rect 15108 15852 15160 15904
rect 19524 15852 19576 15904
rect 19984 15852 20036 15904
rect 20168 15852 20220 15904
rect 24400 16056 24452 16108
rect 22560 15988 22612 16040
rect 23664 15988 23716 16040
rect 23664 15895 23716 15904
rect 23664 15861 23673 15895
rect 23673 15861 23707 15895
rect 23707 15861 23716 15895
rect 23664 15852 23716 15861
rect 3917 15750 3969 15802
rect 3981 15750 4033 15802
rect 4045 15750 4097 15802
rect 4109 15750 4161 15802
rect 4173 15750 4225 15802
rect 9851 15750 9903 15802
rect 9915 15750 9967 15802
rect 9979 15750 10031 15802
rect 10043 15750 10095 15802
rect 10107 15750 10159 15802
rect 15785 15750 15837 15802
rect 15849 15750 15901 15802
rect 15913 15750 15965 15802
rect 15977 15750 16029 15802
rect 16041 15750 16093 15802
rect 21719 15750 21771 15802
rect 21783 15750 21835 15802
rect 21847 15750 21899 15802
rect 21911 15750 21963 15802
rect 21975 15750 22027 15802
rect 2872 15691 2924 15700
rect 2872 15657 2881 15691
rect 2881 15657 2915 15691
rect 2915 15657 2924 15691
rect 2872 15648 2924 15657
rect 3240 15444 3292 15496
rect 4620 15648 4672 15700
rect 4712 15648 4764 15700
rect 7564 15648 7616 15700
rect 9680 15648 9732 15700
rect 10600 15648 10652 15700
rect 12348 15648 12400 15700
rect 16764 15648 16816 15700
rect 18880 15648 18932 15700
rect 3700 15512 3752 15564
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 6368 15512 6420 15564
rect 6828 15555 6880 15564
rect 6828 15521 6837 15555
rect 6837 15521 6871 15555
rect 6871 15521 6880 15555
rect 6828 15512 6880 15521
rect 9036 15512 9088 15564
rect 9312 15512 9364 15564
rect 9680 15512 9732 15564
rect 13360 15512 13412 15564
rect 23848 15648 23900 15700
rect 24124 15691 24176 15700
rect 24124 15657 24133 15691
rect 24133 15657 24167 15691
rect 24167 15657 24176 15691
rect 24124 15648 24176 15657
rect 21640 15580 21692 15632
rect 3516 15444 3568 15496
rect 4160 15444 4212 15496
rect 5356 15444 5408 15496
rect 2320 15351 2372 15360
rect 2320 15317 2329 15351
rect 2329 15317 2363 15351
rect 2363 15317 2372 15351
rect 2320 15308 2372 15317
rect 3240 15351 3292 15360
rect 3240 15317 3249 15351
rect 3249 15317 3283 15351
rect 3283 15317 3292 15351
rect 3240 15308 3292 15317
rect 3700 15308 3752 15360
rect 6368 15308 6420 15360
rect 6552 15308 6604 15360
rect 7012 15444 7064 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 7380 15376 7432 15428
rect 7748 15376 7800 15428
rect 11244 15376 11296 15428
rect 11428 15376 11480 15428
rect 11612 15444 11664 15496
rect 16856 15444 16908 15496
rect 17960 15444 18012 15496
rect 11704 15376 11756 15428
rect 14096 15376 14148 15428
rect 19892 15444 19944 15496
rect 20168 15444 20220 15496
rect 21180 15444 21232 15496
rect 22192 15444 22244 15496
rect 19340 15376 19392 15428
rect 22468 15444 22520 15496
rect 10968 15308 11020 15360
rect 11888 15351 11940 15360
rect 11888 15317 11897 15351
rect 11897 15317 11931 15351
rect 11931 15317 11940 15351
rect 11888 15308 11940 15317
rect 13544 15308 13596 15360
rect 15292 15308 15344 15360
rect 17960 15308 18012 15360
rect 19800 15308 19852 15360
rect 22744 15308 22796 15360
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 6884 15206 6936 15258
rect 6948 15206 7000 15258
rect 7012 15206 7064 15258
rect 7076 15206 7128 15258
rect 7140 15206 7192 15258
rect 12818 15206 12870 15258
rect 12882 15206 12934 15258
rect 12946 15206 12998 15258
rect 13010 15206 13062 15258
rect 13074 15206 13126 15258
rect 18752 15206 18804 15258
rect 18816 15206 18868 15258
rect 18880 15206 18932 15258
rect 18944 15206 18996 15258
rect 19008 15206 19060 15258
rect 24686 15206 24738 15258
rect 24750 15206 24802 15258
rect 24814 15206 24866 15258
rect 24878 15206 24930 15258
rect 24942 15206 24994 15258
rect 2136 15104 2188 15156
rect 2320 15036 2372 15088
rect 3148 15036 3200 15088
rect 3240 15036 3292 15088
rect 4160 15036 4212 15088
rect 1768 15011 1820 15020
rect 1768 14977 1777 15011
rect 1777 14977 1811 15011
rect 1811 14977 1820 15011
rect 1768 14968 1820 14977
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 4620 15104 4672 15156
rect 7288 15104 7340 15156
rect 8852 15104 8904 15156
rect 9956 15104 10008 15156
rect 10140 15104 10192 15156
rect 4988 14968 5040 15020
rect 9312 15036 9364 15088
rect 9680 15036 9732 15088
rect 11796 15036 11848 15088
rect 12624 15104 12676 15156
rect 13176 15104 13228 15156
rect 13544 15104 13596 15156
rect 14648 15104 14700 15156
rect 16396 15104 16448 15156
rect 7472 14968 7524 15020
rect 8668 14968 8720 15020
rect 10232 14968 10284 15020
rect 10876 14968 10928 15020
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12348 14968 12400 15020
rect 13728 14968 13780 15020
rect 14096 14968 14148 15020
rect 17592 15104 17644 15156
rect 19340 15104 19392 15156
rect 22468 15104 22520 15156
rect 22744 15104 22796 15156
rect 17224 15036 17276 15088
rect 17776 15036 17828 15088
rect 17868 15036 17920 15088
rect 19616 15036 19668 15088
rect 18512 14968 18564 15020
rect 6368 14943 6420 14952
rect 1308 14764 1360 14816
rect 2872 14807 2924 14816
rect 2872 14773 2881 14807
rect 2881 14773 2915 14807
rect 2915 14773 2924 14807
rect 2872 14764 2924 14773
rect 3056 14764 3108 14816
rect 3976 14807 4028 14816
rect 3976 14773 3985 14807
rect 3985 14773 4019 14807
rect 4019 14773 4028 14807
rect 3976 14764 4028 14773
rect 4804 14764 4856 14816
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 6920 14900 6972 14952
rect 5080 14832 5132 14884
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 5356 14764 5408 14773
rect 5908 14832 5960 14884
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 7748 14900 7800 14952
rect 11888 14900 11940 14952
rect 13912 14943 13964 14952
rect 13912 14909 13921 14943
rect 13921 14909 13955 14943
rect 13955 14909 13964 14943
rect 13912 14900 13964 14909
rect 19524 15011 19576 15020
rect 19524 14977 19533 15011
rect 19533 14977 19567 15011
rect 19567 14977 19576 15011
rect 19524 14968 19576 14977
rect 19800 15011 19852 15020
rect 19800 14977 19809 15011
rect 19809 14977 19843 15011
rect 19843 14977 19852 15011
rect 19800 14968 19852 14977
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 21180 15036 21232 15088
rect 20812 14968 20864 15020
rect 24216 15104 24268 15156
rect 23664 14968 23716 15020
rect 24216 15011 24268 15020
rect 24216 14977 24225 15011
rect 24225 14977 24259 15011
rect 24259 14977 24268 15011
rect 24216 14968 24268 14977
rect 21272 14900 21324 14952
rect 21548 14900 21600 14952
rect 22836 14900 22888 14952
rect 20260 14832 20312 14884
rect 8668 14764 8720 14816
rect 11428 14764 11480 14816
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 22192 14764 22244 14816
rect 22560 14764 22612 14816
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 3917 14662 3969 14714
rect 3981 14662 4033 14714
rect 4045 14662 4097 14714
rect 4109 14662 4161 14714
rect 4173 14662 4225 14714
rect 9851 14662 9903 14714
rect 9915 14662 9967 14714
rect 9979 14662 10031 14714
rect 10043 14662 10095 14714
rect 10107 14662 10159 14714
rect 15785 14662 15837 14714
rect 15849 14662 15901 14714
rect 15913 14662 15965 14714
rect 15977 14662 16029 14714
rect 16041 14662 16093 14714
rect 21719 14662 21771 14714
rect 21783 14662 21835 14714
rect 21847 14662 21899 14714
rect 21911 14662 21963 14714
rect 21975 14662 22027 14714
rect 2872 14560 2924 14612
rect 3516 14492 3568 14544
rect 2872 14424 2924 14476
rect 1308 14356 1360 14408
rect 2136 14356 2188 14408
rect 2688 14399 2740 14408
rect 2688 14365 2697 14399
rect 2697 14365 2731 14399
rect 2731 14365 2740 14399
rect 2688 14356 2740 14365
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 5080 14560 5132 14612
rect 5908 14560 5960 14612
rect 5356 14492 5408 14544
rect 6552 14492 6604 14544
rect 6828 14492 6880 14544
rect 7564 14560 7616 14612
rect 10508 14560 10560 14612
rect 12072 14560 12124 14612
rect 12348 14560 12400 14612
rect 4436 14424 4488 14476
rect 5448 14424 5500 14476
rect 5908 14424 5960 14476
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 4620 14356 4672 14408
rect 4804 14356 4856 14408
rect 2688 14220 2740 14272
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 4988 14288 5040 14340
rect 5816 14399 5868 14408
rect 5816 14365 5825 14399
rect 5825 14365 5859 14399
rect 5859 14365 5868 14399
rect 5816 14356 5868 14365
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 7564 14424 7616 14476
rect 8208 14424 8260 14476
rect 11244 14467 11296 14476
rect 11244 14433 11253 14467
rect 11253 14433 11287 14467
rect 11287 14433 11296 14467
rect 11244 14424 11296 14433
rect 6736 14356 6788 14408
rect 7012 14356 7064 14408
rect 7472 14356 7524 14408
rect 10876 14356 10928 14408
rect 11520 14399 11572 14408
rect 11520 14365 11527 14399
rect 11527 14365 11561 14399
rect 11561 14365 11572 14399
rect 11520 14356 11572 14365
rect 12624 14399 12676 14408
rect 12624 14365 12633 14399
rect 12633 14365 12667 14399
rect 12667 14365 12676 14399
rect 12624 14356 12676 14365
rect 14924 14560 14976 14612
rect 13360 14492 13412 14544
rect 13636 14492 13688 14544
rect 14740 14492 14792 14544
rect 13728 14424 13780 14476
rect 16580 14560 16632 14612
rect 16948 14560 17000 14612
rect 18512 14560 18564 14612
rect 20260 14560 20312 14612
rect 25504 14696 25556 14748
rect 16120 14424 16172 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 17224 14467 17276 14476
rect 17224 14433 17258 14467
rect 17258 14433 17276 14467
rect 17224 14424 17276 14433
rect 17776 14424 17828 14476
rect 4344 14220 4396 14272
rect 11888 14288 11940 14340
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 16304 14356 16356 14408
rect 16396 14399 16448 14408
rect 16396 14365 16405 14399
rect 16405 14365 16439 14399
rect 16439 14365 16448 14399
rect 16396 14356 16448 14365
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 17408 14399 17460 14408
rect 17408 14365 17417 14399
rect 17417 14365 17451 14399
rect 17451 14365 17460 14399
rect 17408 14356 17460 14365
rect 22468 14492 22520 14544
rect 12072 14220 12124 14272
rect 16120 14331 16172 14340
rect 16120 14297 16129 14331
rect 16129 14297 16163 14331
rect 16163 14297 16172 14331
rect 16120 14288 16172 14297
rect 13176 14220 13228 14272
rect 17316 14220 17368 14272
rect 17868 14220 17920 14272
rect 22192 14356 22244 14408
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 25136 14492 25188 14544
rect 23756 14424 23808 14476
rect 18512 14263 18564 14272
rect 18512 14229 18521 14263
rect 18521 14229 18555 14263
rect 18555 14229 18564 14263
rect 18512 14220 18564 14229
rect 19156 14220 19208 14272
rect 21640 14220 21692 14272
rect 22744 14220 22796 14272
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 24124 14288 24176 14340
rect 24216 14220 24268 14272
rect 6884 14118 6936 14170
rect 6948 14118 7000 14170
rect 7012 14118 7064 14170
rect 7076 14118 7128 14170
rect 7140 14118 7192 14170
rect 12818 14118 12870 14170
rect 12882 14118 12934 14170
rect 12946 14118 12998 14170
rect 13010 14118 13062 14170
rect 13074 14118 13126 14170
rect 18752 14118 18804 14170
rect 18816 14118 18868 14170
rect 18880 14118 18932 14170
rect 18944 14118 18996 14170
rect 19008 14118 19060 14170
rect 24686 14118 24738 14170
rect 24750 14118 24802 14170
rect 24814 14118 24866 14170
rect 24878 14118 24930 14170
rect 24942 14118 24994 14170
rect 1400 14016 1452 14068
rect 2964 14016 3016 14068
rect 6092 14016 6144 14068
rect 6368 14016 6420 14068
rect 12164 14016 12216 14068
rect 12624 14016 12676 14068
rect 12808 14016 12860 14068
rect 13912 14016 13964 14068
rect 6552 13948 6604 14000
rect 7472 13948 7524 14000
rect 11704 13948 11756 14000
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 15292 14016 15344 14068
rect 15476 14016 15528 14068
rect 16764 14016 16816 14068
rect 1952 13880 2004 13932
rect 2412 13880 2464 13932
rect 3700 13923 3752 13932
rect 3700 13889 3709 13923
rect 3709 13889 3743 13923
rect 3743 13889 3752 13923
rect 3700 13880 3752 13889
rect 4344 13923 4396 13932
rect 4344 13889 4353 13923
rect 4353 13889 4387 13923
rect 4387 13889 4396 13923
rect 4344 13880 4396 13889
rect 5080 13880 5132 13932
rect 5264 13880 5316 13932
rect 6736 13880 6788 13932
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2320 13676 2372 13728
rect 2964 13744 3016 13796
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 8116 13880 8168 13932
rect 8852 13880 8904 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9916 13923
rect 9864 13880 9916 13889
rect 7840 13719 7892 13728
rect 7840 13685 7849 13719
rect 7849 13685 7883 13719
rect 7883 13685 7892 13719
rect 7840 13676 7892 13685
rect 9312 13812 9364 13864
rect 12624 13855 12676 13864
rect 12624 13821 12633 13855
rect 12633 13821 12667 13855
rect 12667 13821 12676 13855
rect 12624 13812 12676 13821
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 8944 13744 8996 13796
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 10416 13676 10468 13728
rect 10508 13676 10560 13728
rect 13176 13812 13228 13864
rect 13544 13846 13596 13898
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 14556 13812 14608 13864
rect 15200 13948 15252 14000
rect 17408 14016 17460 14068
rect 17776 14016 17828 14068
rect 20812 14016 20864 14068
rect 22284 14016 22336 14068
rect 23020 14016 23072 14068
rect 23112 14016 23164 14068
rect 14924 13919 14949 13932
rect 14949 13919 14976 13932
rect 14924 13880 14976 13919
rect 16120 13880 16172 13932
rect 16488 13880 16540 13932
rect 18144 13948 18196 14000
rect 14556 13676 14608 13728
rect 17408 13880 17460 13932
rect 19156 13948 19208 14000
rect 22836 13991 22888 14000
rect 22836 13957 22845 13991
rect 22845 13957 22879 13991
rect 22879 13957 22888 13991
rect 22836 13948 22888 13957
rect 17960 13812 18012 13864
rect 20904 13880 20956 13932
rect 22468 13880 22520 13932
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 19156 13812 19208 13864
rect 23112 13880 23164 13932
rect 23296 13880 23348 13932
rect 23388 13855 23440 13864
rect 23388 13821 23397 13855
rect 23397 13821 23431 13855
rect 23431 13821 23440 13855
rect 23388 13812 23440 13821
rect 18880 13744 18932 13796
rect 20444 13744 20496 13796
rect 21272 13676 21324 13728
rect 23480 13787 23532 13796
rect 23480 13753 23489 13787
rect 23489 13753 23523 13787
rect 23523 13753 23532 13787
rect 23480 13744 23532 13753
rect 24400 13719 24452 13728
rect 24400 13685 24409 13719
rect 24409 13685 24443 13719
rect 24443 13685 24452 13719
rect 24400 13676 24452 13685
rect 3917 13574 3969 13626
rect 3981 13574 4033 13626
rect 4045 13574 4097 13626
rect 4109 13574 4161 13626
rect 4173 13574 4225 13626
rect 9851 13574 9903 13626
rect 9915 13574 9967 13626
rect 9979 13574 10031 13626
rect 10043 13574 10095 13626
rect 10107 13574 10159 13626
rect 15785 13574 15837 13626
rect 15849 13574 15901 13626
rect 15913 13574 15965 13626
rect 15977 13574 16029 13626
rect 16041 13574 16093 13626
rect 21719 13574 21771 13626
rect 21783 13574 21835 13626
rect 21847 13574 21899 13626
rect 21911 13574 21963 13626
rect 21975 13574 22027 13626
rect 1216 13472 1268 13524
rect 2780 13472 2832 13524
rect 9128 13472 9180 13524
rect 1676 13447 1728 13456
rect 1676 13413 1685 13447
rect 1685 13413 1719 13447
rect 1719 13413 1728 13447
rect 1676 13404 1728 13413
rect 8208 13404 8260 13456
rect 8392 13404 8444 13456
rect 2044 13336 2096 13388
rect 3240 13336 3292 13388
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 7288 13336 7340 13388
rect 8944 13336 8996 13388
rect 10416 13472 10468 13524
rect 10140 13336 10192 13388
rect 10784 13472 10836 13524
rect 11428 13472 11480 13524
rect 12716 13472 12768 13524
rect 296 13200 348 13252
rect 848 13200 900 13252
rect 1584 13200 1636 13252
rect 2780 13243 2832 13252
rect 2780 13209 2789 13243
rect 2789 13209 2823 13243
rect 2823 13209 2832 13243
rect 2780 13200 2832 13209
rect 3516 13268 3568 13320
rect 4068 13311 4120 13320
rect 4068 13277 4093 13311
rect 4093 13277 4120 13311
rect 4068 13268 4120 13277
rect 4436 13268 4488 13320
rect 5448 13268 5500 13320
rect 8024 13268 8076 13320
rect 9496 13293 9505 13320
rect 9505 13293 9539 13320
rect 9539 13293 9548 13320
rect 9496 13268 9548 13293
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 3792 13132 3844 13184
rect 4436 13132 4488 13184
rect 5264 13132 5316 13184
rect 8392 13132 8444 13184
rect 9956 13200 10008 13252
rect 12164 13336 12216 13388
rect 12348 13336 12400 13388
rect 13636 13515 13688 13524
rect 13636 13481 13645 13515
rect 13645 13481 13679 13515
rect 13679 13481 13688 13515
rect 13636 13472 13688 13481
rect 11612 13268 11664 13320
rect 12808 13268 12860 13320
rect 13820 13268 13872 13320
rect 16856 13472 16908 13524
rect 18512 13472 18564 13524
rect 20444 13472 20496 13524
rect 23204 13472 23256 13524
rect 16948 13404 17000 13456
rect 19524 13404 19576 13456
rect 16488 13336 16540 13388
rect 18972 13336 19024 13388
rect 15200 13268 15252 13320
rect 17776 13268 17828 13320
rect 18880 13268 18932 13320
rect 13544 13200 13596 13252
rect 13636 13200 13688 13252
rect 20352 13311 20404 13320
rect 20352 13277 20361 13311
rect 20361 13277 20395 13311
rect 20395 13277 20404 13311
rect 20352 13268 20404 13277
rect 22284 13447 22336 13456
rect 22284 13413 22293 13447
rect 22293 13413 22327 13447
rect 22327 13413 22336 13447
rect 22284 13404 22336 13413
rect 20812 13311 20864 13320
rect 20812 13277 20821 13311
rect 20821 13277 20855 13311
rect 20855 13277 20864 13311
rect 20812 13268 20864 13277
rect 21180 13268 21232 13320
rect 20168 13243 20220 13252
rect 20168 13209 20177 13243
rect 20177 13209 20211 13243
rect 20211 13209 20220 13243
rect 20168 13200 20220 13209
rect 23480 13268 23532 13320
rect 19248 13132 19300 13184
rect 19340 13132 19392 13184
rect 21456 13132 21508 13184
rect 23204 13200 23256 13252
rect 6884 13030 6936 13082
rect 6948 13030 7000 13082
rect 7012 13030 7064 13082
rect 7076 13030 7128 13082
rect 7140 13030 7192 13082
rect 12818 13030 12870 13082
rect 12882 13030 12934 13082
rect 12946 13030 12998 13082
rect 13010 13030 13062 13082
rect 13074 13030 13126 13082
rect 18752 13030 18804 13082
rect 18816 13030 18868 13082
rect 18880 13030 18932 13082
rect 18944 13030 18996 13082
rect 19008 13030 19060 13082
rect 24686 13030 24738 13082
rect 24750 13030 24802 13082
rect 24814 13030 24866 13082
rect 24878 13030 24930 13082
rect 24942 13030 24994 13082
rect 3792 12928 3844 12980
rect 4344 12928 4396 12980
rect 5540 12928 5592 12980
rect 5816 12928 5868 12980
rect 6000 12928 6052 12980
rect 6828 12928 6880 12980
rect 7196 12928 7248 12980
rect 7932 12928 7984 12980
rect 9496 12928 9548 12980
rect 9956 12928 10008 12980
rect 10232 12928 10284 12980
rect 10876 12928 10928 12980
rect 10968 12928 11020 12980
rect 1860 12903 1912 12912
rect 1860 12869 1869 12903
rect 1869 12869 1903 12903
rect 1903 12869 1912 12903
rect 1860 12860 1912 12869
rect 2412 12860 2464 12912
rect 2964 12860 3016 12912
rect 3884 12860 3936 12912
rect 20168 12928 20220 12980
rect 20812 12928 20864 12980
rect 22192 12971 22244 12980
rect 22192 12937 22201 12971
rect 22201 12937 22235 12971
rect 22235 12937 22244 12971
rect 22192 12928 22244 12937
rect 22652 12928 22704 12980
rect 23388 12971 23440 12980
rect 23388 12937 23397 12971
rect 23397 12937 23431 12971
rect 23431 12937 23440 12971
rect 23388 12928 23440 12937
rect 2228 12656 2280 12708
rect 3240 12792 3292 12844
rect 4712 12835 4764 12844
rect 4712 12801 4746 12835
rect 4746 12801 4764 12835
rect 4712 12792 4764 12801
rect 4896 12835 4948 12844
rect 4896 12801 4905 12835
rect 4905 12801 4939 12835
rect 4939 12801 4948 12835
rect 4896 12792 4948 12801
rect 3056 12724 3108 12776
rect 3332 12724 3384 12776
rect 4068 12724 4120 12776
rect 4436 12724 4488 12776
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 12348 12860 12400 12912
rect 13728 12860 13780 12912
rect 6276 12792 6328 12844
rect 7288 12792 7340 12844
rect 8024 12835 8076 12844
rect 4620 12724 4672 12733
rect 2044 12588 2096 12640
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 6092 12656 6144 12708
rect 7104 12656 7156 12708
rect 6276 12588 6328 12640
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 9036 12835 9088 12844
rect 9036 12801 9070 12835
rect 9070 12801 9088 12835
rect 9036 12792 9088 12801
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 10416 12792 10468 12844
rect 11612 12792 11664 12844
rect 11888 12792 11940 12844
rect 15016 12860 15068 12912
rect 17040 12865 17092 12912
rect 17040 12860 17065 12865
rect 17065 12860 17092 12865
rect 7840 12724 7892 12776
rect 8392 12724 8444 12776
rect 8760 12724 8812 12776
rect 8300 12588 8352 12640
rect 8760 12588 8812 12640
rect 9312 12588 9364 12640
rect 11244 12656 11296 12708
rect 10968 12588 11020 12640
rect 17960 12792 18012 12844
rect 19340 12860 19392 12912
rect 18604 12792 18656 12844
rect 21180 12860 21232 12912
rect 22376 12860 22428 12912
rect 13820 12724 13872 12776
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 19248 12699 19300 12708
rect 19248 12665 19257 12699
rect 19257 12665 19291 12699
rect 19291 12665 19300 12699
rect 19248 12656 19300 12665
rect 22192 12792 22244 12844
rect 24400 12860 24452 12912
rect 22100 12656 22152 12708
rect 17132 12588 17184 12640
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 20352 12588 20404 12640
rect 21456 12588 21508 12640
rect 22652 12588 22704 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 3917 12486 3969 12538
rect 3981 12486 4033 12538
rect 4045 12486 4097 12538
rect 4109 12486 4161 12538
rect 4173 12486 4225 12538
rect 9851 12486 9903 12538
rect 9915 12486 9967 12538
rect 9979 12486 10031 12538
rect 10043 12486 10095 12538
rect 10107 12486 10159 12538
rect 15785 12486 15837 12538
rect 15849 12486 15901 12538
rect 15913 12486 15965 12538
rect 15977 12486 16029 12538
rect 16041 12486 16093 12538
rect 21719 12486 21771 12538
rect 21783 12486 21835 12538
rect 21847 12486 21899 12538
rect 21911 12486 21963 12538
rect 21975 12486 22027 12538
rect 3516 12384 3568 12436
rect 4988 12316 5040 12368
rect 6000 12384 6052 12436
rect 1308 12248 1360 12300
rect 2136 12248 2188 12300
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 2504 12248 2556 12300
rect 2872 12248 2924 12300
rect 3332 12248 3384 12300
rect 5448 12248 5500 12300
rect 5908 12248 5960 12300
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 6920 12248 6972 12300
rect 4344 12180 4396 12232
rect 4528 12180 4580 12232
rect 5264 12180 5316 12232
rect 9772 12384 9824 12436
rect 21548 12384 21600 12436
rect 22284 12384 22336 12436
rect 7472 12359 7524 12368
rect 7472 12325 7481 12359
rect 7481 12325 7515 12359
rect 7515 12325 7524 12359
rect 7472 12316 7524 12325
rect 16304 12316 16356 12368
rect 3516 12044 3568 12096
rect 3700 12044 3752 12096
rect 5908 12044 5960 12096
rect 7196 12180 7248 12232
rect 7840 12291 7892 12300
rect 7840 12257 7874 12291
rect 7874 12257 7892 12291
rect 7840 12248 7892 12257
rect 12532 12248 12584 12300
rect 13912 12248 13964 12300
rect 17040 12291 17092 12300
rect 17040 12257 17049 12291
rect 17049 12257 17083 12291
rect 17083 12257 17092 12291
rect 17040 12248 17092 12257
rect 17776 12248 17828 12300
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 12716 12180 12768 12232
rect 12808 12180 12860 12232
rect 14464 12180 14516 12232
rect 14924 12180 14976 12232
rect 9036 12112 9088 12164
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 8300 12044 8352 12096
rect 11612 12044 11664 12096
rect 12164 12112 12216 12164
rect 12348 12112 12400 12164
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 14004 12112 14056 12164
rect 14740 12112 14792 12164
rect 14188 12044 14240 12096
rect 14464 12044 14516 12096
rect 16488 12180 16540 12232
rect 16764 12180 16816 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20220 12223
rect 20168 12180 20220 12189
rect 21272 12223 21324 12232
rect 21272 12189 21281 12223
rect 21281 12189 21315 12223
rect 21315 12189 21324 12223
rect 21272 12180 21324 12189
rect 20812 12112 20864 12164
rect 22100 12180 22152 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 25136 12384 25188 12436
rect 25228 12316 25280 12368
rect 25688 12248 25740 12300
rect 21640 12112 21692 12164
rect 23848 12180 23900 12232
rect 15384 12087 15436 12096
rect 15384 12053 15393 12087
rect 15393 12053 15427 12087
rect 15427 12053 15436 12087
rect 15384 12044 15436 12053
rect 16396 12044 16448 12096
rect 16580 12044 16632 12096
rect 21824 12044 21876 12096
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 23112 12087 23164 12096
rect 23112 12053 23121 12087
rect 23121 12053 23155 12087
rect 23155 12053 23164 12087
rect 23112 12044 23164 12053
rect 6884 11942 6936 11994
rect 6948 11942 7000 11994
rect 7012 11942 7064 11994
rect 7076 11942 7128 11994
rect 7140 11942 7192 11994
rect 12818 11942 12870 11994
rect 12882 11942 12934 11994
rect 12946 11942 12998 11994
rect 13010 11942 13062 11994
rect 13074 11942 13126 11994
rect 18752 11942 18804 11994
rect 18816 11942 18868 11994
rect 18880 11942 18932 11994
rect 18944 11942 18996 11994
rect 19008 11942 19060 11994
rect 24686 11942 24738 11994
rect 24750 11942 24802 11994
rect 24814 11942 24866 11994
rect 24878 11942 24930 11994
rect 24942 11942 24994 11994
rect 2412 11840 2464 11892
rect 3516 11840 3568 11892
rect 3700 11840 3752 11892
rect 4896 11840 4948 11892
rect 6000 11840 6052 11892
rect 3332 11704 3384 11756
rect 3516 11747 3568 11756
rect 3516 11713 3525 11747
rect 3525 11713 3559 11747
rect 3559 11713 3568 11747
rect 3516 11704 3568 11713
rect 3884 11704 3936 11756
rect 2228 11500 2280 11552
rect 2596 11500 2648 11552
rect 5264 11704 5316 11756
rect 6828 11704 6880 11756
rect 7840 11840 7892 11892
rect 8024 11840 8076 11892
rect 12532 11883 12584 11892
rect 12532 11849 12541 11883
rect 12541 11849 12575 11883
rect 12575 11849 12584 11883
rect 12532 11840 12584 11849
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 7288 11772 7340 11824
rect 8944 11772 8996 11824
rect 4712 11636 4764 11688
rect 8484 11704 8536 11756
rect 5356 11500 5408 11552
rect 8300 11500 8352 11552
rect 9128 11568 9180 11620
rect 10600 11568 10652 11620
rect 8576 11500 8628 11552
rect 8760 11500 8812 11552
rect 9680 11500 9732 11552
rect 11244 11704 11296 11756
rect 12072 11772 12124 11824
rect 14556 11772 14608 11824
rect 13544 11704 13596 11756
rect 15200 11747 15252 11756
rect 15200 11713 15207 11747
rect 15207 11713 15241 11747
rect 15241 11713 15252 11747
rect 15200 11704 15252 11713
rect 16488 11704 16540 11756
rect 17132 11772 17184 11824
rect 16856 11704 16908 11756
rect 17040 11704 17092 11756
rect 22744 11840 22796 11892
rect 22836 11840 22888 11892
rect 23112 11840 23164 11892
rect 23480 11840 23532 11892
rect 17868 11704 17920 11756
rect 17960 11704 18012 11756
rect 21640 11747 21692 11756
rect 21640 11713 21649 11747
rect 21649 11713 21683 11747
rect 21683 11713 21692 11747
rect 21640 11704 21692 11713
rect 21732 11704 21784 11756
rect 21824 11636 21876 11688
rect 23204 11704 23256 11756
rect 23480 11704 23532 11756
rect 12900 11568 12952 11620
rect 16304 11500 16356 11552
rect 19156 11568 19208 11620
rect 18328 11500 18380 11552
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 25228 11500 25280 11552
rect 3917 11398 3969 11450
rect 3981 11398 4033 11450
rect 4045 11398 4097 11450
rect 4109 11398 4161 11450
rect 4173 11398 4225 11450
rect 9851 11398 9903 11450
rect 9915 11398 9967 11450
rect 9979 11398 10031 11450
rect 10043 11398 10095 11450
rect 10107 11398 10159 11450
rect 15785 11398 15837 11450
rect 15849 11398 15901 11450
rect 15913 11398 15965 11450
rect 15977 11398 16029 11450
rect 16041 11398 16093 11450
rect 21719 11398 21771 11450
rect 21783 11398 21835 11450
rect 21847 11398 21899 11450
rect 21911 11398 21963 11450
rect 21975 11398 22027 11450
rect 1768 11339 1820 11348
rect 1768 11305 1777 11339
rect 1777 11305 1811 11339
rect 1811 11305 1820 11339
rect 1768 11296 1820 11305
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3608 11296 3660 11348
rect 3148 11228 3200 11280
rect 6736 11296 6788 11348
rect 7472 11296 7524 11348
rect 10048 11296 10100 11348
rect 1952 11092 2004 11144
rect 480 11024 532 11076
rect 2228 11067 2280 11076
rect 2228 11033 2237 11067
rect 2237 11033 2271 11067
rect 2271 11033 2280 11067
rect 2228 11024 2280 11033
rect 2780 11024 2832 11076
rect 4252 11024 4304 11076
rect 6828 11092 6880 11144
rect 7012 11092 7064 11144
rect 9036 11228 9088 11280
rect 12900 11228 12952 11280
rect 15108 11228 15160 11280
rect 9680 11160 9732 11212
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 15752 11228 15804 11280
rect 15844 11271 15896 11280
rect 15844 11237 15853 11271
rect 15853 11237 15887 11271
rect 15887 11237 15896 11271
rect 15844 11228 15896 11237
rect 9864 11160 9916 11169
rect 16120 11203 16172 11212
rect 16120 11169 16129 11203
rect 16129 11169 16163 11203
rect 16163 11169 16172 11203
rect 16120 11160 16172 11169
rect 16212 11203 16264 11212
rect 16212 11169 16246 11203
rect 16246 11169 16264 11203
rect 16212 11160 16264 11169
rect 18328 11296 18380 11348
rect 19064 11296 19116 11348
rect 19616 11296 19668 11348
rect 21088 11296 21140 11348
rect 7840 11092 7892 11144
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 9312 11092 9364 11144
rect 9956 11135 10008 11144
rect 9956 11101 9990 11135
rect 9990 11101 10008 11135
rect 9956 11092 10008 11101
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 8024 11024 8076 11076
rect 1492 10956 1544 11008
rect 2688 10956 2740 11008
rect 3056 10999 3108 11008
rect 3056 10965 3065 10999
rect 3065 10965 3099 10999
rect 3099 10965 3108 10999
rect 3056 10956 3108 10965
rect 3424 10999 3476 11008
rect 3424 10965 3433 10999
rect 3433 10965 3467 10999
rect 3467 10965 3476 10999
rect 3424 10956 3476 10965
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 4528 10956 4580 11008
rect 5356 10956 5408 11008
rect 7288 10956 7340 11008
rect 8116 10956 8168 11008
rect 12532 11024 12584 11076
rect 14924 11024 14976 11076
rect 17132 11135 17184 11144
rect 17132 11101 17141 11135
rect 17141 11101 17175 11135
rect 17175 11101 17184 11135
rect 17132 11092 17184 11101
rect 17408 11135 17460 11144
rect 17408 11101 17415 11135
rect 17415 11101 17449 11135
rect 17449 11101 17460 11135
rect 17408 11092 17460 11101
rect 17776 11092 17828 11144
rect 18604 11092 18656 11144
rect 19892 11092 19944 11144
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 17040 11024 17092 11076
rect 16856 10956 16908 11008
rect 21364 11024 21416 11076
rect 23204 11296 23256 11348
rect 23480 11296 23532 11348
rect 22468 11092 22520 11144
rect 22652 11092 22704 11144
rect 22928 11092 22980 11144
rect 22284 10956 22336 11008
rect 22744 10956 22796 11008
rect 6884 10854 6936 10906
rect 6948 10854 7000 10906
rect 7012 10854 7064 10906
rect 7076 10854 7128 10906
rect 7140 10854 7192 10906
rect 12818 10854 12870 10906
rect 12882 10854 12934 10906
rect 12946 10854 12998 10906
rect 13010 10854 13062 10906
rect 13074 10854 13126 10906
rect 18752 10854 18804 10906
rect 18816 10854 18868 10906
rect 18880 10854 18932 10906
rect 18944 10854 18996 10906
rect 19008 10854 19060 10906
rect 24686 10854 24738 10906
rect 24750 10854 24802 10906
rect 24814 10854 24866 10906
rect 24878 10854 24930 10906
rect 24942 10854 24994 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2228 10752 2280 10804
rect 4712 10752 4764 10804
rect 5816 10752 5868 10804
rect 6184 10752 6236 10804
rect 6552 10752 6604 10804
rect 7380 10752 7432 10804
rect 9496 10752 9548 10804
rect 10140 10752 10192 10804
rect 1492 10727 1544 10736
rect 1492 10693 1501 10727
rect 1501 10693 1535 10727
rect 1535 10693 1544 10727
rect 1492 10684 1544 10693
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 3516 10480 3568 10532
rect 1952 10455 2004 10464
rect 1952 10421 1961 10455
rect 1961 10421 1995 10455
rect 1995 10421 2004 10455
rect 1952 10412 2004 10421
rect 2320 10412 2372 10464
rect 5816 10616 5868 10668
rect 6552 10616 6604 10668
rect 8576 10616 8628 10668
rect 9588 10684 9640 10736
rect 16212 10752 16264 10804
rect 13636 10727 13688 10736
rect 13636 10693 13645 10727
rect 13645 10693 13679 10727
rect 13679 10693 13688 10727
rect 13636 10684 13688 10693
rect 14188 10684 14240 10736
rect 9404 10616 9456 10668
rect 11244 10616 11296 10668
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4988 10412 5040 10464
rect 7564 10480 7616 10532
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 7472 10412 7524 10464
rect 11888 10616 11940 10668
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 14280 10616 14332 10668
rect 14464 10616 14516 10668
rect 15752 10684 15804 10736
rect 19064 10752 19116 10804
rect 19432 10752 19484 10804
rect 20076 10752 20128 10804
rect 14924 10616 14976 10668
rect 15384 10616 15436 10668
rect 15844 10616 15896 10668
rect 16304 10616 16356 10668
rect 11520 10548 11572 10600
rect 12072 10591 12124 10600
rect 12072 10557 12081 10591
rect 12081 10557 12115 10591
rect 12115 10557 12124 10591
rect 12072 10548 12124 10557
rect 15200 10548 15252 10600
rect 16396 10548 16448 10600
rect 19340 10646 19392 10698
rect 19515 10659 19567 10668
rect 19515 10625 19531 10659
rect 19531 10625 19565 10659
rect 19565 10625 19567 10659
rect 19515 10616 19567 10625
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 20720 10616 20772 10668
rect 22376 10752 22428 10804
rect 22652 10752 22704 10804
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 19064 10548 19116 10600
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 19156 10455 19208 10464
rect 19156 10421 19165 10455
rect 19165 10421 19199 10455
rect 19199 10421 19208 10455
rect 19156 10412 19208 10421
rect 19340 10412 19392 10464
rect 22376 10412 22428 10464
rect 22744 10591 22796 10600
rect 22744 10557 22753 10591
rect 22753 10557 22787 10591
rect 22787 10557 22796 10591
rect 22744 10548 22796 10557
rect 3917 10310 3969 10362
rect 3981 10310 4033 10362
rect 4045 10310 4097 10362
rect 4109 10310 4161 10362
rect 4173 10310 4225 10362
rect 9851 10310 9903 10362
rect 9915 10310 9967 10362
rect 9979 10310 10031 10362
rect 10043 10310 10095 10362
rect 10107 10310 10159 10362
rect 15785 10310 15837 10362
rect 15849 10310 15901 10362
rect 15913 10310 15965 10362
rect 15977 10310 16029 10362
rect 16041 10310 16093 10362
rect 21719 10310 21771 10362
rect 21783 10310 21835 10362
rect 21847 10310 21899 10362
rect 21911 10310 21963 10362
rect 21975 10310 22027 10362
rect 2504 10208 2556 10260
rect 388 10072 440 10124
rect 2044 10072 2096 10124
rect 2412 10115 2464 10124
rect 2412 10081 2421 10115
rect 2421 10081 2455 10115
rect 2455 10081 2464 10115
rect 2412 10072 2464 10081
rect 3516 10072 3568 10124
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 2872 10004 2924 10056
rect 4344 10072 4396 10124
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 7380 10208 7432 10260
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 5540 10140 5592 10192
rect 4896 10072 4948 10124
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 5356 10072 5408 10124
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 5908 10072 5960 10081
rect 6368 10115 6420 10124
rect 6368 10081 6377 10115
rect 6377 10081 6411 10115
rect 6411 10081 6420 10115
rect 6368 10072 6420 10081
rect 6736 10115 6788 10124
rect 6736 10081 6770 10115
rect 6770 10081 6788 10115
rect 6736 10072 6788 10081
rect 11520 10208 11572 10260
rect 14004 10208 14056 10260
rect 17500 10208 17552 10260
rect 18328 10208 18380 10260
rect 18604 10208 18656 10260
rect 19156 10208 19208 10260
rect 19340 10208 19392 10260
rect 19616 10208 19668 10260
rect 20260 10208 20312 10260
rect 11704 10004 11756 10056
rect 12624 10004 12676 10056
rect 14004 10004 14056 10056
rect 10416 9936 10468 9988
rect 10968 9936 11020 9988
rect 5632 9911 5684 9920
rect 5632 9877 5641 9911
rect 5641 9877 5675 9911
rect 5675 9877 5684 9911
rect 5632 9868 5684 9877
rect 5816 9868 5868 9920
rect 8484 9868 8536 9920
rect 9588 9868 9640 9920
rect 11612 9868 11664 9920
rect 11980 9936 12032 9988
rect 12164 9936 12216 9988
rect 12348 9936 12400 9988
rect 12716 9868 12768 9920
rect 13728 9936 13780 9988
rect 19064 10140 19116 10192
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 15752 9936 15804 9988
rect 21180 10004 21232 10056
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 22744 10047 22796 10056
rect 22744 10013 22753 10047
rect 22753 10013 22787 10047
rect 22787 10013 22796 10047
rect 22744 10004 22796 10013
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23072 10047
rect 23020 10004 23072 10013
rect 21456 9936 21508 9988
rect 19892 9868 19944 9920
rect 20628 9868 20680 9920
rect 21180 9868 21232 9920
rect 21548 9868 21600 9920
rect 21824 9911 21876 9920
rect 21824 9877 21833 9911
rect 21833 9877 21867 9911
rect 21867 9877 21876 9911
rect 21824 9868 21876 9877
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 23756 9911 23808 9920
rect 23756 9877 23765 9911
rect 23765 9877 23799 9911
rect 23799 9877 23808 9911
rect 23756 9868 23808 9877
rect 6884 9766 6936 9818
rect 6948 9766 7000 9818
rect 7012 9766 7064 9818
rect 7076 9766 7128 9818
rect 7140 9766 7192 9818
rect 12818 9766 12870 9818
rect 12882 9766 12934 9818
rect 12946 9766 12998 9818
rect 13010 9766 13062 9818
rect 13074 9766 13126 9818
rect 18752 9766 18804 9818
rect 18816 9766 18868 9818
rect 18880 9766 18932 9818
rect 18944 9766 18996 9818
rect 19008 9766 19060 9818
rect 24686 9766 24738 9818
rect 24750 9766 24802 9818
rect 24814 9766 24866 9818
rect 24878 9766 24930 9818
rect 24942 9766 24994 9818
rect 1584 9664 1636 9716
rect 2412 9664 2464 9716
rect 2872 9664 2924 9716
rect 3332 9664 3384 9716
rect 4436 9664 4488 9716
rect 6368 9664 6420 9716
rect 2320 9596 2372 9648
rect 2504 9596 2556 9648
rect 3424 9596 3476 9648
rect 3516 9596 3568 9648
rect 3884 9596 3936 9648
rect 2044 9528 2096 9580
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 4344 9528 4396 9580
rect 5080 9528 5132 9580
rect 7564 9528 7616 9580
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4712 9460 4764 9512
rect 6552 9460 6604 9512
rect 10508 9664 10560 9716
rect 10692 9664 10744 9716
rect 11244 9707 11296 9716
rect 11244 9673 11253 9707
rect 11253 9673 11287 9707
rect 11287 9673 11296 9707
rect 11244 9664 11296 9673
rect 12624 9664 12676 9716
rect 14372 9664 14424 9716
rect 15200 9664 15252 9716
rect 15752 9664 15804 9716
rect 20996 9664 21048 9716
rect 21088 9707 21140 9716
rect 21088 9673 21097 9707
rect 21097 9673 21131 9707
rect 21131 9673 21140 9707
rect 21088 9664 21140 9673
rect 21548 9664 21600 9716
rect 21824 9664 21876 9716
rect 8116 9503 8168 9512
rect 8116 9469 8125 9503
rect 8125 9469 8159 9503
rect 8159 9469 8168 9503
rect 8116 9460 8168 9469
rect 8208 9460 8260 9512
rect 8668 9571 8720 9580
rect 8668 9537 8677 9571
rect 8677 9537 8711 9571
rect 8711 9537 8720 9571
rect 8668 9528 8720 9537
rect 11520 9596 11572 9648
rect 17316 9596 17368 9648
rect 18144 9596 18196 9648
rect 10416 9571 10468 9580
rect 10416 9537 10450 9571
rect 10450 9537 10468 9571
rect 10416 9528 10468 9537
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 9036 9460 9088 9512
rect 9680 9460 9732 9512
rect 10140 9460 10192 9512
rect 10784 9460 10836 9512
rect 10968 9460 11020 9512
rect 16948 9528 17000 9580
rect 18328 9571 18380 9580
rect 18328 9537 18337 9571
rect 18337 9537 18371 9571
rect 18371 9537 18380 9571
rect 18328 9528 18380 9537
rect 20628 9596 20680 9648
rect 22284 9664 22336 9716
rect 22836 9596 22888 9648
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 9128 9392 9180 9444
rect 4252 9324 4304 9376
rect 6000 9324 6052 9376
rect 10324 9324 10376 9376
rect 19708 9503 19760 9512
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 14004 9392 14056 9444
rect 18144 9392 18196 9444
rect 12164 9324 12216 9376
rect 15476 9324 15528 9376
rect 17132 9324 17184 9376
rect 17500 9324 17552 9376
rect 19524 9324 19576 9376
rect 22100 9324 22152 9376
rect 22192 9367 22244 9376
rect 22192 9333 22201 9367
rect 22201 9333 22235 9367
rect 22235 9333 22244 9367
rect 22192 9324 22244 9333
rect 22744 9503 22796 9512
rect 22744 9469 22753 9503
rect 22753 9469 22787 9503
rect 22787 9469 22796 9503
rect 22744 9460 22796 9469
rect 24216 9460 24268 9512
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 3917 9222 3969 9274
rect 3981 9222 4033 9274
rect 4045 9222 4097 9274
rect 4109 9222 4161 9274
rect 4173 9222 4225 9274
rect 9851 9222 9903 9274
rect 9915 9222 9967 9274
rect 9979 9222 10031 9274
rect 10043 9222 10095 9274
rect 10107 9222 10159 9274
rect 15785 9222 15837 9274
rect 15849 9222 15901 9274
rect 15913 9222 15965 9274
rect 15977 9222 16029 9274
rect 16041 9222 16093 9274
rect 21719 9222 21771 9274
rect 21783 9222 21835 9274
rect 21847 9222 21899 9274
rect 21911 9222 21963 9274
rect 21975 9222 22027 9274
rect 1308 9120 1360 9172
rect 3056 9120 3108 9172
rect 1676 9052 1728 9104
rect 2596 8984 2648 9036
rect 1676 8916 1728 8968
rect 2228 8916 2280 8968
rect 3792 9120 3844 9172
rect 7564 9120 7616 9172
rect 1216 8848 1268 8900
rect 664 8780 716 8832
rect 2596 8891 2648 8900
rect 2596 8857 2605 8891
rect 2605 8857 2639 8891
rect 2639 8857 2648 8891
rect 2596 8848 2648 8857
rect 3608 8916 3660 8968
rect 6368 8848 6420 8900
rect 7288 8848 7340 8900
rect 7380 8848 7432 8900
rect 7656 8848 7708 8900
rect 8668 9120 8720 9172
rect 9036 9120 9088 9172
rect 10600 9120 10652 9172
rect 13360 9052 13412 9104
rect 8484 8916 8536 8968
rect 10508 8984 10560 9036
rect 14004 9052 14056 9104
rect 22468 9120 22520 9172
rect 23388 9163 23440 9172
rect 23388 9129 23397 9163
rect 23397 9129 23431 9163
rect 23431 9129 23440 9163
rect 23388 9120 23440 9129
rect 24032 9120 24084 9172
rect 24124 9120 24176 9172
rect 22744 9052 22796 9104
rect 15476 9027 15528 9036
rect 15476 8993 15485 9027
rect 15485 8993 15519 9027
rect 15519 8993 15528 9027
rect 15476 8984 15528 8993
rect 9128 8916 9180 8968
rect 9312 8916 9364 8968
rect 10048 8959 10100 8968
rect 10048 8925 10055 8959
rect 10055 8925 10089 8959
rect 10089 8925 10100 8959
rect 10048 8916 10100 8925
rect 10232 8848 10284 8900
rect 11520 8848 11572 8900
rect 16304 8984 16356 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 14740 8780 14792 8832
rect 15108 8823 15160 8832
rect 15108 8789 15117 8823
rect 15117 8789 15151 8823
rect 15151 8789 15160 8823
rect 15108 8780 15160 8789
rect 15476 8780 15528 8832
rect 17592 8916 17644 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 22284 8916 22336 8968
rect 22376 8916 22428 8968
rect 23572 8916 23624 8968
rect 18604 8848 18656 8900
rect 21180 8848 21232 8900
rect 16120 8780 16172 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 17132 8780 17184 8832
rect 18144 8780 18196 8832
rect 20260 8780 20312 8832
rect 22836 8780 22888 8832
rect 6884 8678 6936 8730
rect 6948 8678 7000 8730
rect 7012 8678 7064 8730
rect 7076 8678 7128 8730
rect 7140 8678 7192 8730
rect 12818 8678 12870 8730
rect 12882 8678 12934 8730
rect 12946 8678 12998 8730
rect 13010 8678 13062 8730
rect 13074 8678 13126 8730
rect 18752 8678 18804 8730
rect 18816 8678 18868 8730
rect 18880 8678 18932 8730
rect 18944 8678 18996 8730
rect 19008 8678 19060 8730
rect 24686 8678 24738 8730
rect 24750 8678 24802 8730
rect 24814 8678 24866 8730
rect 24878 8678 24930 8730
rect 24942 8678 24994 8730
rect 1400 8576 1452 8628
rect 1952 8508 2004 8560
rect 8116 8576 8168 8628
rect 10324 8576 10376 8628
rect 6000 8508 6052 8560
rect 7748 8508 7800 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2872 8440 2924 8492
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7564 8440 7616 8492
rect 848 8372 900 8424
rect 1032 8304 1084 8356
rect 3332 8347 3384 8356
rect 3332 8313 3341 8347
rect 3341 8313 3375 8347
rect 3375 8313 3384 8347
rect 3332 8304 3384 8313
rect 6736 8372 6788 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 11612 8508 11664 8560
rect 11980 8551 12032 8560
rect 11980 8517 11989 8551
rect 11989 8517 12023 8551
rect 12023 8517 12032 8551
rect 11980 8508 12032 8517
rect 12256 8508 12308 8560
rect 12072 8483 12124 8492
rect 12072 8449 12081 8483
rect 12081 8449 12115 8483
rect 12115 8449 12124 8483
rect 12072 8440 12124 8449
rect 12624 8440 12676 8492
rect 13360 8576 13412 8628
rect 16672 8576 16724 8628
rect 13176 8508 13228 8560
rect 13636 8508 13688 8560
rect 13544 8440 13596 8492
rect 14004 8440 14056 8492
rect 14280 8440 14332 8492
rect 14924 8551 14976 8560
rect 14924 8517 14933 8551
rect 14933 8517 14967 8551
rect 14967 8517 14976 8551
rect 14924 8508 14976 8517
rect 15108 8508 15160 8560
rect 17316 8508 17368 8560
rect 22192 8576 22244 8628
rect 18144 8508 18196 8560
rect 23296 8576 23348 8628
rect 23756 8576 23808 8628
rect 17868 8483 17920 8492
rect 17868 8449 17877 8483
rect 17877 8449 17911 8483
rect 17911 8449 17920 8483
rect 17868 8440 17920 8449
rect 8576 8372 8628 8424
rect 11520 8372 11572 8424
rect 13820 8372 13872 8424
rect 8484 8304 8536 8356
rect 10048 8304 10100 8356
rect 10508 8304 10560 8356
rect 10876 8304 10928 8356
rect 15568 8372 15620 8424
rect 17684 8372 17736 8424
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 18788 8440 18840 8492
rect 19340 8440 19392 8492
rect 19524 8440 19576 8492
rect 20168 8483 20220 8492
rect 20168 8449 20177 8483
rect 20177 8449 20211 8483
rect 20211 8449 20220 8483
rect 20168 8440 20220 8449
rect 21548 8440 21600 8492
rect 22100 8440 22152 8492
rect 22468 8508 22520 8560
rect 22744 8508 22796 8560
rect 23020 8440 23072 8492
rect 24032 8483 24084 8492
rect 24032 8449 24041 8483
rect 24041 8449 24075 8483
rect 24075 8449 24084 8483
rect 24032 8440 24084 8449
rect 20628 8372 20680 8424
rect 22468 8372 22520 8424
rect 23572 8372 23624 8424
rect 480 8236 532 8288
rect 2412 8236 2464 8288
rect 2688 8236 2740 8288
rect 11704 8236 11756 8288
rect 18604 8236 18656 8288
rect 18696 8236 18748 8288
rect 19984 8236 20036 8288
rect 22744 8236 22796 8288
rect 24308 8279 24360 8288
rect 24308 8245 24317 8279
rect 24317 8245 24351 8279
rect 24351 8245 24360 8279
rect 24308 8236 24360 8245
rect 24676 8236 24728 8288
rect 3917 8134 3969 8186
rect 3981 8134 4033 8186
rect 4045 8134 4097 8186
rect 4109 8134 4161 8186
rect 4173 8134 4225 8186
rect 9851 8134 9903 8186
rect 9915 8134 9967 8186
rect 9979 8134 10031 8186
rect 10043 8134 10095 8186
rect 10107 8134 10159 8186
rect 15785 8134 15837 8186
rect 15849 8134 15901 8186
rect 15913 8134 15965 8186
rect 15977 8134 16029 8186
rect 16041 8134 16093 8186
rect 21719 8134 21771 8186
rect 21783 8134 21835 8186
rect 21847 8134 21899 8186
rect 21911 8134 21963 8186
rect 21975 8134 22027 8186
rect 1860 8032 1912 8084
rect 2044 8032 2096 8084
rect 2136 7828 2188 7880
rect 4712 7964 4764 8016
rect 3792 7896 3844 7948
rect 2044 7760 2096 7812
rect 2412 7760 2464 7812
rect 4160 7828 4212 7880
rect 4436 7896 4488 7948
rect 5356 8032 5408 8084
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6552 7896 6604 7948
rect 7196 8032 7248 8084
rect 7288 8032 7340 8084
rect 7380 7896 7432 7948
rect 11520 8032 11572 8084
rect 12072 8032 12124 8084
rect 12440 8032 12492 8084
rect 12624 8032 12676 8084
rect 13820 8032 13872 8084
rect 15384 7964 15436 8016
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 6368 7828 6420 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 2504 7692 2556 7744
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 5908 7760 5960 7812
rect 3884 7692 3936 7744
rect 10784 7896 10836 7948
rect 12164 7896 12216 7948
rect 13360 7896 13412 7948
rect 15844 7964 15896 8016
rect 16488 8032 16540 8084
rect 16856 8032 16908 8084
rect 15568 7896 15620 7948
rect 17132 7896 17184 7948
rect 18420 8032 18472 8084
rect 18696 8032 18748 8084
rect 17960 7964 18012 8016
rect 18604 7964 18656 8016
rect 20168 8032 20220 8084
rect 20996 8032 21048 8084
rect 22468 8032 22520 8084
rect 23020 8032 23072 8084
rect 20076 7964 20128 8016
rect 22744 7964 22796 8016
rect 10968 7760 11020 7812
rect 11888 7828 11940 7880
rect 11428 7760 11480 7812
rect 14740 7828 14792 7880
rect 15384 7828 15436 7880
rect 16212 7871 16264 7880
rect 16212 7837 16221 7871
rect 16221 7837 16255 7871
rect 16255 7837 16264 7871
rect 16212 7828 16264 7837
rect 17408 7828 17460 7880
rect 17316 7760 17368 7812
rect 18604 7828 18656 7880
rect 19524 7828 19576 7880
rect 19892 7828 19944 7880
rect 20352 7871 20404 7880
rect 20352 7837 20361 7871
rect 20361 7837 20395 7871
rect 20395 7837 20404 7871
rect 20352 7828 20404 7837
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 21088 7871 21140 7880
rect 21088 7837 21097 7871
rect 21097 7837 21131 7871
rect 21131 7837 21140 7871
rect 21088 7828 21140 7837
rect 22376 7828 22428 7880
rect 17592 7692 17644 7744
rect 17684 7692 17736 7744
rect 19340 7760 19392 7812
rect 19984 7760 20036 7812
rect 23664 7828 23716 7880
rect 20812 7692 20864 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 23940 7760 23992 7812
rect 6884 7590 6936 7642
rect 6948 7590 7000 7642
rect 7012 7590 7064 7642
rect 7076 7590 7128 7642
rect 7140 7590 7192 7642
rect 12818 7590 12870 7642
rect 12882 7590 12934 7642
rect 12946 7590 12998 7642
rect 13010 7590 13062 7642
rect 13074 7590 13126 7642
rect 18752 7590 18804 7642
rect 18816 7590 18868 7642
rect 18880 7590 18932 7642
rect 18944 7590 18996 7642
rect 19008 7590 19060 7642
rect 24686 7590 24738 7642
rect 24750 7590 24802 7642
rect 24814 7590 24866 7642
rect 24878 7590 24930 7642
rect 24942 7590 24994 7642
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 2596 7488 2648 7540
rect 4160 7488 4212 7540
rect 4896 7488 4948 7540
rect 5816 7488 5868 7540
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 388 7284 440 7336
rect 1860 7284 1912 7336
rect 2688 7284 2740 7336
rect 3424 7395 3476 7404
rect 3424 7361 3458 7395
rect 3458 7361 3476 7395
rect 3424 7352 3476 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 6736 7488 6788 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 9312 7488 9364 7540
rect 9680 7488 9732 7540
rect 9772 7488 9824 7540
rect 13360 7488 13412 7540
rect 8668 7352 8720 7404
rect 2964 7284 3016 7336
rect 4436 7284 4488 7336
rect 4528 7327 4580 7336
rect 4528 7293 4537 7327
rect 4537 7293 4571 7327
rect 4571 7293 4580 7327
rect 4528 7284 4580 7293
rect 4620 7284 4672 7336
rect 5080 7284 5132 7336
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 4988 7259 5040 7268
rect 4988 7225 4997 7259
rect 4997 7225 5031 7259
rect 5031 7225 5040 7259
rect 4988 7216 5040 7225
rect 6368 7148 6420 7200
rect 9220 7284 9272 7336
rect 9496 7420 9548 7472
rect 13176 7420 13228 7472
rect 14004 7488 14056 7540
rect 16672 7488 16724 7540
rect 14924 7420 14976 7472
rect 15844 7420 15896 7472
rect 18420 7488 18472 7540
rect 19892 7488 19944 7540
rect 20628 7488 20680 7540
rect 16948 7420 17000 7472
rect 17316 7420 17368 7472
rect 13912 7352 13964 7404
rect 14188 7352 14240 7404
rect 14372 7352 14424 7404
rect 19708 7420 19760 7472
rect 18788 7352 18840 7404
rect 13452 7284 13504 7336
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9496 7148 9548 7200
rect 9772 7148 9824 7200
rect 10324 7148 10376 7200
rect 20904 7352 20956 7404
rect 23572 7488 23624 7540
rect 23664 7488 23716 7540
rect 23940 7488 23992 7540
rect 22560 7425 22612 7472
rect 22560 7420 22585 7425
rect 22585 7420 22612 7425
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 21548 7284 21600 7336
rect 22100 7284 22152 7336
rect 24308 7420 24360 7472
rect 24400 7352 24452 7404
rect 25320 7284 25372 7336
rect 20812 7148 20864 7200
rect 21364 7148 21416 7200
rect 3917 7046 3969 7098
rect 3981 7046 4033 7098
rect 4045 7046 4097 7098
rect 4109 7046 4161 7098
rect 4173 7046 4225 7098
rect 9851 7046 9903 7098
rect 9915 7046 9967 7098
rect 9979 7046 10031 7098
rect 10043 7046 10095 7098
rect 10107 7046 10159 7098
rect 15785 7046 15837 7098
rect 15849 7046 15901 7098
rect 15913 7046 15965 7098
rect 15977 7046 16029 7098
rect 16041 7046 16093 7098
rect 21719 7046 21771 7098
rect 21783 7046 21835 7098
rect 21847 7046 21899 7098
rect 21911 7046 21963 7098
rect 21975 7046 22027 7098
rect 3608 6944 3660 6996
rect 1584 6808 1636 6860
rect 2044 6808 2096 6860
rect 4160 6876 4212 6928
rect 4896 6944 4948 6996
rect 5540 6987 5592 6996
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 5908 6944 5960 6996
rect 9036 6876 9088 6928
rect 10784 6876 10836 6928
rect 13452 6944 13504 6996
rect 17960 6944 18012 6996
rect 18604 6987 18656 6996
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 20352 6987 20404 6996
rect 20352 6953 20361 6987
rect 20361 6953 20395 6987
rect 20395 6953 20404 6987
rect 20352 6944 20404 6953
rect 20812 6944 20864 6996
rect 21088 6987 21140 6996
rect 21088 6953 21097 6987
rect 21097 6953 21131 6987
rect 21131 6953 21140 6987
rect 21088 6944 21140 6953
rect 21272 6987 21324 6996
rect 21272 6953 21281 6987
rect 21281 6953 21315 6987
rect 21315 6953 21324 6987
rect 21272 6944 21324 6953
rect 22192 6944 22244 6996
rect 22284 6944 22336 6996
rect 2228 6740 2280 6792
rect 2964 6740 3016 6792
rect 2596 6719 2621 6724
rect 2621 6719 2648 6724
rect 2596 6672 2648 6719
rect 3424 6672 3476 6724
rect 2044 6604 2096 6656
rect 3700 6604 3752 6656
rect 6736 6808 6788 6860
rect 7564 6808 7616 6860
rect 6184 6740 6236 6792
rect 9496 6808 9548 6860
rect 9864 6851 9916 6860
rect 9864 6817 9873 6851
rect 9873 6817 9907 6851
rect 9907 6817 9916 6851
rect 9864 6808 9916 6817
rect 10324 6808 10376 6860
rect 10048 6740 10100 6792
rect 8392 6672 8444 6724
rect 8944 6672 8996 6724
rect 15384 6808 15436 6860
rect 17868 6808 17920 6860
rect 20628 6876 20680 6928
rect 22744 6876 22796 6928
rect 12808 6783 12860 6792
rect 12808 6749 12815 6783
rect 12815 6749 12849 6783
rect 12849 6749 12860 6783
rect 12808 6740 12860 6749
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 13268 6672 13320 6724
rect 19340 6783 19392 6792
rect 19340 6749 19349 6783
rect 19349 6749 19383 6783
rect 19383 6749 19392 6783
rect 19340 6740 19392 6749
rect 19524 6740 19576 6792
rect 17684 6604 17736 6656
rect 18052 6604 18104 6656
rect 19156 6604 19208 6656
rect 19432 6604 19484 6656
rect 20536 6740 20588 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 21364 6740 21416 6792
rect 21456 6783 21508 6792
rect 21456 6749 21465 6783
rect 21465 6749 21499 6783
rect 21499 6749 21508 6783
rect 21456 6740 21508 6749
rect 21916 6740 21968 6792
rect 21088 6672 21140 6724
rect 20536 6604 20588 6656
rect 21272 6604 21324 6656
rect 21640 6604 21692 6656
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 23204 6740 23256 6792
rect 23388 6783 23440 6792
rect 23388 6749 23397 6783
rect 23397 6749 23431 6783
rect 23431 6749 23440 6783
rect 23388 6740 23440 6749
rect 22284 6672 22336 6724
rect 23572 6740 23624 6792
rect 22836 6604 22888 6656
rect 22928 6604 22980 6656
rect 23204 6647 23256 6656
rect 23204 6613 23213 6647
rect 23213 6613 23247 6647
rect 23247 6613 23256 6647
rect 23204 6604 23256 6613
rect 24032 6604 24084 6656
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 1308 6400 1360 6452
rect 3608 6400 3660 6452
rect 4712 6400 4764 6452
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5632 6400 5684 6452
rect 1216 6332 1268 6384
rect 2688 6332 2740 6384
rect 3240 6332 3292 6384
rect 2136 6264 2188 6316
rect 3792 6264 3844 6316
rect 4160 6264 4212 6316
rect 4344 6264 4396 6316
rect 1308 6128 1360 6180
rect 1400 6060 1452 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 6276 6264 6328 6316
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7380 6307 7432 6316
rect 7380 6273 7414 6307
rect 7414 6273 7432 6307
rect 7380 6264 7432 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 9496 6400 9548 6452
rect 9864 6400 9916 6452
rect 10048 6400 10100 6452
rect 10692 6400 10744 6452
rect 9772 6307 9824 6316
rect 9772 6273 9781 6307
rect 9781 6273 9815 6307
rect 9815 6273 9824 6307
rect 9772 6264 9824 6273
rect 9864 6307 9916 6316
rect 9864 6273 9898 6307
rect 9898 6273 9916 6307
rect 9864 6264 9916 6273
rect 11612 6264 11664 6316
rect 5908 6196 5960 6248
rect 6184 6196 6236 6248
rect 6828 6128 6880 6180
rect 7012 6171 7064 6180
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6920 6060 6972 6112
rect 8944 6196 8996 6248
rect 10232 6196 10284 6248
rect 10600 6196 10652 6248
rect 12440 6400 12492 6452
rect 13912 6400 13964 6452
rect 15568 6400 15620 6452
rect 16764 6400 16816 6452
rect 17868 6400 17920 6452
rect 21456 6400 21508 6452
rect 12532 6264 12584 6316
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 12716 6264 12768 6273
rect 11888 6196 11940 6248
rect 22192 6400 22244 6452
rect 22744 6400 22796 6452
rect 23388 6400 23440 6452
rect 24400 6400 24452 6452
rect 13360 6264 13412 6316
rect 15292 6264 15344 6316
rect 9404 6128 9456 6180
rect 9496 6171 9548 6180
rect 9496 6137 9505 6171
rect 9505 6137 9539 6171
rect 9539 6137 9548 6171
rect 9496 6128 9548 6137
rect 12164 6171 12216 6180
rect 12164 6137 12173 6171
rect 12173 6137 12207 6171
rect 12207 6137 12216 6171
rect 12164 6128 12216 6137
rect 13268 6128 13320 6180
rect 14740 6196 14792 6248
rect 10784 6060 10836 6112
rect 12440 6060 12492 6112
rect 12624 6060 12676 6112
rect 16212 6060 16264 6112
rect 18236 6264 18288 6316
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 20628 6264 20680 6316
rect 20904 6264 20956 6316
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21364 6264 21416 6316
rect 21456 6264 21508 6316
rect 18420 6196 18472 6248
rect 22468 6264 22520 6316
rect 22836 6264 22888 6316
rect 18144 6128 18196 6180
rect 21824 6239 21876 6248
rect 21824 6205 21833 6239
rect 21833 6205 21867 6239
rect 21867 6205 21876 6239
rect 21824 6196 21876 6205
rect 23756 6307 23808 6316
rect 23756 6273 23765 6307
rect 23765 6273 23799 6307
rect 23799 6273 23808 6307
rect 23756 6264 23808 6273
rect 25228 6332 25280 6384
rect 24492 6307 24544 6316
rect 24492 6273 24501 6307
rect 24501 6273 24535 6307
rect 24535 6273 24544 6307
rect 24492 6264 24544 6273
rect 17868 6060 17920 6112
rect 20904 6103 20956 6112
rect 20904 6069 20913 6103
rect 20913 6069 20947 6103
rect 20947 6069 20956 6103
rect 20904 6060 20956 6069
rect 21272 6060 21324 6112
rect 21640 6060 21692 6112
rect 23296 6060 23348 6112
rect 23572 6103 23624 6112
rect 23572 6069 23581 6103
rect 23581 6069 23615 6103
rect 23615 6069 23624 6103
rect 23572 6060 23624 6069
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 1768 5899 1820 5908
rect 1768 5865 1777 5899
rect 1777 5865 1811 5899
rect 1811 5865 1820 5899
rect 1768 5856 1820 5865
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 1032 5788 1084 5840
rect 3884 5856 3936 5908
rect 5356 5856 5408 5908
rect 3332 5788 3384 5840
rect 3700 5720 3752 5772
rect 2320 5695 2372 5704
rect 2320 5661 2329 5695
rect 2329 5661 2363 5695
rect 2363 5661 2372 5695
rect 2320 5652 2372 5661
rect 3884 5652 3936 5704
rect 4712 5788 4764 5840
rect 5908 5856 5960 5908
rect 4160 5652 4212 5704
rect 4252 5695 4304 5704
rect 4252 5661 4259 5695
rect 4259 5661 4293 5695
rect 4293 5661 4304 5695
rect 4252 5652 4304 5661
rect 6368 5856 6420 5908
rect 6552 5856 6604 5908
rect 7472 5856 7524 5908
rect 9496 5856 9548 5908
rect 10600 5856 10652 5908
rect 12164 5856 12216 5908
rect 12716 5856 12768 5908
rect 12440 5788 12492 5840
rect 15476 5788 15528 5840
rect 15568 5788 15620 5840
rect 6828 5720 6880 5772
rect 9220 5720 9272 5772
rect 5356 5584 5408 5636
rect 9588 5652 9640 5704
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 10048 5652 10100 5704
rect 10784 5652 10836 5704
rect 10968 5652 11020 5704
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 2872 5516 2924 5525
rect 4988 5559 5040 5568
rect 4988 5525 4997 5559
rect 4997 5525 5031 5559
rect 5031 5525 5040 5559
rect 4988 5516 5040 5525
rect 5724 5516 5776 5568
rect 6552 5516 6604 5568
rect 7012 5584 7064 5636
rect 7380 5584 7432 5636
rect 8392 5584 8444 5636
rect 8576 5584 8628 5636
rect 9404 5584 9456 5636
rect 11060 5584 11112 5636
rect 11520 5695 11572 5704
rect 11520 5661 11527 5695
rect 11527 5661 11561 5695
rect 11561 5661 11572 5695
rect 11520 5652 11572 5661
rect 12532 5652 12584 5704
rect 15384 5652 15436 5704
rect 16212 5856 16264 5908
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 16304 5763 16356 5772
rect 16304 5729 16338 5763
rect 16338 5729 16356 5763
rect 16304 5720 16356 5729
rect 17132 5720 17184 5772
rect 19524 5856 19576 5908
rect 21088 5856 21140 5908
rect 21180 5899 21232 5908
rect 21180 5865 21189 5899
rect 21189 5865 21223 5899
rect 21223 5865 21232 5899
rect 21180 5856 21232 5865
rect 21364 5856 21416 5908
rect 23572 5856 23624 5908
rect 7656 5516 7708 5568
rect 13912 5584 13964 5636
rect 14924 5584 14976 5636
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 17500 5695 17552 5704
rect 17500 5661 17507 5695
rect 17507 5661 17541 5695
rect 17541 5661 17552 5695
rect 17500 5652 17552 5661
rect 20168 5720 20220 5772
rect 17684 5584 17736 5636
rect 17868 5584 17920 5636
rect 20352 5652 20404 5704
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 22376 5652 22428 5704
rect 22560 5652 22612 5704
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 23756 5652 23808 5704
rect 16580 5516 16632 5568
rect 19340 5516 19392 5568
rect 20904 5516 20956 5568
rect 21824 5627 21876 5636
rect 21824 5593 21858 5627
rect 21858 5593 21876 5627
rect 21824 5584 21876 5593
rect 22100 5584 22152 5636
rect 22652 5584 22704 5636
rect 23388 5584 23440 5636
rect 22192 5516 22244 5568
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 2136 5312 2188 5364
rect 2596 5312 2648 5364
rect 2688 5312 2740 5364
rect 3332 5312 3384 5364
rect 5264 5312 5316 5364
rect 5816 5312 5868 5364
rect 7380 5355 7432 5364
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 10232 5355 10284 5364
rect 10232 5321 10241 5355
rect 10241 5321 10275 5355
rect 10275 5321 10284 5355
rect 10232 5312 10284 5321
rect 10876 5312 10928 5364
rect 1308 5176 1360 5228
rect 2964 5176 3016 5228
rect 3056 5219 3108 5228
rect 3056 5185 3063 5219
rect 3063 5185 3097 5219
rect 3097 5185 3108 5219
rect 3056 5176 3108 5185
rect 4436 5176 4488 5228
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 5264 5219 5316 5228
rect 5264 5185 5273 5219
rect 5273 5185 5307 5219
rect 5307 5185 5316 5219
rect 5264 5176 5316 5185
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6736 5176 6788 5228
rect 10600 5244 10652 5296
rect 9864 5176 9916 5228
rect 10508 5176 10560 5228
rect 10876 5176 10928 5228
rect 4896 5108 4948 5160
rect 4988 5151 5040 5160
rect 4988 5117 4997 5151
rect 4997 5117 5031 5151
rect 5031 5117 5040 5151
rect 4988 5108 5040 5117
rect 5080 5108 5132 5160
rect 8944 5108 8996 5160
rect 10968 5108 11020 5160
rect 2504 4972 2556 5024
rect 4068 5040 4120 5092
rect 4344 5040 4396 5092
rect 3608 4972 3660 5024
rect 6000 4972 6052 5024
rect 12348 5312 12400 5364
rect 13820 5312 13872 5364
rect 13912 5312 13964 5364
rect 17132 5312 17184 5364
rect 18144 5355 18196 5364
rect 18144 5321 18153 5355
rect 18153 5321 18187 5355
rect 18187 5321 18196 5355
rect 18144 5312 18196 5321
rect 18236 5312 18288 5364
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 19156 5312 19208 5364
rect 21916 5312 21968 5364
rect 13084 5176 13136 5228
rect 13360 5083 13412 5092
rect 13360 5049 13369 5083
rect 13369 5049 13403 5083
rect 13403 5049 13412 5083
rect 13360 5040 13412 5049
rect 12348 4972 12400 5024
rect 13820 5108 13872 5160
rect 13912 5151 13964 5160
rect 13912 5117 13921 5151
rect 13921 5117 13955 5151
rect 13955 5117 13964 5151
rect 13912 5108 13964 5117
rect 14924 5108 14976 5160
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 15384 5108 15436 5160
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 15752 5108 15804 5160
rect 16396 5108 16448 5160
rect 17592 5176 17644 5228
rect 17684 5176 17736 5228
rect 17776 5108 17828 5160
rect 15292 5083 15344 5092
rect 15292 5049 15301 5083
rect 15301 5049 15335 5083
rect 15335 5049 15344 5083
rect 15292 5040 15344 5049
rect 16304 5040 16356 5092
rect 17960 5040 18012 5092
rect 18788 5219 18840 5228
rect 18788 5185 18797 5219
rect 18797 5185 18831 5219
rect 18831 5185 18840 5219
rect 18788 5176 18840 5185
rect 19156 5219 19208 5228
rect 19156 5185 19165 5219
rect 19165 5185 19199 5219
rect 19199 5185 19208 5219
rect 19156 5176 19208 5185
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 19708 5244 19760 5296
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 21548 5219 21600 5228
rect 21548 5185 21557 5219
rect 21557 5185 21591 5219
rect 21591 5185 21600 5219
rect 21548 5176 21600 5185
rect 19616 5151 19668 5160
rect 19616 5117 19625 5151
rect 19625 5117 19659 5151
rect 19659 5117 19668 5151
rect 19616 5108 19668 5117
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 21456 5108 21508 5160
rect 21916 5176 21968 5228
rect 22008 5176 22060 5228
rect 22652 5219 22704 5228
rect 22652 5185 22661 5219
rect 22661 5185 22695 5219
rect 22695 5185 22704 5219
rect 22652 5176 22704 5185
rect 22928 5176 22980 5228
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 15752 4972 15804 5024
rect 20720 5040 20772 5092
rect 22560 5040 22612 5092
rect 19616 4972 19668 5024
rect 20076 4972 20128 5024
rect 21364 4972 21416 5024
rect 22376 5015 22428 5024
rect 22376 4981 22385 5015
rect 22385 4981 22419 5015
rect 22419 4981 22428 5015
rect 22376 4972 22428 4981
rect 22468 4972 22520 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 1492 4811 1544 4820
rect 1492 4777 1501 4811
rect 1501 4777 1535 4811
rect 1535 4777 1544 4811
rect 1492 4768 1544 4777
rect 2320 4768 2372 4820
rect 3792 4743 3844 4752
rect 3792 4709 3801 4743
rect 3801 4709 3835 4743
rect 3835 4709 3844 4743
rect 3792 4700 3844 4709
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 12348 4768 12400 4820
rect 13360 4768 13412 4820
rect 14556 4768 14608 4820
rect 16396 4811 16448 4820
rect 16396 4777 16405 4811
rect 16405 4777 16439 4811
rect 16439 4777 16448 4811
rect 16396 4768 16448 4777
rect 18788 4811 18840 4820
rect 18788 4777 18797 4811
rect 18797 4777 18831 4811
rect 18831 4777 18840 4811
rect 18788 4768 18840 4777
rect 19156 4768 19208 4820
rect 19616 4811 19668 4820
rect 19616 4777 19625 4811
rect 19625 4777 19659 4811
rect 19659 4777 19668 4811
rect 19616 4768 19668 4777
rect 20352 4811 20404 4820
rect 20352 4777 20361 4811
rect 20361 4777 20395 4811
rect 20395 4777 20404 4811
rect 20352 4768 20404 4777
rect 14372 4700 14424 4752
rect 2136 4632 2188 4684
rect 2412 4675 2464 4684
rect 2412 4641 2421 4675
rect 2421 4641 2455 4675
rect 2455 4641 2464 4675
rect 2412 4632 2464 4641
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 3516 4632 3568 4684
rect 4344 4632 4396 4684
rect 6368 4632 6420 4684
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 1860 4496 1912 4548
rect 3700 4428 3752 4480
rect 4344 4496 4396 4548
rect 4804 4607 4856 4616
rect 4804 4573 4811 4607
rect 4811 4573 4845 4607
rect 4845 4573 4856 4607
rect 4804 4564 4856 4573
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 12808 4564 12860 4616
rect 13544 4564 13596 4616
rect 6828 4496 6880 4548
rect 20720 4768 20772 4820
rect 21180 4768 21232 4820
rect 21548 4768 21600 4820
rect 22100 4768 22152 4820
rect 23204 4768 23256 4820
rect 25412 4768 25464 4820
rect 19340 4632 19392 4684
rect 14740 4564 14792 4616
rect 15568 4564 15620 4616
rect 16120 4564 16172 4616
rect 16672 4564 16724 4616
rect 18604 4564 18656 4616
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 17868 4496 17920 4548
rect 19800 4564 19852 4616
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20996 4632 21048 4684
rect 20536 4607 20588 4616
rect 20536 4573 20545 4607
rect 20545 4573 20579 4607
rect 20579 4573 20588 4607
rect 20536 4564 20588 4573
rect 20628 4564 20680 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 8024 4428 8076 4480
rect 8668 4428 8720 4480
rect 9128 4428 9180 4480
rect 10416 4428 10468 4480
rect 11888 4428 11940 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 20260 4471 20312 4480
rect 20260 4437 20269 4471
rect 20269 4437 20303 4471
rect 20303 4437 20312 4471
rect 20260 4428 20312 4437
rect 21640 4607 21692 4616
rect 21640 4573 21649 4607
rect 21649 4573 21683 4607
rect 21683 4573 21692 4607
rect 21640 4564 21692 4573
rect 21732 4471 21784 4480
rect 21732 4437 21741 4471
rect 21741 4437 21775 4471
rect 21775 4437 21784 4471
rect 21732 4428 21784 4437
rect 22284 4564 22336 4616
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22796 4607
rect 22744 4564 22796 4573
rect 25228 4564 25280 4616
rect 24216 4496 24268 4548
rect 22836 4428 22888 4480
rect 22928 4428 22980 4480
rect 23296 4428 23348 4480
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 4712 4224 4764 4276
rect 7748 4224 7800 4276
rect 8944 4224 8996 4276
rect 2136 4088 2188 4140
rect 1676 3995 1728 4004
rect 1676 3961 1685 3995
rect 1685 3961 1719 3995
rect 1719 3961 1728 3995
rect 1676 3952 1728 3961
rect 1860 3952 1912 4004
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3332 4131 3384 4140
rect 3332 4097 3341 4131
rect 3341 4097 3375 4131
rect 3375 4097 3384 4131
rect 3332 4088 3384 4097
rect 3516 4088 3568 4140
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 6184 4088 6236 4140
rect 6736 4131 6788 4140
rect 6736 4097 6745 4131
rect 6745 4097 6779 4131
rect 6779 4097 6788 4131
rect 6736 4088 6788 4097
rect 8484 4088 8536 4140
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 8116 4063 8168 4072
rect 8116 4029 8125 4063
rect 8125 4029 8159 4063
rect 8159 4029 8168 4063
rect 8116 4020 8168 4029
rect 8668 4020 8720 4072
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 2504 3884 2556 3936
rect 9680 4020 9732 4072
rect 10416 4156 10468 4208
rect 10600 4156 10652 4208
rect 10692 4088 10744 4140
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12716 4088 12768 4140
rect 15292 4224 15344 4276
rect 17684 4267 17736 4276
rect 17684 4233 17693 4267
rect 17693 4233 17727 4267
rect 17727 4233 17736 4267
rect 17684 4224 17736 4233
rect 15476 4156 15528 4208
rect 18512 4224 18564 4276
rect 18880 4224 18932 4276
rect 19248 4224 19300 4276
rect 20260 4224 20312 4276
rect 20536 4224 20588 4276
rect 21272 4224 21324 4276
rect 21640 4224 21692 4276
rect 22284 4224 22336 4276
rect 23204 4224 23256 4276
rect 14740 4088 14792 4140
rect 24584 4156 24636 4208
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18328 4088 18380 4140
rect 18696 4088 18748 4140
rect 18972 4088 19024 4140
rect 10048 4063 10100 4072
rect 10048 4029 10057 4063
rect 10057 4029 10091 4063
rect 10091 4029 10100 4063
rect 10048 4020 10100 4029
rect 9680 3884 9732 3936
rect 9956 3927 10008 3936
rect 9956 3893 9965 3927
rect 9965 3893 9999 3927
rect 9999 3893 10008 3927
rect 9956 3884 10008 3893
rect 10140 3884 10192 3936
rect 10324 3884 10376 3936
rect 12532 3927 12584 3936
rect 12532 3893 12541 3927
rect 12541 3893 12575 3927
rect 12575 3893 12584 3927
rect 12532 3884 12584 3893
rect 19432 4088 19484 4140
rect 20352 4131 20404 4140
rect 20352 4097 20386 4131
rect 20386 4097 20404 4131
rect 20352 4088 20404 4097
rect 22468 4088 22520 4140
rect 20076 4063 20128 4072
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 22100 4020 22152 4072
rect 22192 4020 22244 4072
rect 22744 4088 22796 4140
rect 23388 4088 23440 4140
rect 24032 4088 24084 4140
rect 18972 3952 19024 4004
rect 19156 3884 19208 3936
rect 19248 3884 19300 3936
rect 22652 3995 22704 4004
rect 22652 3961 22661 3995
rect 22661 3961 22695 3995
rect 22695 3961 22704 3995
rect 22652 3952 22704 3961
rect 24308 3952 24360 4004
rect 20444 3884 20496 3936
rect 20812 3884 20864 3936
rect 21456 3884 21508 3936
rect 22284 3884 22336 3936
rect 23940 3884 23992 3936
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 1768 3723 1820 3732
rect 1768 3689 1777 3723
rect 1777 3689 1811 3723
rect 1811 3689 1820 3723
rect 1768 3680 1820 3689
rect 2136 3680 2188 3732
rect 5356 3680 5408 3732
rect 1400 3612 1452 3664
rect 2780 3612 2832 3664
rect 5080 3612 5132 3664
rect 9404 3680 9456 3732
rect 9496 3680 9548 3732
rect 3700 3544 3752 3596
rect 20 3408 72 3460
rect 2228 3451 2280 3460
rect 2228 3417 2237 3451
rect 2237 3417 2271 3451
rect 2271 3417 2280 3451
rect 2228 3408 2280 3417
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 2780 3476 2832 3528
rect 4620 3476 4672 3528
rect 6736 3544 6788 3596
rect 9680 3612 9732 3664
rect 7288 3476 7340 3528
rect 9956 3587 10008 3596
rect 9956 3553 9990 3587
rect 9990 3553 10008 3587
rect 9956 3544 10008 3553
rect 2044 3340 2096 3392
rect 2596 3340 2648 3392
rect 4528 3340 4580 3392
rect 4896 3383 4948 3392
rect 4896 3349 4905 3383
rect 4905 3349 4939 3383
rect 4939 3349 4948 3383
rect 4896 3340 4948 3349
rect 6000 3408 6052 3460
rect 7656 3476 7708 3528
rect 7840 3476 7892 3528
rect 8116 3476 8168 3528
rect 9036 3476 9088 3528
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 8208 3408 8260 3460
rect 5908 3340 5960 3392
rect 6092 3383 6144 3392
rect 6092 3349 6101 3383
rect 6101 3349 6135 3383
rect 6135 3349 6144 3383
rect 6092 3340 6144 3349
rect 7288 3340 7340 3392
rect 13360 3723 13412 3732
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 13912 3680 13964 3732
rect 17592 3680 17644 3732
rect 18788 3680 18840 3732
rect 12532 3544 12584 3596
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 12256 3408 12308 3460
rect 12440 3451 12492 3460
rect 12440 3417 12449 3451
rect 12449 3417 12483 3451
rect 12483 3417 12492 3451
rect 12440 3408 12492 3417
rect 12532 3408 12584 3460
rect 12900 3408 12952 3460
rect 14372 3519 14424 3528
rect 14372 3485 14379 3519
rect 14379 3485 14413 3519
rect 14413 3485 14424 3519
rect 14372 3476 14424 3485
rect 18144 3544 18196 3596
rect 17960 3495 18012 3504
rect 17960 3461 17969 3495
rect 17969 3461 18003 3495
rect 18003 3461 18012 3495
rect 17960 3452 18012 3461
rect 19156 3612 19208 3664
rect 19984 3680 20036 3732
rect 20628 3723 20680 3732
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 23204 3680 23256 3732
rect 23112 3612 23164 3664
rect 20904 3544 20956 3596
rect 18788 3519 18840 3528
rect 18788 3485 18797 3519
rect 18797 3485 18831 3519
rect 18831 3485 18840 3519
rect 18788 3476 18840 3485
rect 19064 3519 19116 3528
rect 19064 3485 19073 3519
rect 19073 3485 19107 3519
rect 19107 3485 19116 3519
rect 19064 3476 19116 3485
rect 20720 3476 20772 3528
rect 21456 3476 21508 3528
rect 22284 3476 22336 3528
rect 23112 3476 23164 3528
rect 13544 3383 13596 3392
rect 13544 3349 13553 3383
rect 13553 3349 13587 3383
rect 13587 3349 13596 3383
rect 13544 3340 13596 3349
rect 17776 3383 17828 3392
rect 17776 3349 17785 3383
rect 17785 3349 17819 3383
rect 17819 3349 17828 3383
rect 17776 3340 17828 3349
rect 18052 3340 18104 3392
rect 19340 3408 19392 3460
rect 19524 3451 19576 3460
rect 19524 3417 19558 3451
rect 19558 3417 19576 3451
rect 19524 3408 19576 3417
rect 20996 3408 21048 3460
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 18696 3340 18748 3392
rect 19708 3340 19760 3392
rect 22100 3340 22152 3392
rect 24492 3408 24544 3460
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 2228 3136 2280 3188
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 4528 3179 4580 3188
rect 4528 3145 4537 3179
rect 4537 3145 4571 3179
rect 4571 3145 4580 3179
rect 4528 3136 4580 3145
rect 1032 3068 1084 3120
rect 2320 3068 2372 3120
rect 7288 3136 7340 3188
rect 7472 3136 7524 3188
rect 9312 3136 9364 3188
rect 11796 3136 11848 3188
rect 12072 3136 12124 3188
rect 12440 3136 12492 3188
rect 14372 3136 14424 3188
rect 17684 3136 17736 3188
rect 6552 3111 6604 3120
rect 6552 3077 6561 3111
rect 6561 3077 6595 3111
rect 6595 3077 6604 3111
rect 6552 3068 6604 3077
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3056 2932 3108 2984
rect 3332 3000 3384 3052
rect 7748 3068 7800 3120
rect 9588 3068 9640 3120
rect 10140 3068 10192 3120
rect 10324 3111 10376 3120
rect 10324 3077 10333 3111
rect 10333 3077 10367 3111
rect 10367 3077 10376 3111
rect 10324 3068 10376 3077
rect 10416 3068 10468 3120
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7012 3000 7064 3052
rect 4068 2932 4120 2984
rect 6092 2932 6144 2984
rect 7656 2932 7708 2984
rect 3424 2864 3476 2916
rect 3148 2796 3200 2848
rect 9312 3000 9364 3052
rect 10048 3000 10100 3052
rect 10508 3000 10560 3052
rect 11060 3111 11112 3120
rect 11060 3077 11069 3111
rect 11069 3077 11103 3111
rect 11103 3077 11112 3111
rect 11060 3068 11112 3077
rect 11520 3068 11572 3120
rect 10784 2932 10836 2984
rect 12164 3068 12216 3120
rect 16764 3068 16816 3120
rect 18328 3136 18380 3188
rect 19064 3136 19116 3188
rect 19524 3136 19576 3188
rect 20904 3136 20956 3188
rect 18972 3068 19024 3120
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 17868 3000 17920 3052
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 18880 3000 18932 3052
rect 20996 3068 21048 3120
rect 21364 3136 21416 3188
rect 19800 3000 19852 3052
rect 8944 2796 8996 2848
rect 9220 2796 9272 2848
rect 9956 2796 10008 2848
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 13820 2796 13872 2848
rect 17592 2932 17644 2984
rect 19616 2932 19668 2984
rect 19892 2932 19944 2984
rect 21180 3000 21232 3052
rect 23020 3000 23072 3052
rect 24032 3068 24084 3120
rect 23848 3000 23900 3052
rect 21548 2932 21600 2984
rect 17500 2796 17552 2848
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 18696 2864 18748 2916
rect 20720 2864 20772 2916
rect 20812 2864 20864 2916
rect 18972 2796 19024 2848
rect 19156 2796 19208 2848
rect 19984 2796 20036 2848
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 2136 2592 2188 2644
rect 1308 2456 1360 2508
rect 2964 2592 3016 2644
rect 5632 2592 5684 2644
rect 5816 2592 5868 2644
rect 6920 2592 6972 2644
rect 7288 2592 7340 2644
rect 7932 2592 7984 2644
rect 5080 2524 5132 2576
rect 8024 2524 8076 2576
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10784 2592 10836 2644
rect 11060 2524 11112 2576
rect 12256 2592 12308 2644
rect 12532 2524 12584 2576
rect 480 2320 532 2372
rect 2596 2388 2648 2440
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6736 2388 6788 2440
rect 7748 2456 7800 2508
rect 8576 2456 8628 2508
rect 7656 2431 7708 2440
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 7840 2388 7892 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 2688 2320 2740 2372
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 10692 2456 10744 2508
rect 11244 2456 11296 2508
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9496 2388 9548 2440
rect 9864 2431 9916 2440
rect 9864 2397 9873 2431
rect 9873 2397 9907 2431
rect 9907 2397 9916 2431
rect 9864 2388 9916 2397
rect 11152 2388 11204 2440
rect 14096 2456 14148 2508
rect 12072 2431 12124 2440
rect 12072 2397 12081 2431
rect 12081 2397 12115 2431
rect 12115 2397 12124 2431
rect 12072 2388 12124 2397
rect 12164 2388 12216 2440
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 15568 2388 15620 2440
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 16396 2431 16448 2440
rect 16396 2397 16405 2431
rect 16405 2397 16439 2431
rect 16439 2397 16448 2431
rect 16396 2388 16448 2397
rect 17040 2592 17092 2644
rect 17868 2592 17920 2644
rect 23480 2592 23532 2644
rect 23572 2592 23624 2644
rect 18880 2524 18932 2576
rect 19616 2524 19668 2576
rect 17316 2456 17368 2508
rect 17960 2456 18012 2508
rect 16948 2431 17000 2440
rect 16948 2397 16957 2431
rect 16957 2397 16991 2431
rect 16991 2397 17000 2431
rect 16948 2388 17000 2397
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 480 2184 532 2236
rect 5448 2252 5500 2304
rect 5816 2252 5868 2304
rect 6092 2252 6144 2304
rect 6276 2252 6328 2304
rect 7012 2252 7064 2304
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 7564 2252 7616 2304
rect 7840 2252 7892 2304
rect 8208 2252 8260 2304
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 8484 2252 8536 2304
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 9864 2252 9916 2304
rect 10416 2252 10468 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 11704 2252 11756 2304
rect 12164 2295 12216 2304
rect 12164 2261 12173 2295
rect 12173 2261 12207 2295
rect 12207 2261 12216 2295
rect 12164 2252 12216 2261
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 12532 2252 12584 2304
rect 13912 2252 13964 2304
rect 14464 2252 14516 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 17960 2320 18012 2372
rect 18420 2388 18472 2440
rect 18604 2388 18656 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19524 2431 19576 2440
rect 19524 2397 19533 2431
rect 19533 2397 19567 2431
rect 19567 2397 19576 2431
rect 19524 2388 19576 2397
rect 19800 2499 19852 2508
rect 19800 2465 19809 2499
rect 19809 2465 19843 2499
rect 19843 2465 19852 2499
rect 19800 2456 19852 2465
rect 22468 2456 22520 2508
rect 19892 2320 19944 2372
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 16212 2295 16264 2304
rect 16212 2261 16221 2295
rect 16221 2261 16255 2295
rect 16255 2261 16264 2295
rect 16212 2252 16264 2261
rect 16488 2295 16540 2304
rect 16488 2261 16497 2295
rect 16497 2261 16531 2295
rect 16531 2261 16540 2295
rect 16488 2252 16540 2261
rect 17500 2252 17552 2304
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 18420 2252 18472 2304
rect 19248 2295 19300 2304
rect 19248 2261 19257 2295
rect 19257 2261 19291 2295
rect 19291 2261 19300 2295
rect 19248 2252 19300 2261
rect 20720 2388 20772 2440
rect 20904 2388 20956 2440
rect 21548 2431 21600 2440
rect 21548 2397 21557 2431
rect 21557 2397 21591 2431
rect 21591 2397 21600 2431
rect 21548 2388 21600 2397
rect 21824 2388 21876 2440
rect 22652 2388 22704 2440
rect 21548 2252 21600 2304
rect 23480 2252 23532 2304
rect 25596 2252 25648 2304
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 848 2048 900 2100
rect 2412 2048 2464 2100
rect 1308 1912 1360 1964
rect 1400 1955 1452 1964
rect 1400 1921 1409 1955
rect 1409 1921 1443 1955
rect 1443 1921 1452 1955
rect 1400 1912 1452 1921
rect 4528 2091 4580 2100
rect 4528 2057 4537 2091
rect 4537 2057 4571 2091
rect 4571 2057 4580 2091
rect 4528 2048 4580 2057
rect 5448 2048 5500 2100
rect 2044 1912 2096 1964
rect 3240 1955 3292 1964
rect 3240 1921 3249 1955
rect 3249 1921 3283 1955
rect 3283 1921 3292 1955
rect 3240 1912 3292 1921
rect 3700 1955 3752 1964
rect 3700 1921 3709 1955
rect 3709 1921 3743 1955
rect 3743 1921 3752 1955
rect 3700 1912 3752 1921
rect 3792 1844 3844 1896
rect 4712 1912 4764 1964
rect 4804 1955 4856 1964
rect 4804 1921 4813 1955
rect 4813 1921 4847 1955
rect 4847 1921 4856 1955
rect 4804 1912 4856 1921
rect 4620 1844 4672 1896
rect 3056 1708 3108 1760
rect 6184 2023 6236 2032
rect 6184 1989 6193 2023
rect 6193 1989 6227 2023
rect 6227 1989 6236 2023
rect 6184 1980 6236 1989
rect 6552 2091 6604 2100
rect 6552 2057 6561 2091
rect 6561 2057 6595 2091
rect 6595 2057 6604 2091
rect 6552 2048 6604 2057
rect 5724 1912 5776 1964
rect 5908 1912 5960 1964
rect 7564 2048 7616 2100
rect 7748 2048 7800 2100
rect 7840 2048 7892 2100
rect 8116 2048 8168 2100
rect 8392 2091 8444 2100
rect 8392 2057 8401 2091
rect 8401 2057 8435 2091
rect 8435 2057 8444 2091
rect 8392 2048 8444 2057
rect 8484 2048 8536 2100
rect 8576 2048 8628 2100
rect 8852 2048 8904 2100
rect 10232 2048 10284 2100
rect 11612 2048 11664 2100
rect 5816 1844 5868 1896
rect 6460 1844 6512 1896
rect 5540 1708 5592 1760
rect 7288 1819 7340 1828
rect 7288 1785 7297 1819
rect 7297 1785 7331 1819
rect 7331 1785 7340 1819
rect 7288 1776 7340 1785
rect 8484 1912 8536 1964
rect 8668 2023 8720 2032
rect 8668 1989 8677 2023
rect 8677 1989 8711 2023
rect 8711 1989 8720 2023
rect 8668 1980 8720 1989
rect 9220 1985 9272 2032
rect 8944 1955 8996 1964
rect 8944 1921 8953 1955
rect 8953 1921 8987 1955
rect 8987 1921 8996 1955
rect 8944 1912 8996 1921
rect 9220 1980 9245 1985
rect 9245 1980 9272 1985
rect 9404 1980 9456 2032
rect 11704 1980 11756 2032
rect 12440 2048 12492 2100
rect 13544 2048 13596 2100
rect 11796 1955 11848 1964
rect 11796 1921 11805 1955
rect 11805 1921 11839 1955
rect 11839 1921 11848 1955
rect 11796 1912 11848 1921
rect 13544 1955 13596 1964
rect 13544 1921 13553 1955
rect 13553 1921 13587 1955
rect 13587 1921 13596 1955
rect 13544 1912 13596 1921
rect 14740 2048 14792 2100
rect 14924 2048 14976 2100
rect 15476 2048 15528 2100
rect 17960 2048 18012 2100
rect 19248 2048 19300 2100
rect 19524 2048 19576 2100
rect 9680 1844 9732 1896
rect 10508 1844 10560 1896
rect 15384 1955 15436 1964
rect 15384 1921 15393 1955
rect 15393 1921 15427 1955
rect 15427 1921 15436 1955
rect 15384 1912 15436 1921
rect 16764 2023 16816 2032
rect 16764 1989 16773 2023
rect 16773 1989 16807 2023
rect 16807 1989 16816 2023
rect 16764 1980 16816 1989
rect 17776 1980 17828 2032
rect 15016 1844 15068 1896
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 16304 1844 16356 1896
rect 19432 1844 19484 1896
rect 7656 1776 7708 1828
rect 8484 1776 8536 1828
rect 8852 1776 8904 1828
rect 14004 1776 14056 1828
rect 15384 1776 15436 1828
rect 6092 1708 6144 1760
rect 9864 1708 9916 1760
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 10968 1708 11020 1760
rect 11796 1708 11848 1760
rect 12072 1751 12124 1760
rect 12072 1717 12081 1751
rect 12081 1717 12115 1751
rect 12115 1717 12124 1751
rect 12072 1708 12124 1717
rect 12440 1751 12492 1760
rect 12440 1717 12449 1751
rect 12449 1717 12483 1751
rect 12483 1717 12492 1751
rect 12440 1708 12492 1717
rect 12624 1708 12676 1760
rect 13636 1751 13688 1760
rect 13636 1717 13645 1751
rect 13645 1717 13679 1751
rect 13679 1717 13688 1751
rect 13636 1708 13688 1717
rect 14096 1751 14148 1760
rect 14096 1717 14105 1751
rect 14105 1717 14139 1751
rect 14139 1717 14148 1751
rect 14096 1708 14148 1717
rect 14280 1708 14332 1760
rect 14740 1708 14792 1760
rect 15752 1751 15804 1760
rect 15752 1717 15761 1751
rect 15761 1717 15795 1751
rect 15795 1717 15804 1751
rect 15752 1708 15804 1717
rect 16856 1751 16908 1760
rect 16856 1717 16865 1751
rect 16865 1717 16899 1751
rect 16899 1717 16908 1751
rect 16856 1708 16908 1717
rect 17408 1751 17460 1760
rect 17408 1717 17417 1751
rect 17417 1717 17451 1751
rect 17451 1717 17460 1751
rect 17408 1708 17460 1717
rect 17592 1708 17644 1760
rect 19892 1912 19944 1964
rect 20904 1912 20956 1964
rect 21364 1980 21416 2032
rect 21548 1980 21600 2032
rect 22836 2048 22888 2100
rect 23020 1980 23072 2032
rect 25136 1980 25188 2032
rect 20076 1844 20128 1896
rect 21272 1844 21324 1896
rect 21548 1844 21600 1896
rect 21824 1887 21876 1896
rect 21824 1853 21833 1887
rect 21833 1853 21867 1887
rect 21867 1853 21876 1887
rect 21824 1844 21876 1853
rect 23664 1912 23716 1964
rect 20352 1708 20404 1760
rect 20628 1708 20680 1760
rect 23020 1708 23072 1760
rect 24860 1708 24912 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 3332 1504 3384 1556
rect 4896 1504 4948 1556
rect 7288 1504 7340 1556
rect 8668 1547 8720 1556
rect 8668 1513 8677 1547
rect 8677 1513 8711 1547
rect 8711 1513 8720 1547
rect 8668 1504 8720 1513
rect 8852 1504 8904 1556
rect 9496 1504 9548 1556
rect 13728 1504 13780 1556
rect 15108 1504 15160 1556
rect 756 1436 808 1488
rect 5816 1436 5868 1488
rect 6644 1436 6696 1488
rect 6736 1436 6788 1488
rect 11428 1436 11480 1488
rect 10048 1368 10100 1420
rect 11152 1368 11204 1420
rect 1400 1343 1452 1352
rect 1400 1309 1409 1343
rect 1409 1309 1443 1343
rect 1443 1309 1452 1343
rect 1400 1300 1452 1309
rect 1952 1343 2004 1352
rect 1952 1309 1961 1343
rect 1961 1309 1995 1343
rect 1995 1309 2004 1343
rect 1952 1300 2004 1309
rect 2044 1300 2096 1352
rect 1768 1275 1820 1284
rect 1768 1241 1777 1275
rect 1777 1241 1811 1275
rect 1811 1241 1820 1275
rect 1768 1232 1820 1241
rect 2320 1275 2372 1284
rect 2320 1241 2329 1275
rect 2329 1241 2363 1275
rect 2363 1241 2372 1275
rect 2320 1232 2372 1241
rect 3056 1343 3108 1352
rect 3056 1309 3065 1343
rect 3065 1309 3099 1343
rect 3099 1309 3108 1343
rect 3056 1300 3108 1309
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4068 1343 4120 1352
rect 4068 1309 4077 1343
rect 4077 1309 4111 1343
rect 4111 1309 4120 1343
rect 4068 1300 4120 1309
rect 5264 1343 5316 1352
rect 5264 1309 5273 1343
rect 5273 1309 5307 1343
rect 5307 1309 5316 1343
rect 5264 1300 5316 1309
rect 5540 1343 5592 1352
rect 5540 1309 5549 1343
rect 5549 1309 5583 1343
rect 5583 1309 5592 1343
rect 5540 1300 5592 1309
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 7472 1300 7524 1352
rect 7932 1343 7984 1352
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 8300 1300 8352 1352
rect 8392 1343 8444 1352
rect 8392 1309 8401 1343
rect 8401 1309 8435 1343
rect 8435 1309 8444 1343
rect 8392 1300 8444 1309
rect 2780 1207 2832 1216
rect 2780 1173 2789 1207
rect 2789 1173 2823 1207
rect 2823 1173 2832 1207
rect 2780 1164 2832 1173
rect 3424 1207 3476 1216
rect 3424 1173 3433 1207
rect 3433 1173 3467 1207
rect 3467 1173 3476 1207
rect 3424 1164 3476 1173
rect 4528 1232 4580 1284
rect 5632 1232 5684 1284
rect 6460 1232 6512 1284
rect 8852 1232 8904 1284
rect 3976 1164 4028 1216
rect 5172 1164 5224 1216
rect 6552 1207 6604 1216
rect 6552 1173 6561 1207
rect 6561 1173 6595 1207
rect 6595 1173 6604 1207
rect 6552 1164 6604 1173
rect 6736 1164 6788 1216
rect 7472 1207 7524 1216
rect 7472 1173 7481 1207
rect 7481 1173 7515 1207
rect 7515 1173 7524 1207
rect 7472 1164 7524 1173
rect 9680 1300 9732 1352
rect 9956 1300 10008 1352
rect 10416 1300 10468 1352
rect 14096 1436 14148 1488
rect 15200 1436 15252 1488
rect 16304 1547 16356 1556
rect 16304 1513 16313 1547
rect 16313 1513 16347 1547
rect 16347 1513 16356 1547
rect 16304 1504 16356 1513
rect 16672 1504 16724 1556
rect 16120 1436 16172 1488
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 12164 1300 12216 1352
rect 12440 1300 12492 1352
rect 9772 1164 9824 1216
rect 10324 1207 10376 1216
rect 10324 1173 10333 1207
rect 10333 1173 10367 1207
rect 10367 1173 10376 1207
rect 10324 1164 10376 1173
rect 10692 1164 10744 1216
rect 11244 1207 11296 1216
rect 11244 1173 11253 1207
rect 11253 1173 11287 1207
rect 11287 1173 11296 1207
rect 11244 1164 11296 1173
rect 12716 1232 12768 1284
rect 13636 1300 13688 1352
rect 13820 1343 13872 1352
rect 13820 1309 13829 1343
rect 13829 1309 13863 1343
rect 13863 1309 13872 1343
rect 13820 1300 13872 1309
rect 13912 1300 13964 1352
rect 14004 1300 14056 1352
rect 16396 1368 16448 1420
rect 17868 1436 17920 1488
rect 19432 1504 19484 1556
rect 20168 1504 20220 1556
rect 20536 1547 20588 1556
rect 20536 1513 20545 1547
rect 20545 1513 20579 1547
rect 20579 1513 20588 1547
rect 20536 1504 20588 1513
rect 22376 1504 22428 1556
rect 22468 1504 22520 1556
rect 22836 1504 22888 1556
rect 17684 1368 17736 1420
rect 21364 1368 21416 1420
rect 16488 1343 16540 1352
rect 16488 1309 16497 1343
rect 16497 1309 16531 1343
rect 16531 1309 16540 1343
rect 16488 1300 16540 1309
rect 16580 1300 16632 1352
rect 17500 1300 17552 1352
rect 18328 1300 18380 1352
rect 20536 1300 20588 1352
rect 22100 1436 22152 1488
rect 21640 1343 21692 1352
rect 21640 1309 21649 1343
rect 21649 1309 21683 1343
rect 21683 1309 21692 1343
rect 21640 1300 21692 1309
rect 25044 1368 25096 1420
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 12348 1164 12400 1173
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 14464 1232 14516 1284
rect 16212 1232 16264 1284
rect 20996 1232 21048 1284
rect 21180 1275 21232 1284
rect 21180 1241 21189 1275
rect 21189 1241 21223 1275
rect 21223 1241 21232 1275
rect 21180 1232 21232 1241
rect 21916 1275 21968 1284
rect 21916 1241 21925 1275
rect 21925 1241 21959 1275
rect 21959 1241 21968 1275
rect 21916 1232 21968 1241
rect 22100 1275 22152 1284
rect 22100 1241 22109 1275
rect 22109 1241 22143 1275
rect 22143 1241 22152 1275
rect 22100 1232 22152 1241
rect 22468 1343 22520 1352
rect 22468 1309 22477 1343
rect 22477 1309 22511 1343
rect 22511 1309 22520 1343
rect 22468 1300 22520 1309
rect 23756 1300 23808 1352
rect 22928 1232 22980 1284
rect 14004 1164 14056 1216
rect 21088 1164 21140 1216
rect 21272 1207 21324 1216
rect 21272 1173 21281 1207
rect 21281 1173 21315 1207
rect 21315 1173 21324 1207
rect 21272 1164 21324 1173
rect 22192 1164 22244 1216
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 572 960 624 1012
rect 2780 960 2832 1012
rect 3424 960 3476 1012
rect 6276 960 6328 1012
rect 9956 960 10008 1012
rect 12532 960 12584 1012
rect 21180 960 21232 1012
rect 25596 960 25648 1012
rect 9772 892 9824 944
rect 11060 892 11112 944
rect 12256 892 12308 944
rect 21088 892 21140 944
rect 24216 892 24268 944
rect 5172 824 5224 876
rect 21272 824 21324 876
rect 25504 824 25556 876
rect 7472 756 7524 808
rect 14188 756 14240 808
rect 22100 756 22152 808
rect 25228 756 25280 808
rect 1400 688 1452 740
rect 2412 688 2464 740
rect 10324 688 10376 740
rect 11336 688 11388 740
rect 20536 688 20588 740
rect 23204 688 23256 740
rect 11244 620 11296 672
rect 12072 620 12124 672
rect 20996 620 21048 672
rect 22008 620 22060 672
rect 21916 552 21968 604
rect 23756 552 23808 604
rect 18052 484 18104 536
rect 24216 484 24268 536
rect 21180 416 21232 468
rect 22468 416 22520 468
rect 8392 76 8444 128
rect 9404 76 9456 128
<< metal2 >>
rect 202 44463 258 44623
rect 478 44463 534 44623
rect 754 44463 810 44623
rect 1030 44463 1086 44623
rect 1306 44463 1362 44623
rect 1582 44463 1638 44623
rect 1858 44463 1914 44623
rect 2134 44463 2190 44623
rect 2410 44463 2466 44623
rect 2686 44463 2742 44623
rect 2962 44463 3018 44623
rect 3238 44463 3294 44623
rect 3514 44463 3570 44623
rect 3790 44463 3846 44623
rect 4066 44463 4122 44623
rect 4342 44463 4398 44623
rect 4618 44463 4674 44623
rect 4894 44463 4950 44623
rect 5170 44463 5226 44623
rect 5446 44463 5502 44623
rect 5722 44463 5778 44623
rect 5998 44463 6054 44623
rect 6274 44463 6330 44623
rect 6550 44463 6606 44623
rect 6826 44463 6882 44623
rect 7102 44463 7158 44623
rect 7378 44463 7434 44623
rect 7654 44463 7710 44623
rect 7930 44463 7986 44623
rect 8206 44463 8262 44623
rect 8482 44463 8538 44623
rect 8758 44463 8814 44623
rect 9034 44463 9090 44623
rect 9310 44463 9366 44623
rect 9586 44463 9642 44623
rect 9862 44463 9918 44623
rect 10138 44463 10194 44623
rect 10414 44463 10470 44623
rect 10690 44463 10746 44623
rect 10966 44463 11022 44623
rect 11242 44463 11298 44623
rect 11518 44463 11574 44623
rect 11794 44463 11850 44623
rect 12070 44463 12126 44623
rect 12346 44463 12402 44623
rect 12622 44463 12678 44623
rect 12898 44463 12954 44623
rect 13174 44463 13230 44623
rect 13450 44463 13506 44623
rect 13726 44463 13782 44623
rect 14002 44463 14058 44623
rect 14278 44463 14334 44623
rect 14554 44463 14610 44623
rect 14830 44463 14886 44623
rect 15106 44463 15162 44623
rect 15382 44463 15438 44623
rect 15658 44463 15714 44623
rect 15934 44463 15990 44623
rect 16210 44463 16266 44623
rect 16486 44463 16542 44623
rect 16762 44463 16818 44623
rect 17038 44463 17094 44623
rect 17314 44463 17370 44623
rect 17590 44463 17646 44623
rect 17866 44463 17922 44623
rect 18142 44463 18198 44623
rect 18418 44463 18474 44623
rect 18694 44463 18750 44623
rect 18970 44463 19026 44623
rect 19246 44463 19302 44623
rect 19522 44463 19578 44623
rect 19798 44463 19854 44623
rect 20074 44463 20130 44623
rect 20350 44463 20406 44623
rect 20626 44463 20682 44623
rect 20902 44463 20958 44623
rect 21178 44463 21234 44623
rect 21454 44463 21510 44623
rect 21730 44463 21786 44623
rect 22006 44463 22062 44623
rect 22282 44463 22338 44623
rect 22558 44463 22614 44623
rect 22834 44463 22890 44623
rect 23110 44463 23166 44623
rect 23386 44463 23442 44623
rect 23662 44463 23718 44623
rect 23938 44463 23994 44623
rect 24214 44463 24270 44623
rect 24490 44463 24546 44623
rect 24766 44463 24822 44623
rect 25042 44463 25098 44623
rect 25318 44463 25374 44623
rect 25594 44463 25650 44623
rect 216 43874 244 44463
rect 216 43846 428 43874
rect 400 43382 428 43846
rect 388 43376 440 43382
rect 388 43318 440 43324
rect 20 42696 72 42702
rect 20 42638 72 42644
rect 32 3466 60 42638
rect 492 42362 520 44463
rect 480 42356 532 42362
rect 480 42298 532 42304
rect 768 41800 796 44463
rect 1044 42004 1072 44463
rect 1216 43308 1268 43314
rect 1216 43250 1268 43256
rect 1228 42106 1256 43250
rect 1320 42752 1348 44463
rect 1400 42764 1452 42770
rect 1320 42724 1400 42752
rect 1400 42706 1452 42712
rect 1490 42120 1546 42129
rect 1228 42078 1348 42106
rect 1216 42016 1268 42022
rect 1044 41976 1216 42004
rect 1216 41958 1268 41964
rect 940 41812 992 41818
rect 768 41772 940 41800
rect 940 41754 992 41760
rect 480 41064 532 41070
rect 480 41006 532 41012
rect 388 40996 440 41002
rect 388 40938 440 40944
rect 294 36952 350 36961
rect 294 36887 350 36896
rect 204 29436 256 29442
rect 204 29378 256 29384
rect 216 22778 244 29378
rect 204 22772 256 22778
rect 204 22714 256 22720
rect 308 22094 336 36887
rect 400 24721 428 40938
rect 492 27674 520 41006
rect 1032 40928 1084 40934
rect 1032 40870 1084 40876
rect 938 40216 994 40225
rect 938 40151 994 40160
rect 662 40080 718 40089
rect 662 40015 718 40024
rect 676 31754 704 40015
rect 756 38276 808 38282
rect 756 38218 808 38224
rect 768 37913 796 38218
rect 754 37904 810 37913
rect 754 37839 810 37848
rect 756 35080 808 35086
rect 756 35022 808 35028
rect 768 34649 796 35022
rect 754 34640 810 34649
rect 754 34575 810 34584
rect 848 33992 900 33998
rect 848 33934 900 33940
rect 860 31890 888 33934
rect 848 31884 900 31890
rect 848 31826 900 31832
rect 584 31726 704 31754
rect 846 31784 902 31793
rect 584 29442 612 31726
rect 846 31719 902 31728
rect 572 29436 624 29442
rect 572 29378 624 29384
rect 570 29336 626 29345
rect 570 29271 626 29280
rect 664 29300 716 29306
rect 480 27668 532 27674
rect 480 27610 532 27616
rect 386 24712 442 24721
rect 386 24647 442 24656
rect 584 23458 612 29271
rect 664 29242 716 29248
rect 572 23452 624 23458
rect 572 23394 624 23400
rect 676 23338 704 29242
rect 756 28484 808 28490
rect 756 28426 808 28432
rect 768 28393 796 28426
rect 754 28384 810 28393
rect 754 28319 810 28328
rect 756 28076 808 28082
rect 756 28018 808 28024
rect 768 27849 796 28018
rect 754 27840 810 27849
rect 754 27775 810 27784
rect 756 24812 808 24818
rect 756 24754 808 24760
rect 768 23497 796 24754
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 492 23310 704 23338
rect 386 22264 442 22273
rect 386 22199 442 22208
rect 216 22066 336 22094
rect 216 19174 244 22066
rect 294 20088 350 20097
rect 294 20023 350 20032
rect 204 19168 256 19174
rect 204 19110 256 19116
rect 308 13258 336 20023
rect 296 13252 348 13258
rect 296 13194 348 13200
rect 400 12434 428 22199
rect 492 16658 520 23310
rect 572 23248 624 23254
rect 572 23190 624 23196
rect 664 23248 716 23254
rect 664 23190 716 23196
rect 480 16652 532 16658
rect 480 16594 532 16600
rect 308 12406 428 12434
rect 308 4298 336 12406
rect 480 11076 532 11082
rect 480 11018 532 11024
rect 388 10124 440 10130
rect 388 10066 440 10072
rect 400 7342 428 10066
rect 492 8294 520 11018
rect 480 8288 532 8294
rect 480 8230 532 8236
rect 388 7336 440 7342
rect 388 7278 440 7284
rect 386 4312 442 4321
rect 308 4270 386 4298
rect 386 4247 442 4256
rect 20 3460 72 3466
rect 20 3402 72 3408
rect 480 2372 532 2378
rect 400 2332 480 2360
rect 202 82 258 160
rect 400 82 428 2332
rect 480 2314 532 2320
rect 480 2236 532 2242
rect 480 2178 532 2184
rect 492 160 520 2178
rect 584 1018 612 23190
rect 676 18442 704 23190
rect 860 22094 888 31719
rect 952 30598 980 40151
rect 940 30592 992 30598
rect 940 30534 992 30540
rect 938 29744 994 29753
rect 938 29679 994 29688
rect 952 29238 980 29679
rect 940 29232 992 29238
rect 940 29174 992 29180
rect 1044 27962 1072 40870
rect 1216 38208 1268 38214
rect 1214 38176 1216 38185
rect 1268 38176 1270 38185
rect 1214 38111 1270 38120
rect 1124 37800 1176 37806
rect 1124 37742 1176 37748
rect 1136 33590 1164 37742
rect 1216 35624 1268 35630
rect 1216 35566 1268 35572
rect 1228 34406 1256 35566
rect 1216 34400 1268 34406
rect 1216 34342 1268 34348
rect 1216 33924 1268 33930
rect 1216 33866 1268 33872
rect 1124 33584 1176 33590
rect 1228 33561 1256 33866
rect 1124 33526 1176 33532
rect 1214 33552 1270 33561
rect 1214 33487 1270 33496
rect 1216 32768 1268 32774
rect 1216 32710 1268 32716
rect 1124 32564 1176 32570
rect 1124 32506 1176 32512
rect 1136 32201 1164 32506
rect 1228 32473 1256 32710
rect 1214 32464 1270 32473
rect 1214 32399 1270 32408
rect 1216 32224 1268 32230
rect 1122 32192 1178 32201
rect 1216 32166 1268 32172
rect 1122 32127 1178 32136
rect 1228 31929 1256 32166
rect 1214 31920 1270 31929
rect 1214 31855 1270 31864
rect 1320 31754 1348 42078
rect 1490 42055 1546 42064
rect 1504 41614 1532 42055
rect 1492 41608 1544 41614
rect 1492 41550 1544 41556
rect 1596 41478 1624 44463
rect 1872 43450 1900 44463
rect 2148 43602 2176 44463
rect 2148 43574 2268 43602
rect 1860 43444 1912 43450
rect 1860 43386 1912 43392
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1676 43104 1728 43110
rect 1676 43046 1728 43052
rect 1688 41546 1716 43046
rect 1780 42362 1808 43250
rect 2240 42906 2268 43574
rect 2424 43466 2452 44463
rect 2424 43438 2636 43466
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2228 42900 2280 42906
rect 2228 42842 2280 42848
rect 2320 42628 2372 42634
rect 2320 42570 2372 42576
rect 1768 42356 1820 42362
rect 1768 42298 1820 42304
rect 2332 41546 2360 42570
rect 2412 42220 2464 42226
rect 2412 42162 2464 42168
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 2320 41540 2372 41546
rect 2320 41482 2372 41488
rect 1584 41472 1636 41478
rect 1584 41414 1636 41420
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1412 40610 1440 41074
rect 1412 40582 1532 40610
rect 1400 40452 1452 40458
rect 1400 40394 1452 40400
rect 1412 39409 1440 40394
rect 1504 39545 1532 40582
rect 2228 40452 2280 40458
rect 2228 40394 2280 40400
rect 1584 40044 1636 40050
rect 1584 39986 1636 39992
rect 1490 39536 1546 39545
rect 1490 39471 1546 39480
rect 1398 39400 1454 39409
rect 1398 39335 1454 39344
rect 1492 39364 1544 39370
rect 1492 39306 1544 39312
rect 1504 39098 1532 39306
rect 1492 39092 1544 39098
rect 1492 39034 1544 39040
rect 1400 37868 1452 37874
rect 1400 37810 1452 37816
rect 1412 34921 1440 37810
rect 1492 37188 1544 37194
rect 1492 37130 1544 37136
rect 1398 34912 1454 34921
rect 1398 34847 1454 34856
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 1412 33998 1440 34478
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1400 33448 1452 33454
rect 1400 33390 1452 33396
rect 1412 33114 1440 33390
rect 1400 33108 1452 33114
rect 1400 33050 1452 33056
rect 1504 33017 1532 37130
rect 1596 35465 1624 39986
rect 1860 39976 1912 39982
rect 1860 39918 1912 39924
rect 1676 39364 1728 39370
rect 1676 39306 1728 39312
rect 1688 37913 1716 39306
rect 1872 38962 1900 39918
rect 2240 39409 2268 40394
rect 2320 39840 2372 39846
rect 2320 39782 2372 39788
rect 2226 39400 2282 39409
rect 2332 39370 2360 39782
rect 2226 39335 2282 39344
rect 2320 39364 2372 39370
rect 2320 39306 2372 39312
rect 1860 38956 1912 38962
rect 1860 38898 1912 38904
rect 1872 38350 1900 38898
rect 1860 38344 1912 38350
rect 1860 38286 1912 38292
rect 2226 38312 2282 38321
rect 1674 37904 1730 37913
rect 1674 37839 1730 37848
rect 1872 37806 1900 38286
rect 2226 38247 2228 38256
rect 2280 38247 2282 38256
rect 2228 38218 2280 38224
rect 2044 37936 2096 37942
rect 2096 37896 2176 37924
rect 2044 37878 2096 37884
rect 1860 37800 1912 37806
rect 1860 37742 1912 37748
rect 1676 37120 1728 37126
rect 1676 37062 1728 37068
rect 1688 36281 1716 37062
rect 1766 36680 1822 36689
rect 1766 36615 1768 36624
rect 1820 36615 1822 36624
rect 1768 36586 1820 36592
rect 1768 36372 1820 36378
rect 1768 36314 1820 36320
rect 1674 36272 1730 36281
rect 1674 36207 1730 36216
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1582 35456 1638 35465
rect 1582 35391 1638 35400
rect 1584 34604 1636 34610
rect 1688 34592 1716 36110
rect 1636 34564 1716 34592
rect 1584 34546 1636 34552
rect 1490 33008 1546 33017
rect 1490 32943 1546 32952
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1674 32872 1730 32881
rect 1228 31726 1348 31754
rect 1228 30682 1256 31726
rect 1308 31680 1360 31686
rect 1308 31622 1360 31628
rect 1320 31260 1348 31622
rect 1412 31385 1440 32846
rect 1674 32807 1676 32816
rect 1728 32807 1730 32816
rect 1676 32778 1728 32784
rect 1492 32360 1544 32366
rect 1492 32302 1544 32308
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1504 31929 1532 32302
rect 1490 31920 1546 31929
rect 1490 31855 1546 31864
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1400 31272 1452 31278
rect 1320 31232 1400 31260
rect 1400 31214 1452 31220
rect 1308 31136 1360 31142
rect 1308 31078 1360 31084
rect 1320 30841 1348 31078
rect 1306 30832 1362 30841
rect 1306 30767 1362 30776
rect 1228 30654 1348 30682
rect 1216 30592 1268 30598
rect 1216 30534 1268 30540
rect 952 27934 1072 27962
rect 952 24177 980 27934
rect 1228 27826 1256 30534
rect 1320 30326 1348 30654
rect 1308 30320 1360 30326
rect 1308 30262 1360 30268
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 29481 1348 29514
rect 1306 29472 1362 29481
rect 1306 29407 1362 29416
rect 1412 29458 1440 31214
rect 1596 30938 1624 32302
rect 1780 31482 1808 36314
rect 1872 34218 1900 37742
rect 1952 37324 2004 37330
rect 1952 37266 2004 37272
rect 1964 36553 1992 37266
rect 1950 36544 2006 36553
rect 1950 36479 2006 36488
rect 2044 36032 2096 36038
rect 2044 35974 2096 35980
rect 1952 35488 2004 35494
rect 1952 35430 2004 35436
rect 1964 35290 1992 35430
rect 1952 35284 2004 35290
rect 1952 35226 2004 35232
rect 2056 35086 2084 35974
rect 2148 35680 2176 37896
rect 2228 37188 2280 37194
rect 2228 37130 2280 37136
rect 2240 36145 2268 37130
rect 2320 36576 2372 36582
rect 2318 36544 2320 36553
rect 2372 36544 2374 36553
rect 2318 36479 2374 36488
rect 2226 36136 2282 36145
rect 2226 36071 2282 36080
rect 2148 35652 2268 35680
rect 2136 35556 2188 35562
rect 2136 35498 2188 35504
rect 2044 35080 2096 35086
rect 2044 35022 2096 35028
rect 2056 34649 2084 35022
rect 2148 34746 2176 35498
rect 2136 34740 2188 34746
rect 2136 34682 2188 34688
rect 2042 34640 2098 34649
rect 2042 34575 2044 34584
rect 2096 34575 2098 34584
rect 2044 34546 2096 34552
rect 2240 34474 2268 35652
rect 2332 35154 2360 36479
rect 2320 35148 2372 35154
rect 2320 35090 2372 35096
rect 2332 34610 2360 35090
rect 2320 34604 2372 34610
rect 2320 34546 2372 34552
rect 2228 34468 2280 34474
rect 2228 34410 2280 34416
rect 1872 34190 2084 34218
rect 1952 33652 2004 33658
rect 1952 33594 2004 33600
rect 1858 32464 1914 32473
rect 1858 32399 1914 32408
rect 1768 31476 1820 31482
rect 1768 31418 1820 31424
rect 1584 30932 1636 30938
rect 1584 30874 1636 30880
rect 1492 30660 1544 30666
rect 1492 30602 1544 30608
rect 1676 30660 1728 30666
rect 1676 30602 1728 30608
rect 1504 30161 1532 30602
rect 1688 30274 1716 30602
rect 1688 30246 1808 30274
rect 1584 30184 1636 30190
rect 1490 30152 1546 30161
rect 1584 30126 1636 30132
rect 1676 30184 1728 30190
rect 1676 30126 1728 30132
rect 1490 30087 1546 30096
rect 1596 29850 1624 30126
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1584 29640 1636 29646
rect 1584 29582 1636 29588
rect 1596 29481 1624 29582
rect 1688 29510 1716 30126
rect 1676 29504 1728 29510
rect 1582 29472 1638 29481
rect 1412 29430 1582 29458
rect 1044 27798 1256 27826
rect 1044 24970 1072 27798
rect 1412 27538 1440 29430
rect 1676 29446 1728 29452
rect 1582 29407 1638 29416
rect 1492 29164 1544 29170
rect 1492 29106 1544 29112
rect 1504 28801 1532 29106
rect 1490 28792 1546 28801
rect 1490 28727 1546 28736
rect 1584 28756 1636 28762
rect 1584 28698 1636 28704
rect 1596 28422 1624 28698
rect 1780 28642 1808 30246
rect 1872 28762 1900 32399
rect 1964 32042 1992 33594
rect 2056 32212 2084 34190
rect 2136 33856 2188 33862
rect 2136 33798 2188 33804
rect 2148 32366 2176 33798
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2136 32360 2188 32366
rect 2136 32302 2188 32308
rect 2056 32184 2176 32212
rect 1964 32014 2084 32042
rect 1952 31476 2004 31482
rect 1952 31418 2004 31424
rect 1964 29238 1992 31418
rect 2056 29646 2084 32014
rect 2148 30734 2176 32184
rect 2240 31754 2268 33458
rect 2332 32978 2360 34546
rect 2424 34202 2452 42162
rect 2516 41274 2544 43250
rect 2608 41818 2636 43438
rect 2700 42650 2728 44463
rect 2976 43450 3004 44463
rect 3252 43602 3280 44463
rect 3252 43574 3372 43602
rect 2964 43444 3016 43450
rect 2964 43386 3016 43392
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 3068 42673 3096 43250
rect 3344 42906 3372 43574
rect 3424 43376 3476 43382
rect 3424 43318 3476 43324
rect 3332 42900 3384 42906
rect 3332 42842 3384 42848
rect 3054 42664 3110 42673
rect 2700 42622 2820 42650
rect 2792 42566 2820 42622
rect 2872 42628 2924 42634
rect 3054 42599 3110 42608
rect 3240 42628 3292 42634
rect 2872 42570 2924 42576
rect 3240 42570 3292 42576
rect 2780 42560 2832 42566
rect 2780 42502 2832 42508
rect 2780 42220 2832 42226
rect 2780 42162 2832 42168
rect 2792 41818 2820 42162
rect 2596 41812 2648 41818
rect 2596 41754 2648 41760
rect 2780 41812 2832 41818
rect 2780 41754 2832 41760
rect 2884 41698 2912 42570
rect 3252 42362 3280 42570
rect 3240 42356 3292 42362
rect 3240 42298 3292 42304
rect 3436 42242 3464 43318
rect 3344 42214 3464 42242
rect 3148 42152 3200 42158
rect 3148 42094 3200 42100
rect 2792 41670 2912 41698
rect 2792 41274 2820 41670
rect 2964 41540 3016 41546
rect 2964 41482 3016 41488
rect 2976 41274 3004 41482
rect 3160 41414 3188 42094
rect 3344 41818 3372 42214
rect 3528 42090 3556 44463
rect 3608 43104 3660 43110
rect 3608 43046 3660 43052
rect 3620 42362 3648 43046
rect 3700 42764 3752 42770
rect 3700 42706 3752 42712
rect 3608 42356 3660 42362
rect 3608 42298 3660 42304
rect 3516 42084 3568 42090
rect 3516 42026 3568 42032
rect 3608 42084 3660 42090
rect 3608 42026 3660 42032
rect 3620 41818 3648 42026
rect 3332 41812 3384 41818
rect 3332 41754 3384 41760
rect 3608 41812 3660 41818
rect 3608 41754 3660 41760
rect 3712 41614 3740 42706
rect 3804 42362 3832 44463
rect 4080 43092 4108 44463
rect 4356 43450 4384 44463
rect 4344 43444 4396 43450
rect 4344 43386 4396 43392
rect 4436 43104 4488 43110
rect 4080 43064 4292 43092
rect 3917 43004 4225 43013
rect 3917 43002 3923 43004
rect 3979 43002 4003 43004
rect 4059 43002 4083 43004
rect 4139 43002 4163 43004
rect 4219 43002 4225 43004
rect 3979 42950 3981 43002
rect 4161 42950 4163 43002
rect 3917 42948 3923 42950
rect 3979 42948 4003 42950
rect 4059 42948 4083 42950
rect 4139 42948 4163 42950
rect 4219 42948 4225 42950
rect 3917 42939 4225 42948
rect 4264 42786 4292 43064
rect 4488 43064 4568 43092
rect 4436 43046 4488 43052
rect 4264 42770 4384 42786
rect 4264 42764 4396 42770
rect 4264 42758 4344 42764
rect 4344 42706 4396 42712
rect 4252 42696 4304 42702
rect 4252 42638 4304 42644
rect 3792 42356 3844 42362
rect 3792 42298 3844 42304
rect 3884 42220 3936 42226
rect 3804 42180 3884 42208
rect 3804 41682 3832 42180
rect 3884 42162 3936 42168
rect 3917 41916 4225 41925
rect 3917 41914 3923 41916
rect 3979 41914 4003 41916
rect 4059 41914 4083 41916
rect 4139 41914 4163 41916
rect 4219 41914 4225 41916
rect 3979 41862 3981 41914
rect 4161 41862 4163 41914
rect 3917 41860 3923 41862
rect 3979 41860 4003 41862
rect 4059 41860 4083 41862
rect 4139 41860 4163 41862
rect 4219 41860 4225 41862
rect 3917 41851 4225 41860
rect 4264 41818 4292 42638
rect 4436 42628 4488 42634
rect 4436 42570 4488 42576
rect 4448 41818 4476 42570
rect 4252 41812 4304 41818
rect 4252 41754 4304 41760
rect 4436 41812 4488 41818
rect 4436 41754 4488 41760
rect 3792 41676 3844 41682
rect 3792 41618 3844 41624
rect 3332 41608 3384 41614
rect 3332 41550 3384 41556
rect 3608 41608 3660 41614
rect 3608 41550 3660 41556
rect 3700 41608 3752 41614
rect 4252 41608 4304 41614
rect 3700 41550 3752 41556
rect 4158 41576 4214 41585
rect 3068 41386 3188 41414
rect 2504 41268 2556 41274
rect 2504 41210 2556 41216
rect 2780 41268 2832 41274
rect 2780 41210 2832 41216
rect 2964 41268 3016 41274
rect 2964 41210 3016 41216
rect 3068 40730 3096 41386
rect 3240 41132 3292 41138
rect 3240 41074 3292 41080
rect 3056 40724 3108 40730
rect 3056 40666 3108 40672
rect 3148 40656 3200 40662
rect 3148 40598 3200 40604
rect 2780 40452 2832 40458
rect 2780 40394 2832 40400
rect 2688 39500 2740 39506
rect 2688 39442 2740 39448
rect 2596 39364 2648 39370
rect 2596 39306 2648 39312
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 2516 36378 2544 36722
rect 2504 36372 2556 36378
rect 2504 36314 2556 36320
rect 2608 35680 2636 39306
rect 2700 38894 2728 39442
rect 2792 39001 2820 40394
rect 3160 40186 3188 40598
rect 3148 40180 3200 40186
rect 3148 40122 3200 40128
rect 3252 40089 3280 41074
rect 3344 40934 3372 41550
rect 3424 41540 3476 41546
rect 3424 41482 3476 41488
rect 3436 41449 3464 41482
rect 3422 41440 3478 41449
rect 3620 41414 3648 41550
rect 4252 41550 4304 41556
rect 4158 41511 4160 41520
rect 4212 41511 4214 41520
rect 4160 41482 4212 41488
rect 3620 41386 3740 41414
rect 3422 41375 3478 41384
rect 3424 41132 3476 41138
rect 3424 41074 3476 41080
rect 3332 40928 3384 40934
rect 3332 40870 3384 40876
rect 3332 40520 3384 40526
rect 3332 40462 3384 40468
rect 3238 40080 3294 40089
rect 3148 40044 3200 40050
rect 3238 40015 3294 40024
rect 3148 39986 3200 39992
rect 3056 39976 3108 39982
rect 3056 39918 3108 39924
rect 2872 39908 2924 39914
rect 2872 39850 2924 39856
rect 2778 38992 2834 39001
rect 2884 38962 2912 39850
rect 3068 39114 3096 39918
rect 2976 39086 3096 39114
rect 2778 38927 2834 38936
rect 2872 38956 2924 38962
rect 2872 38898 2924 38904
rect 2688 38888 2740 38894
rect 2688 38830 2740 38836
rect 2884 38282 2912 38898
rect 2872 38276 2924 38282
rect 2872 38218 2924 38224
rect 2976 37505 3004 39086
rect 3056 38956 3108 38962
rect 3056 38898 3108 38904
rect 3068 38457 3096 38898
rect 3054 38448 3110 38457
rect 3054 38383 3110 38392
rect 3056 38276 3108 38282
rect 3056 38218 3108 38224
rect 3068 38185 3096 38218
rect 3054 38176 3110 38185
rect 3054 38111 3110 38120
rect 2962 37496 3018 37505
rect 2962 37431 3018 37440
rect 2872 37256 2924 37262
rect 2778 37224 2834 37233
rect 2872 37198 2924 37204
rect 2778 37159 2780 37168
rect 2832 37159 2834 37168
rect 2780 37130 2832 37136
rect 2884 36258 2912 37198
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 2792 36230 2912 36258
rect 2688 36032 2740 36038
rect 2688 35974 2740 35980
rect 2700 35698 2728 35974
rect 2792 35737 2820 36230
rect 2872 36168 2924 36174
rect 2872 36110 2924 36116
rect 2778 35728 2834 35737
rect 2606 35652 2636 35680
rect 2688 35692 2740 35698
rect 2504 35624 2556 35630
rect 2504 35566 2556 35572
rect 2606 35578 2634 35652
rect 2778 35663 2834 35672
rect 2688 35634 2740 35640
rect 2516 35494 2544 35566
rect 2606 35550 2636 35578
rect 2504 35488 2556 35494
rect 2504 35430 2556 35436
rect 2504 34400 2556 34406
rect 2504 34342 2556 34348
rect 2412 34196 2464 34202
rect 2412 34138 2464 34144
rect 2320 32972 2372 32978
rect 2320 32914 2372 32920
rect 2516 32824 2544 34342
rect 2608 34134 2636 35550
rect 2884 34762 2912 36110
rect 2700 34734 2912 34762
rect 2596 34128 2648 34134
rect 2596 34070 2648 34076
rect 2608 33114 2636 34070
rect 2700 33969 2728 34734
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2792 34082 2820 34546
rect 2792 34054 2912 34082
rect 2976 34066 3004 37062
rect 3160 36825 3188 39986
rect 3240 39568 3292 39574
rect 3240 39510 3292 39516
rect 3146 36816 3202 36825
rect 3146 36751 3202 36760
rect 3148 36304 3200 36310
rect 3148 36246 3200 36252
rect 3056 36032 3108 36038
rect 3056 35974 3108 35980
rect 3068 35630 3096 35974
rect 3056 35624 3108 35630
rect 3056 35566 3108 35572
rect 3056 34196 3108 34202
rect 3056 34138 3108 34144
rect 2780 33992 2832 33998
rect 2686 33960 2742 33969
rect 2780 33934 2832 33940
rect 2686 33895 2742 33904
rect 2686 33824 2742 33833
rect 2686 33759 2742 33768
rect 2596 33108 2648 33114
rect 2596 33050 2648 33056
rect 2424 32796 2544 32824
rect 2424 32434 2452 32796
rect 2502 32600 2558 32609
rect 2502 32535 2558 32544
rect 2412 32428 2464 32434
rect 2412 32370 2464 32376
rect 2320 32360 2372 32366
rect 2320 32302 2372 32308
rect 2332 31754 2360 32302
rect 2424 31890 2452 32370
rect 2412 31884 2464 31890
rect 2412 31826 2464 31832
rect 2228 31748 2280 31754
rect 2332 31748 2464 31754
rect 2332 31726 2412 31748
rect 2228 31690 2280 31696
rect 2412 31690 2464 31696
rect 2228 31136 2280 31142
rect 2228 31078 2280 31084
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2240 30190 2268 31078
rect 2320 30932 2372 30938
rect 2320 30874 2372 30880
rect 2228 30184 2280 30190
rect 2134 30152 2190 30161
rect 2228 30126 2280 30132
rect 2134 30087 2190 30096
rect 2044 29640 2096 29646
rect 2044 29582 2096 29588
rect 1952 29232 2004 29238
rect 1952 29174 2004 29180
rect 2148 29102 2176 30087
rect 2228 29504 2280 29510
rect 2228 29446 2280 29452
rect 2136 29096 2188 29102
rect 2136 29038 2188 29044
rect 1952 29028 2004 29034
rect 1952 28970 2004 28976
rect 1860 28756 1912 28762
rect 1860 28698 1912 28704
rect 1964 28665 1992 28970
rect 1950 28656 2006 28665
rect 1780 28614 1900 28642
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1676 28484 1728 28490
rect 1676 28426 1728 28432
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1596 28098 1624 28358
rect 1688 28218 1716 28426
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 1504 28070 1624 28098
rect 1676 28076 1728 28082
rect 1400 27532 1452 27538
rect 1400 27474 1452 27480
rect 1216 27396 1268 27402
rect 1216 27338 1268 27344
rect 1228 26489 1256 27338
rect 1214 26480 1270 26489
rect 1412 26450 1440 27474
rect 1214 26415 1270 26424
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1122 26344 1178 26353
rect 1122 26279 1178 26288
rect 1136 25106 1164 26279
rect 1308 25968 1360 25974
rect 1308 25910 1360 25916
rect 1216 25696 1268 25702
rect 1216 25638 1268 25644
rect 1228 25265 1256 25638
rect 1320 25401 1348 25910
rect 1412 25906 1440 26386
rect 1400 25900 1452 25906
rect 1400 25842 1452 25848
rect 1306 25392 1362 25401
rect 1306 25327 1362 25336
rect 1400 25288 1452 25294
rect 1214 25256 1270 25265
rect 1400 25230 1452 25236
rect 1214 25191 1270 25200
rect 1136 25078 1256 25106
rect 1044 24954 1164 24970
rect 1044 24948 1176 24954
rect 1044 24942 1124 24948
rect 1124 24890 1176 24896
rect 1032 24880 1084 24886
rect 1032 24822 1084 24828
rect 938 24168 994 24177
rect 938 24103 994 24112
rect 1044 23769 1072 24822
rect 1124 24744 1176 24750
rect 1124 24686 1176 24692
rect 1136 24585 1164 24686
rect 1122 24576 1178 24585
rect 1122 24511 1178 24520
rect 1030 23760 1086 23769
rect 1030 23695 1086 23704
rect 1228 22094 1256 25078
rect 1308 24948 1360 24954
rect 1308 24890 1360 24896
rect 1320 23633 1348 24890
rect 1412 24041 1440 25230
rect 1504 24138 1532 28070
rect 1676 28018 1728 28024
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1596 26897 1624 27406
rect 1688 27130 1716 28018
rect 1780 27441 1808 28494
rect 1766 27432 1822 27441
rect 1766 27367 1822 27376
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1582 26888 1638 26897
rect 1582 26823 1638 26832
rect 1766 26888 1822 26897
rect 1766 26823 1822 26832
rect 1582 25800 1638 25809
rect 1582 25735 1638 25744
rect 1596 24954 1624 25735
rect 1676 25288 1728 25294
rect 1676 25230 1728 25236
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1584 24812 1636 24818
rect 1584 24754 1636 24760
rect 1492 24132 1544 24138
rect 1492 24074 1544 24080
rect 1398 24032 1454 24041
rect 1398 23967 1454 23976
rect 1400 23656 1452 23662
rect 1306 23624 1362 23633
rect 1400 23598 1452 23604
rect 1306 23559 1362 23568
rect 1412 23202 1440 23598
rect 1596 23225 1624 24754
rect 1688 24313 1716 25230
rect 1780 24834 1808 26823
rect 1872 25401 1900 28614
rect 2148 28626 2176 29038
rect 1950 28591 2006 28600
rect 2136 28620 2188 28626
rect 2136 28562 2188 28568
rect 2044 28552 2096 28558
rect 2044 28494 2096 28500
rect 1952 28416 2004 28422
rect 1952 28358 2004 28364
rect 1858 25392 1914 25401
rect 1858 25327 1914 25336
rect 1858 25256 1914 25265
rect 1858 25191 1914 25200
rect 1872 25158 1900 25191
rect 1860 25152 1912 25158
rect 1860 25094 1912 25100
rect 1964 24954 1992 28358
rect 2056 27713 2084 28494
rect 2042 27704 2098 27713
rect 2042 27639 2098 27648
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2056 26926 2084 27270
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 2042 26072 2098 26081
rect 2042 26007 2098 26016
rect 2056 25294 2084 26007
rect 2148 25378 2176 28562
rect 2240 27033 2268 29446
rect 2332 28393 2360 30874
rect 2410 30832 2466 30841
rect 2410 30767 2466 30776
rect 2424 30258 2452 30767
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2412 29708 2464 29714
rect 2412 29650 2464 29656
rect 2424 29510 2452 29650
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2318 28384 2374 28393
rect 2318 28319 2374 28328
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2332 27577 2360 28018
rect 2318 27568 2374 27577
rect 2318 27503 2374 27512
rect 2226 27024 2282 27033
rect 2226 26959 2282 26968
rect 2412 26988 2464 26994
rect 2240 25702 2268 26959
rect 2412 26930 2464 26936
rect 2424 26586 2452 26930
rect 2412 26580 2464 26586
rect 2412 26522 2464 26528
rect 2516 26330 2544 32535
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2608 32026 2636 32302
rect 2596 32020 2648 32026
rect 2596 31962 2648 31968
rect 2700 31822 2728 33759
rect 2792 32745 2820 33934
rect 2884 33289 2912 34054
rect 2964 34060 3016 34066
rect 2964 34002 3016 34008
rect 3068 33402 3096 34138
rect 3160 33590 3188 36246
rect 3252 35154 3280 39510
rect 3344 35834 3372 40462
rect 3436 40050 3464 41074
rect 3516 41064 3568 41070
rect 3516 41006 3568 41012
rect 3528 40594 3556 41006
rect 3516 40588 3568 40594
rect 3516 40530 3568 40536
rect 3516 40452 3568 40458
rect 3516 40394 3568 40400
rect 3528 40186 3556 40394
rect 3516 40180 3568 40186
rect 3516 40122 3568 40128
rect 3424 40044 3476 40050
rect 3424 39986 3476 39992
rect 3436 39930 3464 39986
rect 3436 39902 3556 39930
rect 3424 39840 3476 39846
rect 3424 39782 3476 39788
rect 3436 39642 3464 39782
rect 3424 39636 3476 39642
rect 3424 39578 3476 39584
rect 3424 38956 3476 38962
rect 3424 38898 3476 38904
rect 3436 38049 3464 38898
rect 3528 38894 3556 39902
rect 3608 39296 3660 39302
rect 3608 39238 3660 39244
rect 3516 38888 3568 38894
rect 3516 38830 3568 38836
rect 3620 38654 3648 39238
rect 3528 38626 3648 38654
rect 3422 38040 3478 38049
rect 3422 37975 3478 37984
rect 3528 37942 3556 38626
rect 3516 37936 3568 37942
rect 3516 37878 3568 37884
rect 3424 37120 3476 37126
rect 3424 37062 3476 37068
rect 3436 36310 3464 37062
rect 3528 36854 3556 37878
rect 3608 37868 3660 37874
rect 3608 37810 3660 37816
rect 3620 36854 3648 37810
rect 3516 36848 3568 36854
rect 3516 36790 3568 36796
rect 3608 36848 3660 36854
rect 3608 36790 3660 36796
rect 3424 36304 3476 36310
rect 3424 36246 3476 36252
rect 3332 35828 3384 35834
rect 3332 35770 3384 35776
rect 3424 35692 3476 35698
rect 3424 35634 3476 35640
rect 3240 35148 3292 35154
rect 3240 35090 3292 35096
rect 3252 33658 3280 35090
rect 3332 34468 3384 34474
rect 3332 34410 3384 34416
rect 3344 33930 3372 34410
rect 3436 34105 3464 35634
rect 3528 34950 3556 36790
rect 3608 36032 3660 36038
rect 3606 36000 3608 36009
rect 3660 36000 3662 36009
rect 3606 35935 3662 35944
rect 3608 35624 3660 35630
rect 3608 35566 3660 35572
rect 3516 34944 3568 34950
rect 3516 34886 3568 34892
rect 3422 34096 3478 34105
rect 3422 34031 3478 34040
rect 3332 33924 3384 33930
rect 3332 33866 3384 33872
rect 3240 33652 3292 33658
rect 3292 33612 3372 33640
rect 3240 33594 3292 33600
rect 3148 33584 3200 33590
rect 3148 33526 3200 33532
rect 2976 33374 3096 33402
rect 2870 33280 2926 33289
rect 2870 33215 2926 33224
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2976 32366 3004 33374
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 3148 32904 3200 32910
rect 3148 32846 3200 32852
rect 2964 32360 3016 32366
rect 2964 32302 3016 32308
rect 2964 31884 3016 31890
rect 3016 31844 3096 31872
rect 2964 31826 3016 31832
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 2780 31816 2832 31822
rect 2780 31758 2832 31764
rect 2792 31113 2820 31758
rect 2964 31680 3016 31686
rect 2964 31622 3016 31628
rect 2778 31104 2834 31113
rect 2778 31039 2834 31048
rect 2596 30728 2648 30734
rect 2594 30696 2596 30705
rect 2648 30696 2650 30705
rect 2594 30631 2650 30640
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2700 29850 2728 30194
rect 2688 29844 2740 29850
rect 2688 29786 2740 29792
rect 2780 29844 2832 29850
rect 2780 29786 2832 29792
rect 2596 29640 2648 29646
rect 2596 29582 2648 29588
rect 2608 28558 2636 29582
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2596 28552 2648 28558
rect 2594 28520 2596 28529
rect 2648 28520 2650 28529
rect 2594 28455 2650 28464
rect 2700 27577 2728 29446
rect 2792 28150 2820 29786
rect 2976 29782 3004 31622
rect 3068 30054 3096 31844
rect 3160 30433 3188 32846
rect 3146 30424 3202 30433
rect 3146 30359 3202 30368
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 2964 29776 3016 29782
rect 2964 29718 3016 29724
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2686 27568 2742 27577
rect 2686 27503 2742 27512
rect 2596 27056 2648 27062
rect 2596 26998 2648 27004
rect 2608 26625 2636 26998
rect 2594 26616 2650 26625
rect 2594 26551 2650 26560
rect 2332 26302 2544 26330
rect 2228 25696 2280 25702
rect 2228 25638 2280 25644
rect 2228 25492 2280 25498
rect 2332 25480 2360 26302
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2424 25752 2452 25978
rect 2424 25724 2544 25752
rect 2280 25452 2360 25480
rect 2228 25434 2280 25440
rect 2148 25350 2268 25378
rect 2044 25288 2096 25294
rect 2044 25230 2096 25236
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 1780 24806 1992 24834
rect 1768 24608 1820 24614
rect 1768 24550 1820 24556
rect 1674 24304 1730 24313
rect 1674 24239 1730 24248
rect 1780 23769 1808 24550
rect 1860 24132 1912 24138
rect 1860 24074 1912 24080
rect 1872 23866 1900 24074
rect 1860 23860 1912 23866
rect 1860 23802 1912 23808
rect 1766 23760 1822 23769
rect 1766 23695 1822 23704
rect 1582 23216 1638 23225
rect 1412 23174 1532 23202
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1308 23044 1360 23050
rect 1308 22986 1360 22992
rect 1320 22953 1348 22986
rect 1306 22944 1362 22953
rect 1306 22879 1362 22888
rect 1412 22574 1440 23054
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 860 22066 1072 22094
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 768 19854 796 20159
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 756 19848 808 19854
rect 756 19790 808 19796
rect 860 19378 888 19887
rect 848 19372 900 19378
rect 848 19314 900 19320
rect 940 18624 992 18630
rect 940 18566 992 18572
rect 676 18414 796 18442
rect 662 12608 718 12617
rect 662 12543 718 12552
rect 676 8838 704 12543
rect 664 8832 716 8838
rect 664 8774 716 8780
rect 768 7868 796 18414
rect 952 16674 980 18566
rect 1044 17105 1072 22066
rect 1136 22066 1256 22094
rect 1030 17096 1086 17105
rect 1030 17031 1086 17040
rect 1030 16960 1086 16969
rect 1030 16895 1086 16904
rect 1044 16794 1072 16895
rect 1032 16788 1084 16794
rect 1032 16730 1084 16736
rect 952 16646 1072 16674
rect 848 13252 900 13258
rect 848 13194 900 13200
rect 860 13138 888 13194
rect 860 13110 980 13138
rect 846 9344 902 9353
rect 846 9279 902 9288
rect 860 8430 888 9279
rect 848 8424 900 8430
rect 848 8366 900 8372
rect 676 7840 796 7868
rect 676 1476 704 7840
rect 848 2100 900 2106
rect 848 2042 900 2048
rect 756 1488 808 1494
rect 676 1448 756 1476
rect 756 1430 808 1436
rect 572 1012 624 1018
rect 572 954 624 960
rect 202 54 428 82
rect 202 0 258 54
rect 478 0 534 160
rect 754 82 810 160
rect 860 82 888 2042
rect 952 2009 980 13110
rect 1044 9353 1072 16646
rect 1030 9344 1086 9353
rect 1030 9279 1086 9288
rect 1030 9072 1086 9081
rect 1030 9007 1086 9016
rect 1044 8362 1072 9007
rect 1032 8356 1084 8362
rect 1032 8298 1084 8304
rect 1030 6624 1086 6633
rect 1030 6559 1086 6568
rect 1044 5846 1072 6559
rect 1032 5840 1084 5846
rect 1032 5782 1084 5788
rect 1032 3120 1084 3126
rect 1032 3062 1084 3068
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 1044 160 1072 3062
rect 1136 2281 1164 22066
rect 1216 21888 1268 21894
rect 1216 21830 1268 21836
rect 1306 21856 1362 21865
rect 1228 21593 1256 21830
rect 1306 21791 1362 21800
rect 1320 21690 1348 21791
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1214 21584 1270 21593
rect 1412 21554 1440 22510
rect 1504 22409 1532 23174
rect 1582 23151 1638 23160
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1490 22400 1546 22409
rect 1490 22335 1546 22344
rect 1688 21842 1716 22918
rect 1964 22710 1992 24806
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 2056 22094 2084 25230
rect 2148 24857 2176 25230
rect 2134 24848 2190 24857
rect 2134 24783 2190 24792
rect 2240 23662 2268 25350
rect 2320 25220 2372 25226
rect 2320 25162 2372 25168
rect 2332 24682 2360 25162
rect 2320 24676 2372 24682
rect 2320 24618 2372 24624
rect 2412 24268 2464 24274
rect 2412 24210 2464 24216
rect 2228 23656 2280 23662
rect 2228 23598 2280 23604
rect 2134 23488 2190 23497
rect 2134 23423 2190 23432
rect 1872 22066 2084 22094
rect 1766 21992 1822 22001
rect 1766 21927 1768 21936
rect 1820 21927 1822 21936
rect 1768 21898 1820 21904
rect 1596 21814 1716 21842
rect 1214 21519 1270 21528
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1308 21344 1360 21350
rect 1214 21312 1270 21321
rect 1308 21286 1360 21292
rect 1214 21247 1270 21256
rect 1228 21010 1256 21247
rect 1320 21049 1348 21286
rect 1412 21146 1440 21490
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 1306 21040 1362 21049
rect 1216 21004 1268 21010
rect 1306 20975 1362 20984
rect 1216 20946 1268 20952
rect 1400 20936 1452 20942
rect 1214 20904 1270 20913
rect 1400 20878 1452 20884
rect 1214 20839 1270 20848
rect 1308 20868 1360 20874
rect 1228 18630 1256 20839
rect 1308 20810 1360 20816
rect 1320 20777 1348 20810
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1412 20505 1440 20878
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1308 19780 1360 19786
rect 1308 19722 1360 19728
rect 1320 19689 1348 19722
rect 1306 19680 1362 19689
rect 1306 19615 1362 19624
rect 1412 18970 1440 20334
rect 1596 20058 1624 21814
rect 1674 21720 1730 21729
rect 1674 21655 1730 21664
rect 1688 21622 1716 21655
rect 1676 21616 1728 21622
rect 1676 21558 1728 21564
rect 1872 20913 1900 22066
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 1858 20904 1914 20913
rect 1858 20839 1914 20848
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1860 20256 1912 20262
rect 1860 20198 1912 20204
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1582 19816 1638 19825
rect 1582 19751 1638 19760
rect 1596 19514 1624 19751
rect 1584 19508 1636 19514
rect 1584 19450 1636 19456
rect 1766 19408 1822 19417
rect 1766 19343 1822 19352
rect 1676 19304 1728 19310
rect 1674 19272 1676 19281
rect 1728 19272 1730 19281
rect 1674 19207 1730 19216
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 1584 18828 1636 18834
rect 1308 18692 1360 18698
rect 1308 18634 1360 18640
rect 1216 18624 1268 18630
rect 1216 18566 1268 18572
rect 1216 18352 1268 18358
rect 1320 18329 1348 18634
rect 1216 18294 1268 18300
rect 1306 18320 1362 18329
rect 1228 18057 1256 18294
rect 1306 18255 1362 18264
rect 1214 18048 1270 18057
rect 1214 17983 1270 17992
rect 1412 17678 1440 18799
rect 1584 18770 1636 18776
rect 1490 18592 1546 18601
rect 1490 18527 1546 18536
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1504 17490 1532 18527
rect 1596 17864 1624 18770
rect 1688 18290 1716 19207
rect 1780 18290 1808 19343
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1596 17836 1716 17864
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1412 17462 1532 17490
rect 1412 16590 1440 17462
rect 1596 17354 1624 17711
rect 1504 17326 1624 17354
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1308 14816 1360 14822
rect 1308 14758 1360 14764
rect 1320 14414 1348 14758
rect 1308 14408 1360 14414
rect 1308 14350 1360 14356
rect 1216 13524 1268 13530
rect 1216 13466 1268 13472
rect 1228 13161 1256 13466
rect 1214 13152 1270 13161
rect 1214 13087 1270 13096
rect 1320 12306 1348 14350
rect 1400 14068 1452 14074
rect 1504 14056 1532 17326
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1452 14028 1532 14056
rect 1400 14010 1452 14016
rect 1398 13968 1454 13977
rect 1398 13903 1454 13912
rect 1412 12434 1440 13903
rect 1596 13258 1624 16934
rect 1688 15994 1716 17836
rect 1766 17504 1822 17513
rect 1766 17439 1822 17448
rect 1780 16250 1808 17439
rect 1872 17134 1900 20198
rect 1964 19417 1992 20742
rect 2056 20505 2084 21898
rect 2148 21457 2176 23423
rect 2240 22642 2268 23598
rect 2424 23322 2452 24210
rect 2516 24206 2544 25724
rect 2596 25696 2648 25702
rect 2596 25638 2648 25644
rect 2504 24200 2556 24206
rect 2608 24188 2636 25638
rect 2700 24256 2728 27503
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2792 26897 2820 27066
rect 2778 26888 2834 26897
rect 2778 26823 2834 26832
rect 2884 26466 2912 29106
rect 2964 28076 3016 28082
rect 2964 28018 3016 28024
rect 2976 27441 3004 28018
rect 2962 27432 3018 27441
rect 2962 27367 3018 27376
rect 2964 27328 3016 27334
rect 2962 27296 2964 27305
rect 3016 27296 3018 27305
rect 2962 27231 3018 27240
rect 3068 27146 3096 29990
rect 3252 29850 3280 33050
rect 3344 32978 3372 33612
rect 3424 33516 3476 33522
rect 3424 33458 3476 33464
rect 3436 33114 3464 33458
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3332 32972 3384 32978
rect 3332 32914 3384 32920
rect 3424 32836 3476 32842
rect 3424 32778 3476 32784
rect 3436 32366 3464 32778
rect 3424 32360 3476 32366
rect 3424 32302 3476 32308
rect 3332 31272 3384 31278
rect 3332 31214 3384 31220
rect 3344 30938 3372 31214
rect 3332 30932 3384 30938
rect 3332 30874 3384 30880
rect 3424 30252 3476 30258
rect 3344 30212 3424 30240
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3148 29572 3200 29578
rect 3148 29514 3200 29520
rect 3160 28121 3188 29514
rect 3240 29504 3292 29510
rect 3240 29446 3292 29452
rect 3252 29345 3280 29446
rect 3238 29336 3294 29345
rect 3238 29271 3294 29280
rect 3344 29209 3372 30212
rect 3424 30194 3476 30200
rect 3330 29200 3386 29209
rect 3330 29135 3386 29144
rect 3240 29028 3292 29034
rect 3240 28970 3292 28976
rect 3146 28112 3202 28121
rect 3146 28047 3202 28056
rect 3252 28014 3280 28970
rect 3332 28416 3384 28422
rect 3332 28358 3384 28364
rect 3344 28150 3372 28358
rect 3528 28234 3556 34886
rect 3620 34406 3648 35566
rect 3608 34400 3660 34406
rect 3608 34342 3660 34348
rect 3606 34096 3662 34105
rect 3606 34031 3662 34040
rect 3620 29850 3648 34031
rect 3712 31482 3740 41386
rect 3917 40828 4225 40837
rect 3917 40826 3923 40828
rect 3979 40826 4003 40828
rect 4059 40826 4083 40828
rect 4139 40826 4163 40828
rect 4219 40826 4225 40828
rect 3979 40774 3981 40826
rect 4161 40774 4163 40826
rect 3917 40772 3923 40774
rect 3979 40772 4003 40774
rect 4059 40772 4083 40774
rect 4139 40772 4163 40774
rect 4219 40772 4225 40774
rect 3917 40763 4225 40772
rect 3792 40588 3844 40594
rect 3792 40530 3844 40536
rect 3804 40497 3832 40530
rect 3976 40520 4028 40526
rect 3790 40488 3846 40497
rect 3976 40462 4028 40468
rect 3790 40423 3846 40432
rect 3792 40384 3844 40390
rect 3792 40326 3844 40332
rect 3804 39506 3832 40326
rect 3988 39914 4016 40462
rect 4264 40225 4292 41550
rect 4540 41414 4568 43064
rect 4632 42566 4660 44463
rect 4804 43240 4856 43246
rect 4804 43182 4856 43188
rect 4712 43172 4764 43178
rect 4712 43114 4764 43120
rect 4724 42702 4752 43114
rect 4712 42696 4764 42702
rect 4712 42638 4764 42644
rect 4620 42560 4672 42566
rect 4620 42502 4672 42508
rect 4712 42220 4764 42226
rect 4712 42162 4764 42168
rect 4620 41608 4672 41614
rect 4618 41576 4620 41585
rect 4672 41576 4674 41585
rect 4618 41511 4674 41520
rect 4448 41386 4568 41414
rect 4250 40216 4306 40225
rect 4250 40151 4306 40160
rect 4344 39976 4396 39982
rect 4344 39918 4396 39924
rect 3976 39908 4028 39914
rect 3976 39850 4028 39856
rect 4252 39840 4304 39846
rect 4252 39782 4304 39788
rect 3917 39740 4225 39749
rect 3917 39738 3923 39740
rect 3979 39738 4003 39740
rect 4059 39738 4083 39740
rect 4139 39738 4163 39740
rect 4219 39738 4225 39740
rect 3979 39686 3981 39738
rect 4161 39686 4163 39738
rect 3917 39684 3923 39686
rect 3979 39684 4003 39686
rect 4059 39684 4083 39686
rect 4139 39684 4163 39686
rect 4219 39684 4225 39686
rect 3917 39675 4225 39684
rect 3792 39500 3844 39506
rect 4264 39488 4292 39782
rect 3792 39442 3844 39448
rect 4080 39460 4292 39488
rect 4080 39302 4108 39460
rect 4252 39364 4304 39370
rect 4252 39306 4304 39312
rect 4068 39296 4120 39302
rect 4068 39238 4120 39244
rect 4160 39296 4212 39302
rect 4160 39238 4212 39244
rect 4172 39098 4200 39238
rect 4160 39092 4212 39098
rect 4160 39034 4212 39040
rect 3884 38888 3936 38894
rect 3882 38856 3884 38865
rect 3936 38856 3938 38865
rect 3882 38791 3938 38800
rect 3917 38652 4225 38661
rect 3917 38650 3923 38652
rect 3979 38650 4003 38652
rect 4059 38650 4083 38652
rect 4139 38650 4163 38652
rect 4219 38650 4225 38652
rect 3979 38598 3981 38650
rect 4161 38598 4163 38650
rect 3917 38596 3923 38598
rect 3979 38596 4003 38598
rect 4059 38596 4083 38598
rect 4139 38596 4163 38598
rect 4219 38596 4225 38598
rect 3917 38587 4225 38596
rect 4264 37890 4292 39306
rect 4172 37874 4292 37890
rect 4160 37868 4292 37874
rect 4212 37862 4292 37868
rect 4160 37810 4212 37816
rect 3917 37564 4225 37573
rect 3917 37562 3923 37564
rect 3979 37562 4003 37564
rect 4059 37562 4083 37564
rect 4139 37562 4163 37564
rect 4219 37562 4225 37564
rect 3979 37510 3981 37562
rect 4161 37510 4163 37562
rect 3917 37508 3923 37510
rect 3979 37508 4003 37510
rect 4059 37508 4083 37510
rect 4139 37508 4163 37510
rect 4219 37508 4225 37510
rect 3917 37499 4225 37508
rect 3884 37460 3936 37466
rect 3884 37402 3936 37408
rect 3896 37097 3924 37402
rect 4068 37188 4120 37194
rect 4068 37130 4120 37136
rect 3882 37088 3938 37097
rect 3882 37023 3938 37032
rect 4080 36825 4108 37130
rect 4066 36816 4122 36825
rect 4066 36751 4122 36760
rect 3790 36544 3846 36553
rect 3790 36479 3846 36488
rect 3804 36310 3832 36479
rect 3917 36476 4225 36485
rect 3917 36474 3923 36476
rect 3979 36474 4003 36476
rect 4059 36474 4083 36476
rect 4139 36474 4163 36476
rect 4219 36474 4225 36476
rect 3979 36422 3981 36474
rect 4161 36422 4163 36474
rect 3917 36420 3923 36422
rect 3979 36420 4003 36422
rect 4059 36420 4083 36422
rect 4139 36420 4163 36422
rect 4219 36420 4225 36422
rect 3917 36411 4225 36420
rect 3792 36304 3844 36310
rect 3792 36246 3844 36252
rect 3792 36168 3844 36174
rect 3792 36110 3844 36116
rect 3804 35193 3832 36110
rect 4068 36100 4120 36106
rect 4068 36042 4120 36048
rect 4080 36009 4108 36042
rect 4066 36000 4122 36009
rect 4066 35935 4122 35944
rect 3917 35388 4225 35397
rect 3917 35386 3923 35388
rect 3979 35386 4003 35388
rect 4059 35386 4083 35388
rect 4139 35386 4163 35388
rect 4219 35386 4225 35388
rect 3979 35334 3981 35386
rect 4161 35334 4163 35386
rect 3917 35332 3923 35334
rect 3979 35332 4003 35334
rect 4059 35332 4083 35334
rect 4139 35332 4163 35334
rect 4219 35332 4225 35334
rect 3917 35323 4225 35332
rect 3790 35184 3846 35193
rect 3790 35119 3846 35128
rect 4264 35086 4292 37862
rect 4356 36961 4384 39918
rect 4342 36952 4398 36961
rect 4342 36887 4398 36896
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 4356 36242 4384 36722
rect 4344 36236 4396 36242
rect 4344 36178 4396 36184
rect 4252 35080 4304 35086
rect 4252 35022 4304 35028
rect 4344 35012 4396 35018
rect 4344 34954 4396 34960
rect 4250 34912 4306 34921
rect 4250 34847 4306 34856
rect 3884 34604 3936 34610
rect 3884 34546 3936 34552
rect 4160 34604 4212 34610
rect 4160 34546 4212 34552
rect 3896 34406 3924 34546
rect 4066 34504 4122 34513
rect 4172 34490 4200 34546
rect 4122 34462 4200 34490
rect 4066 34439 4122 34448
rect 3884 34400 3936 34406
rect 3884 34342 3936 34348
rect 3917 34300 4225 34309
rect 3917 34298 3923 34300
rect 3979 34298 4003 34300
rect 4059 34298 4083 34300
rect 4139 34298 4163 34300
rect 4219 34298 4225 34300
rect 3979 34246 3981 34298
rect 4161 34246 4163 34298
rect 3917 34244 3923 34246
rect 3979 34244 4003 34246
rect 4059 34244 4083 34246
rect 4139 34244 4163 34246
rect 4219 34244 4225 34246
rect 3917 34235 4225 34244
rect 3976 34128 4028 34134
rect 3976 34070 4028 34076
rect 3792 33652 3844 33658
rect 3792 33594 3844 33600
rect 3804 33114 3832 33594
rect 3988 33590 4016 34070
rect 3976 33584 4028 33590
rect 3976 33526 4028 33532
rect 3917 33212 4225 33221
rect 3917 33210 3923 33212
rect 3979 33210 4003 33212
rect 4059 33210 4083 33212
rect 4139 33210 4163 33212
rect 4219 33210 4225 33212
rect 3979 33158 3981 33210
rect 4161 33158 4163 33210
rect 3917 33156 3923 33158
rect 3979 33156 4003 33158
rect 4059 33156 4083 33158
rect 4139 33156 4163 33158
rect 4219 33156 4225 33158
rect 3917 33147 4225 33156
rect 3792 33108 3844 33114
rect 3792 33050 3844 33056
rect 4264 32366 4292 34847
rect 4356 34746 4384 34954
rect 4344 34740 4396 34746
rect 4344 34682 4396 34688
rect 4342 33688 4398 33697
rect 4342 33623 4398 33632
rect 4356 33454 4384 33623
rect 4344 33448 4396 33454
rect 4344 33390 4396 33396
rect 4344 32836 4396 32842
rect 4344 32778 4396 32784
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 4252 32360 4304 32366
rect 4252 32302 4304 32308
rect 3804 32008 3832 32302
rect 3917 32124 4225 32133
rect 3917 32122 3923 32124
rect 3979 32122 4003 32124
rect 4059 32122 4083 32124
rect 4139 32122 4163 32124
rect 4219 32122 4225 32124
rect 3979 32070 3981 32122
rect 4161 32070 4163 32122
rect 3917 32068 3923 32070
rect 3979 32068 4003 32070
rect 4059 32068 4083 32070
rect 4139 32068 4163 32070
rect 4219 32068 4225 32070
rect 3917 32059 4225 32068
rect 3804 31980 3924 32008
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3804 31657 3832 31758
rect 3790 31648 3846 31657
rect 3790 31583 3846 31592
rect 3896 31498 3924 31980
rect 4356 31754 4384 32778
rect 3700 31476 3752 31482
rect 3700 31418 3752 31424
rect 3804 31470 3924 31498
rect 4264 31726 4384 31754
rect 3804 30920 3832 31470
rect 3917 31036 4225 31045
rect 3917 31034 3923 31036
rect 3979 31034 4003 31036
rect 4059 31034 4083 31036
rect 4139 31034 4163 31036
rect 4219 31034 4225 31036
rect 3979 30982 3981 31034
rect 4161 30982 4163 31034
rect 3917 30980 3923 30982
rect 3979 30980 4003 30982
rect 4059 30980 4083 30982
rect 4139 30980 4163 30982
rect 4219 30980 4225 30982
rect 3917 30971 4225 30980
rect 3804 30892 4016 30920
rect 3792 30728 3844 30734
rect 3792 30670 3844 30676
rect 3698 30560 3754 30569
rect 3698 30495 3754 30504
rect 3712 30258 3740 30495
rect 3804 30297 3832 30670
rect 3882 30424 3938 30433
rect 3988 30394 4016 30892
rect 4160 30728 4212 30734
rect 4160 30670 4212 30676
rect 3882 30359 3938 30368
rect 3976 30388 4028 30394
rect 3790 30288 3846 30297
rect 3700 30252 3752 30258
rect 3896 30258 3924 30359
rect 3976 30330 4028 30336
rect 3790 30223 3846 30232
rect 3884 30252 3936 30258
rect 3700 30194 3752 30200
rect 3884 30194 3936 30200
rect 4172 30190 4200 30670
rect 4264 30598 4292 31726
rect 4448 31521 4476 41386
rect 4528 40928 4580 40934
rect 4528 40870 4580 40876
rect 4540 39438 4568 40870
rect 4528 39432 4580 39438
rect 4528 39374 4580 39380
rect 4528 39296 4580 39302
rect 4528 39238 4580 39244
rect 4540 37942 4568 39238
rect 4724 38729 4752 42162
rect 4816 39982 4844 43182
rect 4908 42770 4936 44463
rect 4896 42764 4948 42770
rect 4896 42706 4948 42712
rect 5184 42362 5212 44463
rect 5460 43874 5488 44463
rect 5460 43846 5580 43874
rect 5356 43648 5408 43654
rect 5356 43590 5408 43596
rect 5264 43308 5316 43314
rect 5264 43250 5316 43256
rect 5172 42356 5224 42362
rect 5172 42298 5224 42304
rect 5080 42084 5132 42090
rect 5080 42026 5132 42032
rect 5092 41682 5120 42026
rect 5276 41818 5304 43250
rect 5264 41812 5316 41818
rect 5264 41754 5316 41760
rect 4988 41676 5040 41682
rect 4988 41618 5040 41624
rect 5080 41676 5132 41682
rect 5080 41618 5132 41624
rect 4896 41064 4948 41070
rect 4896 41006 4948 41012
rect 4908 40594 4936 41006
rect 4896 40588 4948 40594
rect 4896 40530 4948 40536
rect 4908 39982 4936 40530
rect 5000 40440 5028 41618
rect 5264 41132 5316 41138
rect 5264 41074 5316 41080
rect 5276 40730 5304 41074
rect 5264 40724 5316 40730
rect 5264 40666 5316 40672
rect 5000 40412 5212 40440
rect 4804 39976 4856 39982
rect 4804 39918 4856 39924
rect 4896 39976 4948 39982
rect 4896 39918 4948 39924
rect 5080 39500 5132 39506
rect 5080 39442 5132 39448
rect 4896 39296 4948 39302
rect 4896 39238 4948 39244
rect 4908 39098 4936 39238
rect 4896 39092 4948 39098
rect 4896 39034 4948 39040
rect 4710 38720 4766 38729
rect 4710 38655 4766 38664
rect 4804 38208 4856 38214
rect 4804 38150 4856 38156
rect 4816 38010 4844 38150
rect 4804 38004 4856 38010
rect 4804 37946 4856 37952
rect 4528 37936 4580 37942
rect 4908 37890 4936 39034
rect 5092 38350 5120 39442
rect 5080 38344 5132 38350
rect 5080 38286 5132 38292
rect 4528 37878 4580 37884
rect 4540 36242 4568 37878
rect 4816 37874 4936 37890
rect 4804 37868 4936 37874
rect 4856 37862 4936 37868
rect 4988 37868 5040 37874
rect 4804 37810 4856 37816
rect 4988 37810 5040 37816
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 4632 36802 4660 37062
rect 4632 36786 4752 36802
rect 4632 36780 4764 36786
rect 4632 36774 4712 36780
rect 4712 36722 4764 36728
rect 4816 36718 4844 37810
rect 4896 37800 4948 37806
rect 4896 37742 4948 37748
rect 4908 37369 4936 37742
rect 5000 37466 5028 37810
rect 4988 37460 5040 37466
rect 4988 37402 5040 37408
rect 4894 37360 4950 37369
rect 4894 37295 4950 37304
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 4804 36712 4856 36718
rect 4856 36672 4936 36700
rect 4804 36654 4856 36660
rect 4620 36576 4672 36582
rect 4620 36518 4672 36524
rect 4804 36576 4856 36582
rect 4804 36518 4856 36524
rect 4632 36310 4660 36518
rect 4816 36310 4844 36518
rect 4620 36304 4672 36310
rect 4620 36246 4672 36252
rect 4804 36304 4856 36310
rect 4804 36246 4856 36252
rect 4528 36236 4580 36242
rect 4528 36178 4580 36184
rect 4712 36236 4764 36242
rect 4712 36178 4764 36184
rect 4528 35828 4580 35834
rect 4528 35770 4580 35776
rect 4540 35494 4568 35770
rect 4620 35624 4672 35630
rect 4620 35566 4672 35572
rect 4528 35488 4580 35494
rect 4528 35430 4580 35436
rect 4540 34626 4568 35430
rect 4632 34746 4660 35566
rect 4724 35018 4752 36178
rect 4804 36168 4856 36174
rect 4804 36110 4856 36116
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4540 34598 4752 34626
rect 4528 34536 4580 34542
rect 4528 34478 4580 34484
rect 4540 34066 4568 34478
rect 4620 34468 4672 34474
rect 4620 34410 4672 34416
rect 4528 34060 4580 34066
rect 4528 34002 4580 34008
rect 4540 33386 4568 34002
rect 4632 33590 4660 34410
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4528 33380 4580 33386
rect 4528 33322 4580 33328
rect 4632 32570 4660 33526
rect 4724 32774 4752 34598
rect 4712 32768 4764 32774
rect 4712 32710 4764 32716
rect 4620 32564 4672 32570
rect 4620 32506 4672 32512
rect 4620 32360 4672 32366
rect 4618 32328 4620 32337
rect 4672 32328 4674 32337
rect 4618 32263 4674 32272
rect 4724 32212 4752 32710
rect 4632 32184 4752 32212
rect 4434 31512 4490 31521
rect 4434 31447 4490 31456
rect 4344 31408 4396 31414
rect 4344 31350 4396 31356
rect 4436 31408 4488 31414
rect 4436 31350 4488 31356
rect 4528 31408 4580 31414
rect 4528 31350 4580 31356
rect 4356 30666 4384 31350
rect 4448 31249 4476 31350
rect 4434 31240 4490 31249
rect 4434 31175 4490 31184
rect 4540 31192 4568 31350
rect 4540 31164 4582 31192
rect 4554 30954 4582 31164
rect 4540 30938 4582 30954
rect 4528 30932 4582 30938
rect 4580 30926 4582 30932
rect 4528 30874 4580 30880
rect 4436 30728 4488 30734
rect 4436 30670 4488 30676
rect 4344 30660 4396 30666
rect 4344 30602 4396 30608
rect 4252 30592 4304 30598
rect 4448 30546 4476 30670
rect 4252 30534 4304 30540
rect 3792 30184 3844 30190
rect 3792 30126 3844 30132
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3804 29782 3832 30126
rect 3917 29948 4225 29957
rect 3917 29946 3923 29948
rect 3979 29946 4003 29948
rect 4059 29946 4083 29948
rect 4139 29946 4163 29948
rect 4219 29946 4225 29948
rect 3979 29894 3981 29946
rect 4161 29894 4163 29946
rect 3917 29892 3923 29894
rect 3979 29892 4003 29894
rect 4059 29892 4083 29894
rect 4139 29892 4163 29894
rect 4219 29892 4225 29894
rect 3917 29883 4225 29892
rect 3700 29776 3752 29782
rect 3700 29718 3752 29724
rect 3792 29776 3844 29782
rect 3792 29718 3844 29724
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3620 28937 3648 29106
rect 3606 28928 3662 28937
rect 3606 28863 3662 28872
rect 3712 28642 3740 29718
rect 3917 28860 4225 28869
rect 3917 28858 3923 28860
rect 3979 28858 4003 28860
rect 4059 28858 4083 28860
rect 4139 28858 4163 28860
rect 4219 28858 4225 28860
rect 3979 28806 3981 28858
rect 4161 28806 4163 28858
rect 3917 28804 3923 28806
rect 3979 28804 4003 28806
rect 4059 28804 4083 28806
rect 4139 28804 4163 28806
rect 4219 28804 4225 28806
rect 3917 28795 4225 28804
rect 3712 28614 3924 28642
rect 3792 28552 3844 28558
rect 3896 28540 3924 28614
rect 4160 28552 4212 28558
rect 3896 28520 4160 28540
rect 4212 28520 4214 28529
rect 3896 28512 4158 28520
rect 3792 28494 3844 28500
rect 3436 28206 3556 28234
rect 3332 28144 3384 28150
rect 3332 28086 3384 28092
rect 3240 28008 3292 28014
rect 3240 27950 3292 27956
rect 3332 27668 3384 27674
rect 3332 27610 3384 27616
rect 2964 27124 3016 27130
rect 3068 27118 3280 27146
rect 3344 27130 3372 27610
rect 2964 27066 3016 27072
rect 2792 26438 2912 26466
rect 2792 26081 2820 26438
rect 2872 26376 2924 26382
rect 2872 26318 2924 26324
rect 2778 26072 2834 26081
rect 2778 26007 2834 26016
rect 2780 25900 2832 25906
rect 2780 25842 2832 25848
rect 2792 25702 2820 25842
rect 2780 25696 2832 25702
rect 2884 25673 2912 26318
rect 2780 25638 2832 25644
rect 2870 25664 2926 25673
rect 2870 25599 2926 25608
rect 2870 24712 2926 24721
rect 2870 24647 2926 24656
rect 2780 24608 2832 24614
rect 2780 24550 2832 24556
rect 2792 24410 2820 24550
rect 2884 24410 2912 24647
rect 2780 24404 2832 24410
rect 2780 24346 2832 24352
rect 2872 24404 2924 24410
rect 2872 24346 2924 24352
rect 2700 24228 2912 24256
rect 2608 24160 2728 24188
rect 2504 24142 2556 24148
rect 2596 24064 2648 24070
rect 2596 24006 2648 24012
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2412 22432 2464 22438
rect 2412 22374 2464 22380
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 21690 2360 22034
rect 2424 22030 2452 22374
rect 2412 22024 2464 22030
rect 2412 21966 2464 21972
rect 2608 21690 2636 24006
rect 2700 22556 2728 24160
rect 2778 23896 2834 23905
rect 2778 23831 2834 23840
rect 2792 23730 2820 23831
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2792 23168 2820 23666
rect 2884 23322 2912 24228
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2872 23180 2924 23186
rect 2792 23140 2872 23168
rect 2872 23122 2924 23128
rect 2872 23044 2924 23050
rect 2872 22986 2924 22992
rect 2884 22681 2912 22986
rect 2870 22672 2926 22681
rect 2870 22607 2926 22616
rect 2700 22528 2912 22556
rect 2780 22432 2832 22438
rect 2780 22374 2832 22380
rect 2320 21684 2372 21690
rect 2320 21626 2372 21632
rect 2596 21684 2648 21690
rect 2596 21626 2648 21632
rect 2134 21448 2190 21457
rect 2134 21383 2190 21392
rect 2148 20942 2176 21383
rect 2594 21040 2650 21049
rect 2594 20975 2650 20984
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2318 20768 2374 20777
rect 2318 20703 2374 20712
rect 2042 20496 2098 20505
rect 2042 20431 2098 20440
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2044 19508 2096 19514
rect 2044 19450 2096 19456
rect 1950 19408 2006 19417
rect 1950 19343 2006 19352
rect 1964 18426 1992 19343
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1964 17134 1992 17546
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1872 16833 1900 17070
rect 1858 16824 1914 16833
rect 1858 16759 1914 16768
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1964 16028 1992 17070
rect 2056 16182 2084 19450
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 2148 16522 2176 18362
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 1964 16000 2084 16028
rect 1688 15966 1900 15994
rect 1674 15872 1730 15881
rect 1674 15807 1730 15816
rect 1688 13462 1716 15807
rect 1872 15026 1900 15966
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1780 14385 1808 14962
rect 1858 14648 1914 14657
rect 1858 14583 1914 14592
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1766 14240 1822 14249
rect 1766 14175 1822 14184
rect 1676 13456 1728 13462
rect 1676 13398 1728 13404
rect 1584 13252 1636 13258
rect 1584 13194 1636 13200
rect 1412 12406 1624 12434
rect 1308 12300 1360 12306
rect 1308 12242 1360 12248
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1214 9616 1270 9625
rect 1214 9551 1270 9560
rect 1228 8906 1256 9551
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1216 8900 1268 8906
rect 1216 8842 1268 8848
rect 1320 8537 1348 9114
rect 1412 8634 1440 11999
rect 1492 11008 1544 11014
rect 1492 10950 1544 10956
rect 1504 10742 1532 10950
rect 1596 10810 1624 12406
rect 1780 11354 1808 14175
rect 1872 12918 1900 14583
rect 1950 14240 2006 14249
rect 1950 14175 2006 14184
rect 1964 13938 1992 14175
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 1858 11520 1914 11529
rect 1858 11455 1914 11464
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1674 10976 1730 10985
rect 1674 10911 1730 10920
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1492 10736 1544 10742
rect 1492 10678 1544 10684
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 8922 1532 9862
rect 1584 9716 1636 9722
rect 1584 9658 1636 9664
rect 1596 9489 1624 9658
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1688 9110 1716 10911
rect 1766 9888 1822 9897
rect 1766 9823 1822 9832
rect 1676 9104 1728 9110
rect 1676 9046 1728 9052
rect 1676 8968 1728 8974
rect 1504 8916 1676 8922
rect 1504 8910 1728 8916
rect 1504 8894 1716 8910
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1306 8528 1362 8537
rect 1306 8463 1362 8472
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1228 6390 1256 6831
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 1216 6384 1268 6390
rect 1320 6361 1348 6394
rect 1216 6326 1268 6332
rect 1306 6352 1362 6361
rect 1306 6287 1362 6296
rect 1308 6180 1360 6186
rect 1308 6122 1360 6128
rect 1320 5817 1348 6122
rect 1412 6118 1440 8191
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1306 5808 1362 5817
rect 1306 5743 1362 5752
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1320 2514 1348 5170
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1412 3670 1440 4927
rect 1504 4826 1532 7346
rect 1596 6866 1624 8735
rect 1674 7712 1730 7721
rect 1674 7647 1730 7656
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1582 6080 1638 6089
rect 1582 6015 1638 6024
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 1400 3664 1452 3670
rect 1400 3606 1452 3612
rect 1596 3194 1624 6015
rect 1688 4010 1716 7647
rect 1780 7546 1808 9823
rect 1872 8090 1900 11455
rect 1964 11150 1992 13670
rect 2056 13394 2084 16000
rect 2148 15162 2176 16186
rect 2240 16182 2268 19858
rect 2332 18766 2360 20703
rect 2608 20466 2636 20975
rect 2792 20942 2820 22374
rect 2884 21078 2912 22528
rect 2872 21072 2924 21078
rect 2872 21014 2924 21020
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2332 18290 2360 18702
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2424 17134 2452 20198
rect 2608 19854 2636 20402
rect 2792 20058 2820 20878
rect 2976 20806 3004 27066
rect 3252 26874 3280 27118
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 3436 26908 3464 28206
rect 3516 28076 3568 28082
rect 3516 28018 3568 28024
rect 3068 26846 3280 26874
rect 3344 26880 3464 26908
rect 3068 24818 3096 26846
rect 3240 26784 3292 26790
rect 3240 26726 3292 26732
rect 3252 26314 3280 26726
rect 3240 26308 3292 26314
rect 3240 26250 3292 26256
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3056 24812 3108 24818
rect 3056 24754 3108 24760
rect 3068 24410 3096 24754
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3160 22778 3188 25638
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3252 22778 3280 24754
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3068 22234 3096 22714
rect 3146 22672 3202 22681
rect 3146 22607 3202 22616
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2964 20800 3016 20806
rect 2964 20742 3016 20748
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2976 20233 3004 20334
rect 2962 20224 3018 20233
rect 2962 20159 3018 20168
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2596 19848 2648 19854
rect 3068 19825 3096 21830
rect 2596 19790 2648 19796
rect 3054 19816 3110 19825
rect 2608 19378 2636 19790
rect 3054 19751 3110 19760
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2594 18456 2650 18465
rect 2516 18414 2594 18442
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 15201 2360 15302
rect 2318 15192 2374 15201
rect 2136 15156 2188 15162
rect 2318 15127 2374 15136
rect 2136 15098 2188 15104
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 11506 2084 12582
rect 2148 12306 2176 14350
rect 2332 13734 2360 15030
rect 2516 14532 2544 18414
rect 2594 18391 2650 18400
rect 2594 18320 2650 18329
rect 2594 18255 2650 18264
rect 2608 17660 2636 18255
rect 2700 17882 2728 19110
rect 2872 18624 2924 18630
rect 2872 18566 2924 18572
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2792 17678 2820 17818
rect 2688 17672 2740 17678
rect 2608 17632 2688 17660
rect 2608 17134 2636 17632
rect 2688 17614 2740 17620
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 17354 2820 17614
rect 2700 17326 2820 17354
rect 2596 17128 2648 17134
rect 2596 17070 2648 17076
rect 2424 14504 2544 14532
rect 2424 13938 2452 14504
rect 2608 14362 2636 17070
rect 2700 16674 2728 17326
rect 2884 17202 2912 18566
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17678 3004 18022
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2870 16688 2926 16697
rect 2700 16646 2820 16674
rect 2688 16448 2740 16454
rect 2686 16416 2688 16425
rect 2740 16416 2742 16425
rect 2686 16351 2742 16360
rect 2792 16114 2820 16646
rect 2870 16623 2926 16632
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2884 15706 2912 16623
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2976 16250 3004 16458
rect 3056 16448 3108 16454
rect 3056 16390 3108 16396
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3068 16153 3096 16390
rect 3054 16144 3110 16153
rect 3054 16079 3110 16088
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 14618 2912 14758
rect 2976 14634 3004 15982
rect 3054 15600 3110 15609
rect 3054 15535 3110 15544
rect 3068 14822 3096 15535
rect 3160 15094 3188 22607
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3252 22137 3280 22170
rect 3238 22128 3294 22137
rect 3238 22063 3294 22072
rect 3238 21856 3294 21865
rect 3238 21791 3294 21800
rect 3252 15502 3280 21791
rect 3344 19836 3372 26880
rect 3528 26586 3556 28018
rect 3804 26994 3832 28494
rect 4158 28455 4214 28464
rect 3976 28212 4028 28218
rect 3976 28154 4028 28160
rect 3988 28098 4016 28154
rect 4264 28150 4292 30534
rect 4356 30518 4476 30546
rect 4160 28144 4212 28150
rect 4066 28112 4122 28121
rect 3988 28070 4066 28098
rect 4160 28086 4212 28092
rect 4252 28144 4304 28150
rect 4252 28086 4304 28092
rect 4066 28047 4122 28056
rect 4172 27996 4200 28086
rect 4172 27985 4292 27996
rect 4172 27976 4306 27985
rect 4172 27968 4250 27976
rect 4250 27911 4306 27920
rect 3917 27772 4225 27781
rect 3917 27770 3923 27772
rect 3979 27770 4003 27772
rect 4059 27770 4083 27772
rect 4139 27770 4163 27772
rect 4219 27770 4225 27772
rect 3979 27718 3981 27770
rect 4161 27718 4163 27770
rect 3917 27716 3923 27718
rect 3979 27716 4003 27718
rect 4059 27716 4083 27718
rect 4139 27716 4163 27718
rect 4219 27716 4225 27718
rect 3917 27707 4225 27716
rect 3792 26988 3844 26994
rect 3712 26948 3792 26976
rect 3608 26920 3660 26926
rect 3608 26862 3660 26868
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 3516 26444 3568 26450
rect 3516 26386 3568 26392
rect 3424 26376 3476 26382
rect 3424 26318 3476 26324
rect 3436 25945 3464 26318
rect 3422 25936 3478 25945
rect 3422 25871 3478 25880
rect 3528 25294 3556 26386
rect 3516 25288 3568 25294
rect 3516 25230 3568 25236
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3436 24206 3464 24754
rect 3516 24744 3568 24750
rect 3516 24686 3568 24692
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3528 23866 3556 24686
rect 3620 24290 3648 26862
rect 3712 25702 3740 26948
rect 3792 26930 3844 26936
rect 3917 26684 4225 26693
rect 3917 26682 3923 26684
rect 3979 26682 4003 26684
rect 4059 26682 4083 26684
rect 4139 26682 4163 26684
rect 4219 26682 4225 26684
rect 3979 26630 3981 26682
rect 4161 26630 4163 26682
rect 3917 26628 3923 26630
rect 3979 26628 4003 26630
rect 4059 26628 4083 26630
rect 4139 26628 4163 26630
rect 4219 26628 4225 26630
rect 3917 26619 4225 26628
rect 4264 26450 4292 27911
rect 4252 26444 4304 26450
rect 4252 26386 4304 26392
rect 3792 26376 3844 26382
rect 3792 26318 3844 26324
rect 3804 26217 3832 26318
rect 3790 26208 3846 26217
rect 3790 26143 3846 26152
rect 4252 25900 4304 25906
rect 4356 25888 4384 30518
rect 4436 30388 4488 30394
rect 4436 30330 4488 30336
rect 4448 27849 4476 30330
rect 4528 30252 4580 30258
rect 4528 30194 4580 30200
rect 4540 29306 4568 30194
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4528 28144 4580 28150
rect 4528 28086 4580 28092
rect 4434 27840 4490 27849
rect 4434 27775 4490 27784
rect 4448 27554 4476 27775
rect 4540 27674 4568 28086
rect 4528 27668 4580 27674
rect 4528 27610 4580 27616
rect 4448 27526 4568 27554
rect 4436 27464 4488 27470
rect 4436 27406 4488 27412
rect 4304 25860 4384 25888
rect 4252 25842 4304 25848
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3712 25430 3740 25638
rect 3917 25596 4225 25605
rect 3917 25594 3923 25596
rect 3979 25594 4003 25596
rect 4059 25594 4083 25596
rect 4139 25594 4163 25596
rect 4219 25594 4225 25596
rect 3979 25542 3981 25594
rect 4161 25542 4163 25594
rect 3917 25540 3923 25542
rect 3979 25540 4003 25542
rect 4059 25540 4083 25542
rect 4139 25540 4163 25542
rect 4219 25540 4225 25542
rect 3917 25531 4225 25540
rect 3700 25424 3752 25430
rect 3700 25366 3752 25372
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3884 25152 3936 25158
rect 3884 25094 3936 25100
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 3712 24954 3740 25094
rect 3700 24948 3752 24954
rect 3700 24890 3752 24896
rect 3896 24886 3924 25094
rect 3884 24880 3936 24886
rect 3884 24822 3936 24828
rect 4080 24682 4108 25094
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3917 24508 4225 24517
rect 3917 24506 3923 24508
rect 3979 24506 4003 24508
rect 4059 24506 4083 24508
rect 4139 24506 4163 24508
rect 4219 24506 4225 24508
rect 3979 24454 3981 24506
rect 4161 24454 4163 24506
rect 3917 24452 3923 24454
rect 3979 24452 4003 24454
rect 4059 24452 4083 24454
rect 4139 24452 4163 24454
rect 4219 24452 4225 24454
rect 3917 24443 4225 24452
rect 3620 24262 3832 24290
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3608 23792 3660 23798
rect 3608 23734 3660 23740
rect 3516 23588 3568 23594
rect 3516 23530 3568 23536
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 3436 21729 3464 23258
rect 3528 23254 3556 23530
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3620 22234 3648 23734
rect 3516 22228 3568 22234
rect 3516 22170 3568 22176
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3528 22012 3556 22170
rect 3608 22024 3660 22030
rect 3528 21984 3608 22012
rect 3608 21966 3660 21972
rect 3422 21720 3478 21729
rect 3422 21655 3478 21664
rect 3712 20482 3740 24142
rect 3804 22234 3832 24262
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4066 24168 4122 24177
rect 4066 24103 4122 24112
rect 4080 23866 4108 24103
rect 4172 24070 4200 24210
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 3917 23420 4225 23429
rect 3917 23418 3923 23420
rect 3979 23418 4003 23420
rect 4059 23418 4083 23420
rect 4139 23418 4163 23420
rect 4219 23418 4225 23420
rect 3979 23366 3981 23418
rect 4161 23366 4163 23418
rect 3917 23364 3923 23366
rect 3979 23364 4003 23366
rect 4059 23364 4083 23366
rect 4139 23364 4163 23366
rect 4219 23364 4225 23366
rect 3917 23355 4225 23364
rect 4264 23304 4292 25842
rect 4448 25820 4476 27406
rect 4540 27062 4568 27526
rect 4528 27056 4580 27062
rect 4528 26998 4580 27004
rect 4528 26920 4580 26926
rect 4528 26862 4580 26868
rect 4540 26450 4568 26862
rect 4528 26444 4580 26450
rect 4528 26386 4580 26392
rect 4172 23276 4292 23304
rect 4356 25792 4476 25820
rect 3976 23248 4028 23254
rect 3976 23190 4028 23196
rect 3988 22953 4016 23190
rect 3974 22944 4030 22953
rect 3974 22879 4030 22888
rect 4172 22556 4200 23276
rect 4356 22778 4384 25792
rect 4436 25696 4488 25702
rect 4436 25638 4488 25644
rect 4448 25226 4476 25638
rect 4436 25220 4488 25226
rect 4436 25162 4488 25168
rect 4632 24682 4660 32184
rect 4712 30388 4764 30394
rect 4712 30330 4764 30336
rect 4724 29850 4752 30330
rect 4712 29844 4764 29850
rect 4712 29786 4764 29792
rect 4710 29744 4766 29753
rect 4710 29679 4766 29688
rect 4724 24954 4752 29679
rect 4816 28082 4844 36110
rect 4908 36038 4936 36672
rect 4896 36032 4948 36038
rect 4896 35974 4948 35980
rect 4896 35556 4948 35562
rect 4896 35498 4948 35504
rect 4908 33674 4936 35498
rect 5000 34921 5028 37198
rect 5092 36174 5120 38286
rect 5080 36168 5132 36174
rect 5080 36110 5132 36116
rect 5080 36032 5132 36038
rect 5080 35974 5132 35980
rect 5092 34950 5120 35974
rect 5080 34944 5132 34950
rect 4986 34912 5042 34921
rect 5080 34886 5132 34892
rect 4986 34847 5042 34856
rect 5092 34746 5120 34886
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 5080 34740 5132 34746
rect 5080 34682 5132 34688
rect 5000 34474 5028 34682
rect 5078 34640 5134 34649
rect 5078 34575 5080 34584
rect 5132 34575 5134 34584
rect 5080 34546 5132 34552
rect 4988 34468 5040 34474
rect 4988 34410 5040 34416
rect 4908 33646 5120 33674
rect 4896 33584 4948 33590
rect 4896 33526 4948 33532
rect 4908 33046 4936 33526
rect 4896 33040 4948 33046
rect 4896 32982 4948 32988
rect 4988 32564 5040 32570
rect 4988 32506 5040 32512
rect 4896 31816 4948 31822
rect 4896 31758 4948 31764
rect 4908 31113 4936 31758
rect 4894 31104 4950 31113
rect 4894 31039 4950 31048
rect 4908 30433 4936 31039
rect 4894 30424 4950 30433
rect 4894 30359 4950 30368
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4908 29102 4936 29990
rect 5000 29594 5028 32506
rect 5092 30138 5120 33646
rect 5184 32026 5212 40412
rect 5276 39137 5304 40666
rect 5368 39846 5396 43590
rect 5552 43450 5580 43846
rect 5540 43444 5592 43450
rect 5540 43386 5592 43392
rect 5540 42832 5592 42838
rect 5460 42792 5540 42820
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5460 39506 5488 42792
rect 5540 42774 5592 42780
rect 5540 42696 5592 42702
rect 5540 42638 5592 42644
rect 5552 41818 5580 42638
rect 5736 42566 5764 44463
rect 6012 43602 6040 44463
rect 6012 43574 6132 43602
rect 6000 43308 6052 43314
rect 6000 43250 6052 43256
rect 6012 42752 6040 43250
rect 6104 42906 6132 43574
rect 6288 43450 6316 44463
rect 6276 43444 6328 43450
rect 6276 43386 6328 43392
rect 6564 43330 6592 44463
rect 6840 44418 6868 44463
rect 6748 44390 6868 44418
rect 6748 43432 6776 44390
rect 7116 43738 7144 44463
rect 7392 43874 7420 44463
rect 7392 43846 7512 43874
rect 7116 43710 7420 43738
rect 6884 43548 7192 43557
rect 6884 43546 6890 43548
rect 6946 43546 6970 43548
rect 7026 43546 7050 43548
rect 7106 43546 7130 43548
rect 7186 43546 7192 43548
rect 6946 43494 6948 43546
rect 7128 43494 7130 43546
rect 6884 43492 6890 43494
rect 6946 43492 6970 43494
rect 7026 43492 7050 43494
rect 7106 43492 7130 43494
rect 7186 43492 7192 43494
rect 6884 43483 7192 43492
rect 6828 43444 6880 43450
rect 6748 43404 6828 43432
rect 6828 43386 6880 43392
rect 6276 43308 6328 43314
rect 6564 43302 6868 43330
rect 6276 43250 6328 43256
rect 6092 42900 6144 42906
rect 6092 42842 6144 42848
rect 6012 42724 6132 42752
rect 6000 42628 6052 42634
rect 6000 42570 6052 42576
rect 5724 42560 5776 42566
rect 5724 42502 5776 42508
rect 5908 42560 5960 42566
rect 5908 42502 5960 42508
rect 5724 42220 5776 42226
rect 5776 42180 5856 42208
rect 5724 42162 5776 42168
rect 5632 42084 5684 42090
rect 5632 42026 5684 42032
rect 5540 41812 5592 41818
rect 5540 41754 5592 41760
rect 5644 41614 5672 42026
rect 5724 42016 5776 42022
rect 5724 41958 5776 41964
rect 5736 41614 5764 41958
rect 5632 41608 5684 41614
rect 5632 41550 5684 41556
rect 5724 41608 5776 41614
rect 5724 41550 5776 41556
rect 5828 41414 5856 42180
rect 5920 41818 5948 42502
rect 6012 41818 6040 42570
rect 5908 41812 5960 41818
rect 5908 41754 5960 41760
rect 6000 41812 6052 41818
rect 6000 41754 6052 41760
rect 6104 41478 6132 42724
rect 6288 42362 6316 43250
rect 6840 42906 6868 43302
rect 7288 43308 7340 43314
rect 7288 43250 7340 43256
rect 6828 42900 6880 42906
rect 6828 42842 6880 42848
rect 7300 42752 7328 43250
rect 7392 42906 7420 43710
rect 7380 42900 7432 42906
rect 7380 42842 7432 42848
rect 7300 42724 7420 42752
rect 7288 42628 7340 42634
rect 7288 42570 7340 42576
rect 6884 42460 7192 42469
rect 6884 42458 6890 42460
rect 6946 42458 6970 42460
rect 7026 42458 7050 42460
rect 7106 42458 7130 42460
rect 7186 42458 7192 42460
rect 6946 42406 6948 42458
rect 7128 42406 7130 42458
rect 6884 42404 6890 42406
rect 6946 42404 6970 42406
rect 7026 42404 7050 42406
rect 7106 42404 7130 42406
rect 7186 42404 7192 42406
rect 6884 42395 7192 42404
rect 6276 42356 6328 42362
rect 6276 42298 6328 42304
rect 7012 42356 7064 42362
rect 7012 42298 7064 42304
rect 6184 42220 6236 42226
rect 6184 42162 6236 42168
rect 6552 42220 6604 42226
rect 6552 42162 6604 42168
rect 6196 41857 6224 42162
rect 6460 42084 6512 42090
rect 6460 42026 6512 42032
rect 6182 41848 6238 41857
rect 6182 41783 6238 41792
rect 6092 41472 6144 41478
rect 6092 41414 6144 41420
rect 6472 41414 6500 42026
rect 6564 41721 6592 42162
rect 6920 42016 6972 42022
rect 6920 41958 6972 41964
rect 6932 41818 6960 41958
rect 6920 41812 6972 41818
rect 6920 41754 6972 41760
rect 6550 41712 6606 41721
rect 6550 41647 6606 41656
rect 6736 41608 6788 41614
rect 6734 41576 6736 41585
rect 6788 41576 6790 41585
rect 7024 41546 7052 42298
rect 7196 42152 7248 42158
rect 7196 42094 7248 42100
rect 7208 41698 7236 42094
rect 7300 41818 7328 42570
rect 7392 42362 7420 42724
rect 7484 42566 7512 43846
rect 7668 43450 7696 44463
rect 7944 43450 7972 44463
rect 7656 43444 7708 43450
rect 7656 43386 7708 43392
rect 7932 43444 7984 43450
rect 7932 43386 7984 43392
rect 8116 43308 8168 43314
rect 8116 43250 8168 43256
rect 7564 42696 7616 42702
rect 7564 42638 7616 42644
rect 7472 42560 7524 42566
rect 7472 42502 7524 42508
rect 7380 42356 7432 42362
rect 7380 42298 7432 42304
rect 7380 42220 7432 42226
rect 7380 42162 7432 42168
rect 7392 42129 7420 42162
rect 7378 42120 7434 42129
rect 7378 42055 7434 42064
rect 7380 42016 7432 42022
rect 7380 41958 7432 41964
rect 7472 42016 7524 42022
rect 7472 41958 7524 41964
rect 7392 41818 7420 41958
rect 7484 41818 7512 41958
rect 7576 41818 7604 42638
rect 7656 42220 7708 42226
rect 7656 42162 7708 42168
rect 7932 42220 7984 42226
rect 7932 42162 7984 42168
rect 7668 41857 7696 42162
rect 7840 42152 7892 42158
rect 7840 42094 7892 42100
rect 7748 42016 7800 42022
rect 7748 41958 7800 41964
rect 7654 41848 7710 41857
rect 7288 41812 7340 41818
rect 7288 41754 7340 41760
rect 7380 41812 7432 41818
rect 7380 41754 7432 41760
rect 7472 41812 7524 41818
rect 7472 41754 7524 41760
rect 7564 41812 7616 41818
rect 7760 41818 7788 41958
rect 7654 41783 7710 41792
rect 7748 41812 7800 41818
rect 7564 41754 7616 41760
rect 7748 41754 7800 41760
rect 7208 41670 7328 41698
rect 6734 41511 6790 41520
rect 7012 41540 7064 41546
rect 7012 41482 7064 41488
rect 7300 41478 7328 41670
rect 7288 41472 7340 41478
rect 7288 41414 7340 41420
rect 5736 41386 5856 41414
rect 6380 41386 6500 41414
rect 5448 39500 5500 39506
rect 5448 39442 5500 39448
rect 5356 39296 5408 39302
rect 5356 39238 5408 39244
rect 5262 39128 5318 39137
rect 5368 39098 5396 39238
rect 5262 39063 5318 39072
rect 5356 39092 5408 39098
rect 5276 38962 5304 39063
rect 5356 39034 5408 39040
rect 5264 38956 5316 38962
rect 5264 38898 5316 38904
rect 5264 38752 5316 38758
rect 5264 38694 5316 38700
rect 5276 38554 5304 38694
rect 5264 38548 5316 38554
rect 5264 38490 5316 38496
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5630 38312 5686 38321
rect 5356 38208 5408 38214
rect 5356 38150 5408 38156
rect 5264 37664 5316 37670
rect 5264 37606 5316 37612
rect 5276 36224 5304 37606
rect 5368 37262 5396 38150
rect 5552 37369 5580 38286
rect 5630 38247 5686 38256
rect 5644 37466 5672 38247
rect 5736 37890 5764 41386
rect 5816 40928 5868 40934
rect 5816 40870 5868 40876
rect 6000 40928 6052 40934
rect 6000 40870 6052 40876
rect 5828 40633 5856 40870
rect 5814 40624 5870 40633
rect 5814 40559 5870 40568
rect 5828 40526 5856 40559
rect 5816 40520 5868 40526
rect 5816 40462 5868 40468
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5920 39642 5948 39782
rect 5908 39636 5960 39642
rect 5908 39578 5960 39584
rect 5908 38888 5960 38894
rect 5908 38830 5960 38836
rect 5814 37904 5870 37913
rect 5736 37862 5814 37890
rect 5814 37839 5870 37848
rect 5632 37460 5684 37466
rect 5632 37402 5684 37408
rect 5538 37360 5594 37369
rect 5538 37295 5594 37304
rect 5356 37256 5408 37262
rect 5356 37198 5408 37204
rect 5724 37256 5776 37262
rect 5920 37210 5948 38830
rect 6012 38486 6040 40870
rect 6380 40458 6408 41386
rect 6884 41372 7192 41381
rect 6884 41370 6890 41372
rect 6946 41370 6970 41372
rect 7026 41370 7050 41372
rect 7106 41370 7130 41372
rect 7186 41370 7192 41372
rect 6946 41318 6948 41370
rect 7128 41318 7130 41370
rect 6884 41316 6890 41318
rect 6946 41316 6970 41318
rect 7026 41316 7050 41318
rect 7106 41316 7130 41318
rect 7186 41316 7192 41318
rect 6884 41307 7192 41316
rect 6828 40520 6880 40526
rect 6826 40488 6828 40497
rect 6880 40488 6882 40497
rect 6092 40452 6144 40458
rect 6092 40394 6144 40400
rect 6368 40452 6420 40458
rect 6368 40394 6420 40400
rect 6748 40446 6826 40474
rect 6000 38480 6052 38486
rect 6000 38422 6052 38428
rect 6104 37806 6132 40394
rect 6644 40384 6696 40390
rect 6644 40326 6696 40332
rect 6656 39506 6684 40326
rect 6748 39794 6776 40446
rect 6826 40423 6882 40432
rect 6884 40284 7192 40293
rect 6884 40282 6890 40284
rect 6946 40282 6970 40284
rect 7026 40282 7050 40284
rect 7106 40282 7130 40284
rect 7186 40282 7192 40284
rect 6946 40230 6948 40282
rect 7128 40230 7130 40282
rect 6884 40228 6890 40230
rect 6946 40228 6970 40230
rect 7026 40228 7050 40230
rect 7106 40228 7130 40230
rect 7186 40228 7192 40230
rect 6884 40219 7192 40228
rect 6748 39766 6868 39794
rect 6736 39636 6788 39642
rect 6736 39578 6788 39584
rect 6644 39500 6696 39506
rect 6644 39442 6696 39448
rect 6368 39432 6420 39438
rect 6368 39374 6420 39380
rect 6380 39098 6408 39374
rect 6368 39092 6420 39098
rect 6368 39034 6420 39040
rect 6276 38344 6328 38350
rect 6276 38286 6328 38292
rect 6552 38344 6604 38350
rect 6552 38286 6604 38292
rect 6092 37800 6144 37806
rect 6092 37742 6144 37748
rect 5724 37198 5776 37204
rect 5448 37120 5500 37126
rect 5448 37062 5500 37068
rect 5460 36310 5488 37062
rect 5448 36304 5500 36310
rect 5448 36246 5500 36252
rect 5356 36236 5408 36242
rect 5276 36196 5356 36224
rect 5276 35834 5304 36196
rect 5356 36178 5408 36184
rect 5264 35828 5316 35834
rect 5264 35770 5316 35776
rect 5264 35624 5316 35630
rect 5264 35566 5316 35572
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 5276 34950 5304 35566
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 5276 30240 5304 34886
rect 5368 32774 5396 35566
rect 5460 35494 5488 36246
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5448 35488 5500 35494
rect 5448 35430 5500 35436
rect 5448 35216 5500 35222
rect 5446 35184 5448 35193
rect 5500 35184 5502 35193
rect 5446 35119 5502 35128
rect 5448 35080 5500 35086
rect 5448 35022 5500 35028
rect 5460 34950 5488 35022
rect 5448 34944 5500 34950
rect 5448 34886 5500 34892
rect 5460 34610 5488 34886
rect 5448 34604 5500 34610
rect 5448 34546 5500 34552
rect 5552 34513 5580 35974
rect 5630 35592 5686 35601
rect 5630 35527 5686 35536
rect 5644 35086 5672 35527
rect 5632 35080 5684 35086
rect 5632 35022 5684 35028
rect 5538 34504 5594 34513
rect 5538 34439 5594 34448
rect 5448 34400 5500 34406
rect 5448 34342 5500 34348
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5460 32586 5488 34342
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5552 32978 5580 33798
rect 5540 32972 5592 32978
rect 5540 32914 5592 32920
rect 5368 32558 5488 32586
rect 5368 32230 5396 32558
rect 5644 32298 5672 35022
rect 5736 34950 5764 37198
rect 5828 37182 5948 37210
rect 5724 34944 5776 34950
rect 5724 34886 5776 34892
rect 5724 34604 5776 34610
rect 5724 34546 5776 34552
rect 5736 34202 5764 34546
rect 5724 34196 5776 34202
rect 5724 34138 5776 34144
rect 5828 32858 5856 37182
rect 5908 37120 5960 37126
rect 5908 37062 5960 37068
rect 5920 35057 5948 37062
rect 6000 36168 6052 36174
rect 6000 36110 6052 36116
rect 6012 35494 6040 36110
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 6104 35136 6132 37742
rect 6288 37670 6316 38286
rect 6564 38010 6592 38286
rect 6552 38004 6604 38010
rect 6552 37946 6604 37952
rect 6276 37664 6328 37670
rect 6276 37606 6328 37612
rect 6552 37460 6604 37466
rect 6552 37402 6604 37408
rect 6460 36236 6512 36242
rect 6380 36196 6460 36224
rect 6380 35562 6408 36196
rect 6460 36178 6512 36184
rect 6368 35556 6420 35562
rect 6368 35498 6420 35504
rect 6380 35290 6408 35498
rect 6460 35488 6512 35494
rect 6460 35430 6512 35436
rect 6368 35284 6420 35290
rect 6368 35226 6420 35232
rect 6012 35108 6132 35136
rect 5906 35048 5962 35057
rect 5906 34983 5962 34992
rect 5920 33522 5948 34983
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 5920 32910 5948 33254
rect 5736 32830 5856 32858
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 5736 32502 5764 32830
rect 5908 32768 5960 32774
rect 5908 32710 5960 32716
rect 5724 32496 5776 32502
rect 5724 32438 5776 32444
rect 5632 32292 5684 32298
rect 5632 32234 5684 32240
rect 5356 32224 5408 32230
rect 5356 32166 5408 32172
rect 5368 30734 5396 32166
rect 5540 31816 5592 31822
rect 5920 31793 5948 32710
rect 5540 31758 5592 31764
rect 5906 31784 5962 31793
rect 5552 31498 5580 31758
rect 5906 31719 5962 31728
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5828 31498 5856 31622
rect 6012 31498 6040 35108
rect 6184 34536 6236 34542
rect 6184 34478 6236 34484
rect 6196 33969 6224 34478
rect 6368 34060 6420 34066
rect 6368 34002 6420 34008
rect 6182 33960 6238 33969
rect 6182 33895 6238 33904
rect 6276 33924 6328 33930
rect 6196 32978 6224 33895
rect 6276 33866 6328 33872
rect 6288 33289 6316 33866
rect 6274 33280 6330 33289
rect 6274 33215 6330 33224
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6104 32570 6132 32710
rect 6092 32564 6144 32570
rect 6092 32506 6144 32512
rect 6092 32428 6144 32434
rect 6092 32370 6144 32376
rect 6104 31822 6132 32370
rect 6196 32042 6224 32914
rect 6276 32768 6328 32774
rect 6276 32710 6328 32716
rect 6288 32570 6316 32710
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 6196 32014 6316 32042
rect 6092 31816 6144 31822
rect 6092 31758 6144 31764
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 5552 31470 5856 31498
rect 5448 31408 5500 31414
rect 5446 31376 5448 31385
rect 5500 31376 5502 31385
rect 5446 31311 5502 31320
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 5448 31204 5500 31210
rect 5448 31146 5500 31152
rect 5460 30841 5488 31146
rect 5446 30832 5502 30841
rect 5446 30767 5502 30776
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5276 30212 5488 30240
rect 5092 30110 5304 30138
rect 5172 30048 5224 30054
rect 5172 29990 5224 29996
rect 5184 29714 5212 29990
rect 5172 29708 5224 29714
rect 5172 29650 5224 29656
rect 5000 29566 5120 29594
rect 4988 29504 5040 29510
rect 4988 29446 5040 29452
rect 5000 29238 5028 29446
rect 4988 29232 5040 29238
rect 4988 29174 5040 29180
rect 4896 29096 4948 29102
rect 4896 29038 4948 29044
rect 4986 28792 5042 28801
rect 4986 28727 5042 28736
rect 5000 28529 5028 28727
rect 4986 28520 5042 28529
rect 4986 28455 5042 28464
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4620 24676 4672 24682
rect 4620 24618 4672 24624
rect 4528 24268 4580 24274
rect 4528 24210 4580 24216
rect 4436 24132 4488 24138
rect 4436 24074 4488 24080
rect 4448 22778 4476 24074
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4252 22704 4304 22710
rect 4304 22652 4476 22658
rect 4252 22646 4476 22652
rect 4264 22630 4476 22646
rect 4172 22528 4384 22556
rect 3917 22332 4225 22341
rect 3917 22330 3923 22332
rect 3979 22330 4003 22332
rect 4059 22330 4083 22332
rect 4139 22330 4163 22332
rect 4219 22330 4225 22332
rect 3979 22278 3981 22330
rect 4161 22278 4163 22330
rect 3917 22276 3923 22278
rect 3979 22276 4003 22278
rect 4059 22276 4083 22278
rect 4139 22276 4163 22278
rect 4219 22276 4225 22278
rect 3917 22267 4225 22276
rect 3792 22228 3844 22234
rect 3792 22170 3844 22176
rect 3804 20602 3832 22170
rect 3974 22128 4030 22137
rect 3974 22063 4030 22072
rect 3988 21962 4016 22063
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 4080 21690 4108 21830
rect 4068 21684 4120 21690
rect 4068 21626 4120 21632
rect 3917 21244 4225 21253
rect 3917 21242 3923 21244
rect 3979 21242 4003 21244
rect 4059 21242 4083 21244
rect 4139 21242 4163 21244
rect 4219 21242 4225 21244
rect 3979 21190 3981 21242
rect 4161 21190 4163 21242
rect 3917 21188 3923 21190
rect 3979 21188 4003 21190
rect 4059 21188 4083 21190
rect 4139 21188 4163 21190
rect 4219 21188 4225 21190
rect 3917 21179 4225 21188
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 4068 20800 4120 20806
rect 4172 20777 4200 20878
rect 4068 20742 4120 20748
rect 4158 20768 4214 20777
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3712 20466 3924 20482
rect 4080 20466 4108 20742
rect 4158 20703 4214 20712
rect 3712 20460 3936 20466
rect 3712 20454 3884 20460
rect 3516 20324 3568 20330
rect 3516 20266 3568 20272
rect 3528 20058 3556 20266
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3344 19808 3464 19836
rect 3332 19372 3384 19378
rect 3332 19314 3384 19320
rect 3344 19145 3372 19314
rect 3330 19136 3386 19145
rect 3330 19071 3386 19080
rect 3436 17728 3464 19808
rect 3712 17882 3740 20454
rect 3884 20402 3936 20408
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 3917 20156 4225 20165
rect 3917 20154 3923 20156
rect 3979 20154 4003 20156
rect 4059 20154 4083 20156
rect 4139 20154 4163 20156
rect 4219 20154 4225 20156
rect 3979 20102 3981 20154
rect 4161 20102 4163 20154
rect 3917 20100 3923 20102
rect 3979 20100 4003 20102
rect 4059 20100 4083 20102
rect 4139 20100 4163 20102
rect 4219 20100 4225 20102
rect 3917 20091 4225 20100
rect 4264 19310 4292 20334
rect 4252 19304 4304 19310
rect 4252 19246 4304 19252
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 3917 19068 4225 19077
rect 3917 19066 3923 19068
rect 3979 19066 4003 19068
rect 4059 19066 4083 19068
rect 4139 19066 4163 19068
rect 4219 19066 4225 19068
rect 3979 19014 3981 19066
rect 4161 19014 4163 19066
rect 3917 19012 3923 19014
rect 3979 19012 4003 19014
rect 4059 19012 4083 19014
rect 4139 19012 4163 19014
rect 4219 19012 4225 19014
rect 3917 19003 4225 19012
rect 3974 18864 4030 18873
rect 4030 18822 4108 18850
rect 3974 18799 4030 18808
rect 4080 18766 4108 18822
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3976 18624 4028 18630
rect 3976 18566 4028 18572
rect 3896 18204 3924 18566
rect 3988 18426 4016 18566
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3976 18216 4028 18222
rect 3896 18184 3976 18204
rect 4028 18184 4030 18193
rect 3896 18176 3974 18184
rect 3974 18119 4030 18128
rect 4080 18068 4108 18702
rect 4158 18456 4214 18465
rect 4264 18426 4292 19110
rect 4158 18391 4214 18400
rect 4252 18420 4304 18426
rect 4172 18272 4200 18391
rect 4252 18362 4304 18368
rect 4252 18284 4304 18290
rect 4172 18244 4252 18272
rect 4252 18226 4304 18232
rect 4080 18040 4292 18068
rect 3917 17980 4225 17989
rect 3917 17978 3923 17980
rect 3979 17978 4003 17980
rect 4059 17978 4083 17980
rect 4139 17978 4163 17980
rect 4219 17978 4225 17980
rect 3979 17926 3981 17978
rect 4161 17926 4163 17978
rect 3917 17924 3923 17926
rect 3979 17924 4003 17926
rect 4059 17924 4083 17926
rect 4139 17924 4163 17926
rect 4219 17924 4225 17926
rect 3917 17915 4225 17924
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3608 17808 3660 17814
rect 3974 17776 4030 17785
rect 3660 17756 3740 17762
rect 3608 17750 3740 17756
rect 3516 17740 3568 17746
rect 3436 17700 3516 17728
rect 3620 17734 3740 17750
rect 3516 17682 3568 17688
rect 3608 17536 3660 17542
rect 3608 17478 3660 17484
rect 3620 17338 3648 17478
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3330 17232 3386 17241
rect 3330 17167 3386 17176
rect 3344 16794 3372 17167
rect 3516 16992 3568 16998
rect 3436 16952 3516 16980
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3332 16584 3384 16590
rect 3332 16526 3384 16532
rect 3344 16454 3372 16526
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3330 16280 3386 16289
rect 3330 16215 3386 16224
rect 3344 16182 3372 16215
rect 3332 16176 3384 16182
rect 3332 16118 3384 16124
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15094 3280 15302
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3240 15088 3292 15094
rect 3240 15030 3292 15036
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2872 14612 2924 14618
rect 2976 14606 3096 14634
rect 2872 14554 2924 14560
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 2872 14476 2924 14482
rect 2688 14408 2740 14414
rect 2608 14356 2688 14362
rect 2608 14350 2740 14356
rect 2608 14334 2728 14350
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13002 2360 13670
rect 2332 12974 2452 13002
rect 2424 12918 2452 12974
rect 2412 12912 2464 12918
rect 2318 12880 2374 12889
rect 2412 12854 2464 12860
rect 2318 12815 2374 12824
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2240 11558 2268 12650
rect 2228 11552 2280 11558
rect 2056 11478 2176 11506
rect 2228 11494 2280 11500
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 2042 11112 2098 11121
rect 2042 11047 2098 11056
rect 2056 10554 2084 11047
rect 2148 10674 2176 11478
rect 2240 11234 2268 11494
rect 2332 11354 2360 12815
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2504 12300 2556 12306
rect 2608 12288 2636 14334
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 2556 12260 2636 12288
rect 2504 12242 2556 12248
rect 2424 11898 2452 12242
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2240 11206 2360 11234
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10810 2268 11018
rect 2228 10804 2280 10810
rect 2228 10746 2280 10752
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2056 10526 2176 10554
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 8566 1992 10406
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 2056 10033 2084 10066
rect 2042 10024 2098 10033
rect 2042 9959 2098 9968
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2056 9353 2084 9522
rect 2042 9344 2098 9353
rect 2042 9279 2098 9288
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2056 8090 2084 8434
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2148 7970 2176 10526
rect 2332 10470 2360 11206
rect 2320 10464 2372 10470
rect 2320 10406 2372 10412
rect 2332 9654 2360 10406
rect 2516 10266 2544 12242
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9722 2452 10066
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 1964 7942 2176 7970
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1766 7440 1822 7449
rect 1766 7375 1822 7384
rect 1780 5914 1808 7375
rect 1860 7336 1912 7342
rect 1860 7278 1912 7284
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1766 5400 1822 5409
rect 1766 5335 1822 5344
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1780 3738 1808 5335
rect 1872 4554 1900 7278
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1872 4010 1900 4490
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1768 3732 1820 3738
rect 1768 3674 1820 3680
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1872 3097 1900 3946
rect 1858 3088 1914 3097
rect 1858 3023 1914 3032
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1122 2272 1178 2281
rect 1122 2207 1178 2216
rect 1320 1970 1348 2450
rect 1308 1964 1360 1970
rect 1308 1906 1360 1912
rect 1400 1964 1452 1970
rect 1400 1906 1452 1912
rect 1412 1442 1440 1906
rect 1320 1414 1440 1442
rect 1320 160 1348 1414
rect 1964 1358 1992 7942
rect 2136 7880 2188 7886
rect 2134 7848 2136 7857
rect 2188 7848 2190 7857
rect 2044 7812 2096 7818
rect 2134 7783 2190 7792
rect 2044 7754 2096 7760
rect 2056 6866 2084 7754
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2148 6610 2176 7783
rect 2240 6798 2268 8910
rect 2332 8401 2360 9590
rect 2318 8392 2374 8401
rect 2318 8327 2374 8336
rect 2412 8288 2464 8294
rect 2412 8230 2464 8236
rect 2424 7818 2452 8230
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2516 7750 2544 9590
rect 2608 9042 2636 11494
rect 2700 11014 2728 14214
rect 2792 13530 2820 14447
rect 2872 14418 2924 14424
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 11937 2820 13194
rect 2884 12306 2912 14418
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 14074 3004 14350
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2976 12918 3004 13738
rect 2964 12912 3016 12918
rect 2964 12854 3016 12860
rect 3068 12782 3096 14606
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3252 12850 3280 13330
rect 3344 13297 3372 16118
rect 3330 13288 3386 13297
rect 3330 13223 3386 13232
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3056 12776 3108 12782
rect 3332 12776 3384 12782
rect 3056 12718 3108 12724
rect 3252 12724 3332 12730
rect 3252 12718 3384 12724
rect 3252 12702 3372 12718
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 3252 12220 3280 12702
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12306 3372 12582
rect 3332 12300 3384 12306
rect 3332 12242 3384 12248
rect 2962 12200 3018 12209
rect 2962 12135 3018 12144
rect 3068 12192 3280 12220
rect 2870 12064 2926 12073
rect 2870 11999 2926 12008
rect 2778 11928 2834 11937
rect 2778 11863 2834 11872
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2686 10024 2742 10033
rect 2686 9959 2742 9968
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2608 7546 2636 8842
rect 2700 8294 2728 9959
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2700 7342 2728 8230
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 2594 6760 2650 6769
rect 2594 6695 2596 6704
rect 2648 6695 2650 6704
rect 2596 6666 2648 6672
rect 2056 3398 2084 6598
rect 2148 6582 2268 6610
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 5914 2176 6258
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2148 4690 2176 5306
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2134 4448 2190 4457
rect 2134 4383 2190 4392
rect 2148 4146 2176 4383
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3738 2176 3878
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2240 3618 2268 6582
rect 2688 6384 2740 6390
rect 2608 6344 2688 6372
rect 2320 5704 2372 5710
rect 2318 5672 2320 5681
rect 2372 5672 2374 5681
rect 2318 5607 2374 5616
rect 2608 5370 2636 6344
rect 2688 6326 2740 6332
rect 2596 5364 2648 5370
rect 2596 5306 2648 5312
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2148 3590 2268 3618
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 2148 2774 2176 3590
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 2240 3194 2268 3402
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2332 3126 2360 4762
rect 2412 4684 2464 4690
rect 2412 4626 2464 4632
rect 2320 3120 2372 3126
rect 2320 3062 2372 3068
rect 2056 2746 2176 2774
rect 2056 1970 2084 2746
rect 2134 2680 2190 2689
rect 2134 2615 2136 2624
rect 2188 2615 2190 2624
rect 2136 2586 2188 2592
rect 2424 2106 2452 4626
rect 2516 3942 2544 4966
rect 2608 4146 2636 5306
rect 2700 4690 2728 5306
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2792 3670 2820 11018
rect 2884 10062 2912 11999
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2884 8498 2912 9658
rect 2976 9058 3004 12135
rect 3068 11098 3096 12192
rect 3146 11792 3202 11801
rect 3146 11727 3202 11736
rect 3332 11756 3384 11762
rect 3160 11286 3188 11727
rect 3332 11698 3384 11704
rect 3344 11665 3372 11698
rect 3330 11656 3386 11665
rect 3330 11591 3386 11600
rect 3238 11520 3294 11529
rect 3238 11455 3294 11464
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 3068 11070 3188 11098
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 3068 10169 3096 10950
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3068 9178 3096 9318
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2976 9030 3096 9058
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7342 3004 7686
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5273 2912 5510
rect 2870 5264 2926 5273
rect 2976 5234 3004 6734
rect 3068 5234 3096 9030
rect 3160 8616 3188 11070
rect 3252 9586 3280 11455
rect 3436 11132 3464 16952
rect 3516 16934 3568 16940
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 16250 3648 16526
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3712 16046 3740 17734
rect 3974 17711 4030 17720
rect 3988 17678 4016 17711
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4264 17338 4292 18040
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 3804 16522 3832 16934
rect 3917 16892 4225 16901
rect 3917 16890 3923 16892
rect 3979 16890 4003 16892
rect 4059 16890 4083 16892
rect 4139 16890 4163 16892
rect 4219 16890 4225 16892
rect 3979 16838 3981 16890
rect 4161 16838 4163 16890
rect 3917 16836 3923 16838
rect 3979 16836 4003 16838
rect 4059 16836 4083 16838
rect 4139 16836 4163 16838
rect 4219 16836 4225 16838
rect 3917 16827 4225 16836
rect 3792 16516 3844 16522
rect 3792 16458 3844 16464
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3514 15600 3570 15609
rect 3712 15570 3740 15846
rect 3917 15804 4225 15813
rect 3917 15802 3923 15804
rect 3979 15802 4003 15804
rect 4059 15802 4083 15804
rect 4139 15802 4163 15804
rect 4219 15802 4225 15804
rect 3979 15750 3981 15802
rect 4161 15750 4163 15802
rect 3917 15748 3923 15750
rect 3979 15748 4003 15750
rect 4059 15748 4083 15750
rect 4139 15748 4163 15750
rect 4219 15748 4225 15750
rect 3917 15739 4225 15748
rect 3514 15535 3570 15544
rect 3700 15564 3752 15570
rect 3528 15502 3556 15535
rect 3700 15506 3752 15512
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3712 15366 3740 15506
rect 4160 15496 4212 15502
rect 3974 15464 4030 15473
rect 4160 15438 4212 15444
rect 3974 15399 4030 15408
rect 3700 15360 3752 15366
rect 3700 15302 3752 15308
rect 3988 14822 4016 15399
rect 4172 15094 4200 15438
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3917 14716 4225 14725
rect 3917 14714 3923 14716
rect 3979 14714 4003 14716
rect 4059 14714 4083 14716
rect 4139 14714 4163 14716
rect 4219 14714 4225 14716
rect 3979 14662 3981 14714
rect 4161 14662 4163 14714
rect 3917 14660 3923 14662
rect 3979 14660 4003 14662
rect 4059 14660 4083 14662
rect 4139 14660 4163 14662
rect 4219 14660 4225 14662
rect 3917 14651 4225 14660
rect 4264 14600 4292 16390
rect 4356 16153 4384 22528
rect 4448 21185 4476 22630
rect 4434 21176 4490 21185
rect 4434 21111 4490 21120
rect 4436 20936 4488 20942
rect 4436 20878 4488 20884
rect 4448 19786 4476 20878
rect 4436 19780 4488 19786
rect 4436 19722 4488 19728
rect 4448 17134 4476 19722
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4342 16144 4398 16153
rect 4448 16114 4476 17070
rect 4540 16114 4568 24210
rect 4632 24138 4660 24618
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4620 23180 4672 23186
rect 4620 23122 4672 23128
rect 4632 22817 4660 23122
rect 4618 22808 4674 22817
rect 4618 22743 4674 22752
rect 4632 22710 4660 22743
rect 4620 22704 4672 22710
rect 4620 22646 4672 22652
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4632 22273 4660 22374
rect 4618 22264 4674 22273
rect 4618 22199 4674 22208
rect 4632 21690 4660 22199
rect 4724 22094 4752 24686
rect 4816 24274 4844 28018
rect 5000 28014 5028 28358
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 5000 27334 5028 27406
rect 4988 27328 5040 27334
rect 4988 27270 5040 27276
rect 4988 27056 5040 27062
rect 4988 26998 5040 27004
rect 5000 25673 5028 26998
rect 4986 25664 5042 25673
rect 4986 25599 5042 25608
rect 5092 25294 5120 29566
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5184 29073 5212 29106
rect 5170 29064 5226 29073
rect 5170 28999 5226 29008
rect 5276 28994 5304 30110
rect 5276 28966 5396 28994
rect 5264 28484 5316 28490
rect 5264 28426 5316 28432
rect 5172 28416 5224 28422
rect 5172 28358 5224 28364
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4804 24268 4856 24274
rect 4804 24210 4856 24216
rect 4908 23866 4936 24550
rect 5000 24206 5028 24890
rect 5092 24750 5120 25230
rect 5080 24744 5132 24750
rect 5080 24686 5132 24692
rect 5184 24732 5212 28358
rect 5276 28121 5304 28426
rect 5368 28150 5396 28966
rect 5460 28422 5488 30212
rect 5448 28416 5500 28422
rect 5448 28358 5500 28364
rect 5552 28257 5580 31282
rect 5828 29578 5856 31470
rect 5920 31470 6040 31498
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5724 29572 5776 29578
rect 5724 29514 5776 29520
rect 5816 29572 5868 29578
rect 5816 29514 5868 29520
rect 5644 29306 5672 29514
rect 5632 29300 5684 29306
rect 5632 29242 5684 29248
rect 5630 29064 5686 29073
rect 5630 28999 5686 29008
rect 5538 28248 5594 28257
rect 5538 28183 5594 28192
rect 5356 28144 5408 28150
rect 5262 28112 5318 28121
rect 5644 28098 5672 28999
rect 5356 28086 5408 28092
rect 5262 28047 5318 28056
rect 5448 28076 5500 28082
rect 5448 28018 5500 28024
rect 5552 28070 5672 28098
rect 5460 27130 5488 28018
rect 5552 27316 5580 28070
rect 5632 28008 5684 28014
rect 5630 27976 5632 27985
rect 5684 27976 5686 27985
rect 5630 27911 5686 27920
rect 5552 27288 5672 27316
rect 5448 27124 5500 27130
rect 5448 27066 5500 27072
rect 5356 26240 5408 26246
rect 5356 26182 5408 26188
rect 5538 26208 5594 26217
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5276 25362 5304 25638
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5276 24954 5304 25094
rect 5264 24948 5316 24954
rect 5264 24890 5316 24896
rect 5264 24744 5316 24750
rect 5184 24704 5264 24732
rect 5078 24304 5134 24313
rect 5184 24290 5212 24704
rect 5264 24686 5316 24692
rect 5134 24262 5212 24290
rect 5264 24268 5316 24274
rect 5078 24239 5134 24248
rect 5264 24210 5316 24216
rect 4988 24200 5040 24206
rect 4988 24142 5040 24148
rect 5276 24138 5304 24210
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4986 23488 5042 23497
rect 4986 23423 5042 23432
rect 4896 22636 4948 22642
rect 4896 22578 4948 22584
rect 4724 22066 4844 22094
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4618 21584 4674 21593
rect 4618 21519 4674 21528
rect 4632 21418 4660 21519
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4724 21078 4752 21830
rect 4816 21350 4844 22066
rect 4804 21344 4856 21350
rect 4908 21321 4936 22578
rect 4804 21286 4856 21292
rect 4894 21312 4950 21321
rect 4712 21072 4764 21078
rect 4712 21014 4764 21020
rect 4712 20256 4764 20262
rect 4712 20198 4764 20204
rect 4618 20088 4674 20097
rect 4618 20023 4674 20032
rect 4632 19514 4660 20023
rect 4724 19514 4752 20198
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4816 19394 4844 21286
rect 4894 21247 4950 21256
rect 4894 20904 4950 20913
rect 4894 20839 4950 20848
rect 4632 19366 4844 19394
rect 4632 18970 4660 19366
rect 4620 18964 4672 18970
rect 4620 18906 4672 18912
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4724 17882 4752 18838
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4816 16794 4844 17138
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4342 16079 4398 16088
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4172 14572 4292 14600
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 13326 3556 14486
rect 3608 14272 3660 14278
rect 4172 14260 4200 14572
rect 4250 14512 4306 14521
rect 4448 14482 4476 16050
rect 4540 14498 4568 16050
rect 4908 16046 4936 20839
rect 5000 18193 5028 23423
rect 5276 23118 5304 24074
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22098 5212 22374
rect 5262 22128 5318 22137
rect 5172 22092 5224 22098
rect 5262 22063 5318 22072
rect 5172 22034 5224 22040
rect 5276 22030 5304 22063
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 5092 21690 5120 21966
rect 5172 21956 5224 21962
rect 5172 21898 5224 21904
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5078 21176 5134 21185
rect 5078 21111 5134 21120
rect 5092 20806 5120 21111
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 5092 18850 5120 20742
rect 5184 20058 5212 21898
rect 5368 21468 5396 26182
rect 5538 26143 5594 26152
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 5460 24342 5488 24686
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 5460 23225 5488 23666
rect 5446 23216 5502 23225
rect 5446 23151 5502 23160
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5276 21440 5396 21468
rect 5276 20942 5304 21440
rect 5460 21400 5488 23054
rect 5368 21372 5488 21400
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5264 20528 5316 20534
rect 5264 20470 5316 20476
rect 5172 20052 5224 20058
rect 5172 19994 5224 20000
rect 5184 19394 5212 19994
rect 5276 19514 5304 20470
rect 5368 20346 5396 21372
rect 5552 21298 5580 26143
rect 5644 24426 5672 27288
rect 5736 24721 5764 29514
rect 5828 26246 5856 29514
rect 5816 26240 5868 26246
rect 5816 26182 5868 26188
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5722 24712 5778 24721
rect 5722 24647 5778 24656
rect 5724 24608 5776 24614
rect 5828 24596 5856 25638
rect 5776 24568 5856 24596
rect 5724 24550 5776 24556
rect 5644 24398 5764 24426
rect 5630 24304 5686 24313
rect 5630 24239 5686 24248
rect 5644 23254 5672 24239
rect 5736 23322 5764 24398
rect 5828 24342 5856 24568
rect 5816 24336 5868 24342
rect 5816 24278 5868 24284
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5632 23248 5684 23254
rect 5920 23202 5948 31470
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 6012 25974 6040 30874
rect 6104 29617 6132 31758
rect 6196 31210 6224 31758
rect 6288 31754 6316 32014
rect 6276 31748 6328 31754
rect 6276 31690 6328 31696
rect 6184 31204 6236 31210
rect 6184 31146 6236 31152
rect 6182 30968 6238 30977
rect 6182 30903 6238 30912
rect 6090 29608 6146 29617
rect 6090 29543 6146 29552
rect 6104 29073 6132 29543
rect 6090 29064 6146 29073
rect 6090 28999 6146 29008
rect 6090 27976 6146 27985
rect 6090 27911 6146 27920
rect 6000 25968 6052 25974
rect 6000 25910 6052 25916
rect 6104 24426 6132 27911
rect 6196 25888 6224 30903
rect 6288 30802 6316 31690
rect 6380 31686 6408 34002
rect 6472 31822 6500 35430
rect 6564 33590 6592 37402
rect 6644 36236 6696 36242
rect 6644 36178 6696 36184
rect 6656 35834 6684 36178
rect 6644 35828 6696 35834
rect 6644 35770 6696 35776
rect 6644 35148 6696 35154
rect 6644 35090 6696 35096
rect 6552 33584 6604 33590
rect 6552 33526 6604 33532
rect 6656 33454 6684 35090
rect 6748 34950 6776 39578
rect 6840 39506 6868 39766
rect 6828 39500 6880 39506
rect 6828 39442 6880 39448
rect 6884 39196 7192 39205
rect 6884 39194 6890 39196
rect 6946 39194 6970 39196
rect 7026 39194 7050 39196
rect 7106 39194 7130 39196
rect 7186 39194 7192 39196
rect 6946 39142 6948 39194
rect 7128 39142 7130 39194
rect 6884 39140 6890 39142
rect 6946 39140 6970 39142
rect 7026 39140 7050 39142
rect 7106 39140 7130 39142
rect 7186 39140 7192 39142
rect 6884 39131 7192 39140
rect 6828 38888 6880 38894
rect 6828 38830 6880 38836
rect 6840 38214 6868 38830
rect 6828 38208 6880 38214
rect 6828 38150 6880 38156
rect 6884 38108 7192 38117
rect 6884 38106 6890 38108
rect 6946 38106 6970 38108
rect 7026 38106 7050 38108
rect 7106 38106 7130 38108
rect 7186 38106 7192 38108
rect 6946 38054 6948 38106
rect 7128 38054 7130 38106
rect 6884 38052 6890 38054
rect 6946 38052 6970 38054
rect 7026 38052 7050 38054
rect 7106 38052 7130 38054
rect 7186 38052 7192 38054
rect 6884 38043 7192 38052
rect 6884 37020 7192 37029
rect 6884 37018 6890 37020
rect 6946 37018 6970 37020
rect 7026 37018 7050 37020
rect 7106 37018 7130 37020
rect 7186 37018 7192 37020
rect 6946 36966 6948 37018
rect 7128 36966 7130 37018
rect 6884 36964 6890 36966
rect 6946 36964 6970 36966
rect 7026 36964 7050 36966
rect 7106 36964 7130 36966
rect 7186 36964 7192 36966
rect 6884 36955 7192 36964
rect 6920 36780 6972 36786
rect 6920 36722 6972 36728
rect 7012 36780 7064 36786
rect 7012 36722 7064 36728
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 6932 36378 6960 36722
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 7024 36038 7052 36722
rect 7116 36174 7144 36722
rect 7104 36168 7156 36174
rect 7104 36110 7156 36116
rect 7012 36032 7064 36038
rect 7012 35974 7064 35980
rect 6884 35932 7192 35941
rect 6884 35930 6890 35932
rect 6946 35930 6970 35932
rect 7026 35930 7050 35932
rect 7106 35930 7130 35932
rect 7186 35930 7192 35932
rect 6946 35878 6948 35930
rect 7128 35878 7130 35930
rect 6884 35876 6890 35878
rect 6946 35876 6970 35878
rect 7026 35876 7050 35878
rect 7106 35876 7130 35878
rect 7186 35876 7192 35878
rect 6884 35867 7192 35876
rect 6736 34944 6788 34950
rect 6736 34886 6788 34892
rect 6748 33998 6776 34886
rect 6884 34844 7192 34853
rect 6884 34842 6890 34844
rect 6946 34842 6970 34844
rect 7026 34842 7050 34844
rect 7106 34842 7130 34844
rect 7186 34842 7192 34844
rect 6946 34790 6948 34842
rect 7128 34790 7130 34842
rect 6884 34788 6890 34790
rect 6946 34788 6970 34790
rect 7026 34788 7050 34790
rect 7106 34788 7130 34790
rect 7186 34788 7192 34790
rect 6884 34779 7192 34788
rect 6736 33992 6788 33998
rect 6736 33934 6788 33940
rect 6884 33756 7192 33765
rect 6884 33754 6890 33756
rect 6946 33754 6970 33756
rect 7026 33754 7050 33756
rect 7106 33754 7130 33756
rect 7186 33754 7192 33756
rect 6946 33702 6948 33754
rect 7128 33702 7130 33754
rect 6884 33700 6890 33702
rect 6946 33700 6970 33702
rect 7026 33700 7050 33702
rect 7106 33700 7130 33702
rect 7186 33700 7192 33702
rect 6884 33691 7192 33700
rect 6736 33584 6788 33590
rect 6736 33526 6788 33532
rect 6644 33448 6696 33454
rect 6644 33390 6696 33396
rect 6552 33312 6604 33318
rect 6552 33254 6604 33260
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6368 31680 6420 31686
rect 6368 31622 6420 31628
rect 6380 31414 6408 31622
rect 6368 31408 6420 31414
rect 6368 31350 6420 31356
rect 6460 31408 6512 31414
rect 6564 31396 6592 33254
rect 6656 32609 6684 33390
rect 6642 32600 6698 32609
rect 6642 32535 6698 32544
rect 6748 32314 6776 33526
rect 7012 33448 7064 33454
rect 6918 33416 6974 33425
rect 7196 33448 7248 33454
rect 7012 33390 7064 33396
rect 7194 33416 7196 33425
rect 7248 33416 7250 33425
rect 6918 33351 6974 33360
rect 6932 32910 6960 33351
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 7024 32842 7052 33390
rect 7194 33351 7250 33360
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 6884 32668 7192 32677
rect 6884 32666 6890 32668
rect 6946 32666 6970 32668
rect 7026 32666 7050 32668
rect 7106 32666 7130 32668
rect 7186 32666 7192 32668
rect 6946 32614 6948 32666
rect 7128 32614 7130 32666
rect 6884 32612 6890 32614
rect 6946 32612 6970 32614
rect 7026 32612 7050 32614
rect 7106 32612 7130 32614
rect 7186 32612 7192 32614
rect 6884 32603 7192 32612
rect 6748 32286 6868 32314
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6748 31958 6776 32166
rect 6736 31952 6788 31958
rect 6642 31920 6698 31929
rect 6736 31894 6788 31900
rect 6642 31855 6698 31864
rect 6512 31368 6592 31396
rect 6460 31350 6512 31356
rect 6276 30796 6328 30802
rect 6276 30738 6328 30744
rect 6288 30054 6316 30738
rect 6472 30326 6500 31350
rect 6552 31136 6604 31142
rect 6552 31078 6604 31084
rect 6460 30320 6512 30326
rect 6460 30262 6512 30268
rect 6460 30184 6512 30190
rect 6460 30126 6512 30132
rect 6276 30048 6328 30054
rect 6276 29990 6328 29996
rect 6288 28014 6316 29990
rect 6472 29481 6500 30126
rect 6458 29472 6514 29481
rect 6458 29407 6514 29416
rect 6472 29170 6500 29407
rect 6460 29164 6512 29170
rect 6460 29106 6512 29112
rect 6564 28994 6592 31078
rect 6472 28966 6592 28994
rect 6276 28008 6328 28014
rect 6276 27950 6328 27956
rect 6288 27334 6316 27950
rect 6368 27668 6420 27674
rect 6368 27610 6420 27616
rect 6380 27334 6408 27610
rect 6472 27334 6500 28966
rect 6552 28416 6604 28422
rect 6552 28358 6604 28364
rect 6564 27470 6592 28358
rect 6552 27464 6604 27470
rect 6552 27406 6604 27412
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 6276 25900 6328 25906
rect 6196 25860 6276 25888
rect 6276 25842 6328 25848
rect 6184 25356 6236 25362
rect 6184 25298 6236 25304
rect 5632 23190 5684 23196
rect 5736 23174 5948 23202
rect 6012 24398 6132 24426
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5644 21962 5672 22714
rect 5632 21956 5684 21962
rect 5632 21898 5684 21904
rect 5736 21672 5764 23174
rect 6012 23066 6040 24398
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6104 23798 6132 24142
rect 6092 23792 6144 23798
rect 6092 23734 6144 23740
rect 5644 21644 5764 21672
rect 5828 23038 6040 23066
rect 5644 21418 5672 21644
rect 5632 21412 5684 21418
rect 5632 21354 5684 21360
rect 5552 21270 5672 21298
rect 5368 20318 5488 20346
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5264 19508 5316 19514
rect 5264 19450 5316 19456
rect 5368 19394 5396 19790
rect 5184 19366 5396 19394
rect 5460 19334 5488 20318
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5552 19514 5580 19722
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5460 19306 5580 19334
rect 5354 19272 5410 19281
rect 5410 19230 5488 19258
rect 5354 19207 5410 19216
rect 5356 19168 5408 19174
rect 5354 19136 5356 19145
rect 5408 19136 5410 19145
rect 5354 19071 5410 19080
rect 5092 18822 5304 18850
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17678 5028 18022
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5184 16969 5212 18226
rect 5170 16960 5226 16969
rect 5170 16895 5226 16904
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 15706 4660 15846
rect 4724 15706 4752 15982
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4618 15192 4674 15201
rect 4618 15127 4620 15136
rect 4672 15127 4674 15136
rect 4620 15098 4672 15104
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4250 14447 4306 14456
rect 4436 14476 4488 14482
rect 4264 14414 4292 14447
rect 4540 14470 4752 14498
rect 4436 14418 4488 14424
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4344 14272 4396 14278
rect 4172 14232 4292 14260
rect 3608 14214 3660 14220
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3514 13016 3570 13025
rect 3514 12951 3570 12960
rect 3528 12442 3556 12951
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11898 3556 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3514 11792 3570 11801
rect 3514 11727 3516 11736
rect 3568 11727 3570 11736
rect 3516 11698 3568 11704
rect 3620 11529 3648 14214
rect 3700 13932 3752 13938
rect 3700 13874 3752 13880
rect 3712 12424 3740 13874
rect 3792 13728 3844 13734
rect 3790 13696 3792 13705
rect 3844 13696 3846 13705
rect 3790 13631 3846 13640
rect 3917 13628 4225 13637
rect 3917 13626 3923 13628
rect 3979 13626 4003 13628
rect 4059 13626 4083 13628
rect 4139 13626 4163 13628
rect 4219 13626 4225 13628
rect 3979 13574 3981 13626
rect 4161 13574 4163 13626
rect 3917 13572 3923 13574
rect 3979 13572 4003 13574
rect 4059 13572 4083 13574
rect 4139 13572 4163 13574
rect 4219 13572 4225 13574
rect 3917 13563 4225 13572
rect 3790 13424 3846 13433
rect 3790 13359 3792 13368
rect 3844 13359 3846 13368
rect 3792 13330 3844 13336
rect 4068 13320 4120 13326
rect 4066 13288 4068 13297
rect 4120 13288 4122 13297
rect 4066 13223 4122 13232
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12986 3832 13126
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3884 12912 3936 12918
rect 3882 12880 3884 12889
rect 3936 12880 3938 12889
rect 3882 12815 3938 12824
rect 4068 12776 4120 12782
rect 4066 12744 4068 12753
rect 4120 12744 4122 12753
rect 4066 12679 4122 12688
rect 3917 12540 4225 12549
rect 3917 12538 3923 12540
rect 3979 12538 4003 12540
rect 4059 12538 4083 12540
rect 4139 12538 4163 12540
rect 4219 12538 4225 12540
rect 3979 12486 3981 12538
rect 4161 12486 4163 12538
rect 3917 12484 3923 12486
rect 3979 12484 4003 12486
rect 4059 12484 4083 12486
rect 4139 12484 4163 12486
rect 4219 12484 4225 12486
rect 3917 12475 4225 12484
rect 4264 12434 4292 14232
rect 4344 14214 4396 14220
rect 4356 13938 4384 14214
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4448 13326 4476 14418
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 3712 12396 3832 12424
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3712 12102 3740 12271
rect 3700 12096 3752 12102
rect 3700 12038 3752 12044
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3606 11520 3662 11529
rect 3606 11455 3662 11464
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3620 11257 3648 11290
rect 3606 11248 3662 11257
rect 3606 11183 3662 11192
rect 3436 11104 3648 11132
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3330 10432 3386 10441
rect 3330 10367 3386 10376
rect 3344 9722 3372 10367
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3436 9654 3464 10950
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 10130 3556 10474
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3424 9648 3476 9654
rect 3330 9616 3386 9625
rect 3240 9580 3292 9586
rect 3424 9590 3476 9596
rect 3516 9648 3568 9654
rect 3516 9590 3568 9596
rect 3330 9551 3386 9560
rect 3240 9522 3292 9528
rect 3160 8588 3280 8616
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2870 5199 2926 5208
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3528 2740 3534
rect 2686 3496 2688 3505
rect 2780 3528 2832 3534
rect 2740 3496 2742 3505
rect 2780 3470 2832 3476
rect 2686 3431 2742 3440
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2608 2446 2636 3334
rect 2792 3058 2820 3470
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2976 2650 3004 4558
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2688 2372 2740 2378
rect 2688 2314 2740 2320
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 1952 1352 2004 1358
rect 1952 1294 2004 1300
rect 2044 1352 2096 1358
rect 2044 1294 2096 1300
rect 1412 746 1440 1294
rect 1768 1284 1820 1290
rect 1768 1226 1820 1232
rect 1400 740 1452 746
rect 1400 682 1452 688
rect 754 54 888 82
rect 754 0 810 54
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 82 1638 160
rect 1780 82 1808 1226
rect 1582 54 1808 82
rect 1858 82 1914 160
rect 2056 82 2084 1294
rect 2320 1284 2372 1290
rect 2320 1226 2372 1232
rect 1858 54 2084 82
rect 2134 82 2190 160
rect 2332 82 2360 1226
rect 2412 740 2464 746
rect 2412 682 2464 688
rect 2424 160 2452 682
rect 2700 160 2728 2314
rect 3068 1766 3096 2926
rect 3160 2854 3188 8434
rect 3252 6390 3280 8588
rect 3344 8480 3372 9551
rect 3528 9518 3556 9590
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3344 8452 3464 8480
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3344 7993 3372 8298
rect 3330 7984 3386 7993
rect 3330 7919 3386 7928
rect 3436 7410 3464 8452
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3528 7290 3556 9454
rect 3620 8974 3648 11104
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3712 8650 3740 11834
rect 3804 9178 3832 12396
rect 4172 12406 4292 12434
rect 3882 12200 3938 12209
rect 3882 12135 3938 12144
rect 3896 11762 3924 12135
rect 4172 12073 4200 12406
rect 4250 12336 4306 12345
rect 4250 12271 4306 12280
rect 4158 12064 4214 12073
rect 4158 11999 4214 12008
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3917 11452 4225 11461
rect 3917 11450 3923 11452
rect 3979 11450 4003 11452
rect 4059 11450 4083 11452
rect 4139 11450 4163 11452
rect 4219 11450 4225 11452
rect 3979 11398 3981 11450
rect 4161 11398 4163 11450
rect 3917 11396 3923 11398
rect 3979 11396 4003 11398
rect 4059 11396 4083 11398
rect 4139 11396 4163 11398
rect 4219 11396 4225 11398
rect 3917 11387 4225 11396
rect 4264 11200 4292 12271
rect 4356 12238 4384 12922
rect 4448 12782 4476 13126
rect 4632 12900 4660 14350
rect 4540 12872 4660 12900
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4540 12434 4568 12872
rect 4724 12850 4752 14470
rect 4816 14414 4844 14758
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4908 14226 4936 15982
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 5000 14346 5028 14962
rect 5080 14884 5132 14890
rect 5080 14826 5132 14832
rect 5092 14618 5120 14826
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 4908 14198 5028 14226
rect 4802 13424 4858 13433
rect 4802 13359 4858 13368
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4448 12406 4568 12434
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4264 11172 4384 11200
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3988 10713 4016 10950
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 4068 10600 4120 10606
rect 4066 10568 4068 10577
rect 4120 10568 4122 10577
rect 4066 10503 4122 10512
rect 3917 10364 4225 10373
rect 3917 10362 3923 10364
rect 3979 10362 4003 10364
rect 4059 10362 4083 10364
rect 4139 10362 4163 10364
rect 4219 10362 4225 10364
rect 3979 10310 3981 10362
rect 4161 10310 4163 10362
rect 3917 10308 3923 10310
rect 3979 10308 4003 10310
rect 4059 10308 4083 10310
rect 4139 10308 4163 10310
rect 4219 10308 4225 10310
rect 3917 10299 4225 10308
rect 3974 10160 4030 10169
rect 3896 10118 3974 10146
rect 3896 9654 3924 10118
rect 3974 10095 4030 10104
rect 3976 10056 4028 10062
rect 3974 10024 3976 10033
rect 4028 10024 4030 10033
rect 3974 9959 4030 9968
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 4264 9382 4292 11018
rect 4356 10130 4384 11172
rect 4448 10826 4476 12406
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4540 11014 4568 12174
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4448 10798 4568 10826
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4448 9722 4476 10066
rect 4436 9716 4488 9722
rect 4436 9658 4488 9664
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 3917 9276 4225 9285
rect 3917 9274 3923 9276
rect 3979 9274 4003 9276
rect 4059 9274 4083 9276
rect 4139 9274 4163 9276
rect 4219 9274 4225 9276
rect 3979 9222 3981 9274
rect 4161 9222 4163 9274
rect 3917 9220 3923 9222
rect 3979 9220 4003 9222
rect 4059 9220 4083 9222
rect 4139 9220 4163 9222
rect 4219 9220 4225 9222
rect 3917 9211 4225 9220
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3712 8622 3832 8650
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3344 7262 3556 7290
rect 3240 6384 3292 6390
rect 3238 6352 3240 6361
rect 3292 6352 3294 6361
rect 3238 6287 3294 6296
rect 3344 5846 3372 7262
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 3424 6724 3476 6730
rect 3424 6666 3476 6672
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3344 4146 3372 5306
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3330 4040 3386 4049
rect 3330 3975 3386 3984
rect 3344 3194 3372 3975
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3056 1760 3108 1766
rect 3056 1702 3108 1708
rect 3056 1352 3108 1358
rect 3056 1294 3108 1300
rect 2780 1216 2832 1222
rect 2780 1158 2832 1164
rect 2792 1018 2820 1158
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 2134 54 2360 82
rect 1582 0 1638 54
rect 1858 0 1914 54
rect 2134 0 2190 54
rect 2410 0 2466 160
rect 2686 0 2742 160
rect 2962 82 3018 160
rect 3068 82 3096 1294
rect 3252 160 3280 1906
rect 3344 1562 3372 2994
rect 3436 2922 3464 6666
rect 3528 6440 3556 7103
rect 3620 7002 3648 7346
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3712 6662 3740 8434
rect 3804 7954 3832 8622
rect 3917 8188 4225 8197
rect 3917 8186 3923 8188
rect 3979 8186 4003 8188
rect 4059 8186 4083 8188
rect 4139 8186 4163 8188
rect 4219 8186 4225 8188
rect 3979 8134 3981 8186
rect 4161 8134 4163 8186
rect 3917 8132 3923 8134
rect 3979 8132 4003 8134
rect 4059 8132 4083 8134
rect 4139 8132 4163 8134
rect 4219 8132 4225 8134
rect 3917 8123 4225 8132
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3884 7744 3936 7750
rect 3804 7704 3884 7732
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6452 3660 6458
rect 3528 6412 3608 6440
rect 3804 6440 3832 7704
rect 3884 7686 3936 7692
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3917 7100 4225 7109
rect 3917 7098 3923 7100
rect 3979 7098 4003 7100
rect 4059 7098 4083 7100
rect 4139 7098 4163 7100
rect 4219 7098 4225 7100
rect 3979 7046 3981 7098
rect 4161 7046 4163 7098
rect 3917 7044 3923 7046
rect 3979 7044 4003 7046
rect 4059 7044 4083 7046
rect 4139 7044 4163 7046
rect 4219 7044 4225 7046
rect 3917 7035 4225 7044
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4250 6896 4306 6905
rect 3608 6394 3660 6400
rect 3712 6412 3832 6440
rect 3712 5778 3740 6412
rect 4172 6322 4200 6870
rect 4250 6831 4306 6840
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3528 4146 3556 4626
rect 3620 4146 3648 4966
rect 3804 4758 3832 6258
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3896 5710 3924 5850
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 4080 5098 4108 5743
rect 4264 5710 4292 6831
rect 4356 6322 4384 9522
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4448 7342 4476 7890
rect 4540 7342 4568 10798
rect 4632 7342 4660 12718
rect 4816 12594 4844 13359
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4724 12566 4844 12594
rect 4724 11801 4752 12566
rect 4802 12472 4858 12481
rect 4802 12407 4858 12416
rect 4710 11792 4766 11801
rect 4710 11727 4766 11736
rect 4724 11694 4752 11727
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4724 10810 4752 11630
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4724 9518 4752 10746
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 8022 4752 9454
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4160 5704 4212 5710
rect 4160 5646 4212 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4172 5556 4200 5646
rect 4172 5528 4292 5556
rect 4068 5092 4120 5098
rect 4068 5034 4120 5040
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3976 4616 4028 4622
rect 3974 4584 3976 4593
rect 4028 4584 4030 4593
rect 4264 4570 4292 5528
rect 4448 5234 4476 7278
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4540 5166 4568 7278
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4724 5846 4752 6394
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4356 4690 4384 5034
rect 4540 5001 4568 5102
rect 4526 4992 4582 5001
rect 4526 4927 4582 4936
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4816 4622 4844 12407
rect 4908 11898 4936 12786
rect 5000 12434 5028 14198
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5092 12617 5120 13874
rect 5078 12608 5134 12617
rect 5078 12543 5134 12552
rect 5000 12406 5120 12434
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5000 10554 5028 12310
rect 4908 10526 5028 10554
rect 4908 10130 4936 10526
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 5000 10130 5028 10406
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5092 9586 5120 12406
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4894 8392 4950 8401
rect 4894 8327 4950 8336
rect 4908 7886 4936 8327
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 4908 7546 4936 7822
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4908 7002 4936 7482
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 5000 6458 5028 7210
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4894 5264 4950 5273
rect 4894 5199 4950 5208
rect 4908 5166 4936 5199
rect 5000 5166 5028 5510
rect 5092 5166 5120 7278
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4804 4616 4856 4622
rect 4264 4554 4384 4570
rect 4804 4558 4856 4564
rect 4264 4548 4396 4554
rect 4264 4542 4344 4548
rect 3974 4519 4030 4528
rect 4344 4490 4396 4496
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3712 3602 3740 4422
rect 4434 4312 4490 4321
rect 4434 4247 4490 4256
rect 4712 4276 4764 4282
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 3700 3596 3752 3602
rect 3700 3538 3752 3544
rect 4068 2984 4120 2990
rect 4066 2952 4068 2961
rect 4120 2952 4122 2961
rect 3424 2916 3476 2922
rect 4066 2887 4122 2896
rect 3424 2858 3476 2864
rect 4448 2774 4476 4247
rect 4712 4218 4764 4224
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 3194 4568 3334
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 4448 2746 4568 2774
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 3700 1964 3752 1970
rect 3700 1906 3752 1912
rect 3332 1556 3384 1562
rect 3332 1498 3384 1504
rect 3424 1216 3476 1222
rect 3424 1158 3476 1164
rect 3436 1018 3464 1158
rect 3424 1012 3476 1018
rect 3424 954 3476 960
rect 2962 54 3096 82
rect 2962 0 3018 54
rect 3238 0 3294 160
rect 3514 82 3570 160
rect 3712 82 3740 1906
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3804 1442 3832 1838
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 3804 1414 3924 1442
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3804 160 3832 1294
rect 3514 54 3740 82
rect 3514 0 3570 54
rect 3790 0 3846 160
rect 3896 82 3924 1414
rect 4068 1352 4120 1358
rect 3974 1320 4030 1329
rect 4068 1294 4120 1300
rect 3974 1255 4030 1264
rect 3988 1222 4016 1255
rect 3976 1216 4028 1222
rect 4080 1193 4108 1294
rect 3976 1158 4028 1164
rect 4066 1184 4122 1193
rect 4066 1119 4122 1128
rect 4066 82 4122 160
rect 3896 54 4122 82
rect 4066 0 4122 54
rect 4342 82 4398 160
rect 4448 82 4476 2382
rect 4540 2106 4568 2746
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4632 1902 4660 3470
rect 4724 1970 4752 4218
rect 5078 3768 5134 3777
rect 5078 3703 5134 3712
rect 5092 3670 5120 3703
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4896 3392 4948 3398
rect 4894 3360 4896 3369
rect 4948 3360 4950 3369
rect 4894 3295 4950 3304
rect 5184 2774 5212 16895
rect 5276 13938 5304 18822
rect 5368 18465 5396 19071
rect 5354 18456 5410 18465
rect 5354 18391 5410 18400
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17746 5396 18022
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5368 15502 5396 17206
rect 5460 15978 5488 19230
rect 5552 16454 5580 19306
rect 5540 16448 5592 16454
rect 5540 16390 5592 16396
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 15570 5488 15914
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14550 5396 14758
rect 5644 14657 5672 21270
rect 5828 20346 5856 23038
rect 6196 22642 6224 25298
rect 6288 24886 6316 25842
rect 6368 25152 6420 25158
rect 6368 25094 6420 25100
rect 6276 24880 6328 24886
rect 6276 24822 6328 24828
rect 6380 24750 6408 25094
rect 6368 24744 6420 24750
rect 6368 24686 6420 24692
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6184 22636 6236 22642
rect 6184 22578 6236 22584
rect 6196 22166 6224 22578
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6182 21856 6238 21865
rect 5908 21412 5960 21418
rect 5908 21354 5960 21360
rect 5920 21162 5948 21354
rect 6012 21350 6040 21830
rect 6182 21791 6238 21800
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 6104 21457 6132 21626
rect 6090 21448 6146 21457
rect 6090 21383 6146 21392
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5920 21134 6040 21162
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5736 20318 5856 20346
rect 5630 14648 5686 14657
rect 5630 14583 5686 14592
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5448 14476 5500 14482
rect 5736 14464 5764 20318
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5828 19922 5856 20198
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5920 19854 5948 20946
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 6012 19281 6040 21134
rect 5998 19272 6054 19281
rect 5998 19207 6054 19216
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5828 18358 5856 18702
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5828 17678 5856 18294
rect 6000 17808 6052 17814
rect 5998 17776 6000 17785
rect 6052 17776 6054 17785
rect 5998 17711 6054 17720
rect 5816 17672 5868 17678
rect 5816 17614 5868 17620
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5828 14793 5856 17478
rect 5920 17202 5948 17546
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5814 14784 5870 14793
rect 5814 14719 5870 14728
rect 5920 14618 5948 14826
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 5448 14418 5500 14424
rect 5552 14436 5764 14464
rect 5908 14476 5960 14482
rect 5354 14376 5410 14385
rect 5354 14311 5410 14320
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5276 12238 5304 13126
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5262 11792 5318 11801
rect 5262 11727 5264 11736
rect 5316 11727 5318 11736
rect 5264 11698 5316 11704
rect 5276 11234 5304 11698
rect 5368 11558 5396 14311
rect 5460 14113 5488 14418
rect 5446 14104 5502 14113
rect 5446 14039 5502 14048
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12306 5488 13262
rect 5552 12986 5580 14436
rect 5908 14418 5960 14424
rect 5816 14408 5868 14414
rect 5644 14368 5816 14396
rect 5644 13977 5672 14368
rect 5816 14350 5868 14356
rect 5920 14113 5948 14418
rect 5906 14104 5962 14113
rect 5906 14039 5962 14048
rect 5630 13968 5686 13977
rect 5630 13903 5686 13912
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5446 11248 5502 11257
rect 5276 11206 5446 11234
rect 5446 11183 5502 11192
rect 5356 11008 5408 11014
rect 5356 10950 5408 10956
rect 5368 10130 5396 10950
rect 5540 10192 5592 10198
rect 5644 10180 5672 13903
rect 5906 13560 5962 13569
rect 5906 13495 5962 13504
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5828 12288 5856 12922
rect 5920 12594 5948 13495
rect 6012 12986 6040 16662
rect 6196 16538 6224 21791
rect 6288 17116 6316 24550
rect 6380 24274 6408 24686
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6368 23792 6420 23798
rect 6368 23734 6420 23740
rect 6380 21622 6408 23734
rect 6472 23168 6500 27270
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6564 25362 6592 26386
rect 6552 25356 6604 25362
rect 6552 25298 6604 25304
rect 6552 24676 6604 24682
rect 6552 24618 6604 24624
rect 6564 23526 6592 24618
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6472 23140 6592 23168
rect 6458 23080 6514 23089
rect 6458 23015 6514 23024
rect 6368 21616 6420 21622
rect 6368 21558 6420 21564
rect 6380 18329 6408 21558
rect 6366 18320 6422 18329
rect 6366 18255 6422 18264
rect 6380 17338 6408 18255
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6472 17270 6500 23015
rect 6564 22778 6592 23140
rect 6656 22982 6684 31855
rect 6736 31680 6788 31686
rect 6840 31668 6868 32286
rect 7102 31920 7158 31929
rect 7102 31855 7158 31864
rect 6736 31622 6788 31628
rect 6822 31640 6868 31668
rect 7116 31668 7144 31855
rect 7300 31754 7328 41414
rect 7852 41274 7880 42094
rect 7944 41721 7972 42162
rect 8024 42016 8076 42022
rect 8024 41958 8076 41964
rect 7930 41712 7986 41721
rect 7930 41647 7986 41656
rect 8036 41414 8064 41958
rect 8128 41750 8156 43250
rect 8220 42362 8248 44463
rect 8496 43450 8524 44463
rect 8484 43444 8536 43450
rect 8484 43386 8536 43392
rect 8576 43376 8628 43382
rect 8576 43318 8628 43324
rect 8390 42800 8446 42809
rect 8390 42735 8446 42744
rect 8484 42764 8536 42770
rect 8404 42702 8432 42735
rect 8484 42706 8536 42712
rect 8392 42696 8444 42702
rect 8392 42638 8444 42644
rect 8208 42356 8260 42362
rect 8208 42298 8260 42304
rect 8208 42220 8260 42226
rect 8208 42162 8260 42168
rect 8116 41744 8168 41750
rect 8116 41686 8168 41692
rect 7944 41386 8064 41414
rect 7840 41268 7892 41274
rect 7840 41210 7892 41216
rect 7944 41138 7972 41386
rect 7932 41132 7984 41138
rect 7932 41074 7984 41080
rect 7656 40724 7708 40730
rect 7656 40666 7708 40672
rect 7668 40610 7696 40666
rect 7576 40582 7696 40610
rect 7470 40216 7526 40225
rect 7470 40151 7472 40160
rect 7524 40151 7526 40160
rect 7472 40122 7524 40128
rect 7576 40118 7604 40582
rect 7656 40520 7708 40526
rect 7656 40462 7708 40468
rect 7564 40112 7616 40118
rect 7564 40054 7616 40060
rect 7380 39500 7432 39506
rect 7380 39442 7432 39448
rect 7392 38962 7420 39442
rect 7576 39438 7604 40054
rect 7668 40050 7696 40462
rect 7932 40384 7984 40390
rect 7932 40326 7984 40332
rect 7656 40044 7708 40050
rect 7656 39986 7708 39992
rect 7944 39982 7972 40326
rect 8024 40180 8076 40186
rect 8024 40122 8076 40128
rect 8036 40050 8064 40122
rect 8024 40044 8076 40050
rect 8024 39986 8076 39992
rect 8116 40044 8168 40050
rect 8116 39986 8168 39992
rect 7932 39976 7984 39982
rect 7932 39918 7984 39924
rect 7564 39432 7616 39438
rect 7564 39374 7616 39380
rect 7380 38956 7432 38962
rect 7380 38898 7432 38904
rect 7472 38208 7524 38214
rect 7472 38150 7524 38156
rect 7380 37664 7432 37670
rect 7380 37606 7432 37612
rect 7392 37398 7420 37606
rect 7380 37392 7432 37398
rect 7380 37334 7432 37340
rect 7484 36854 7512 38150
rect 7576 37874 7604 39374
rect 8024 39364 8076 39370
rect 8024 39306 8076 39312
rect 8036 39098 8064 39306
rect 8024 39092 8076 39098
rect 8024 39034 8076 39040
rect 7656 38344 7708 38350
rect 7656 38286 7708 38292
rect 7564 37868 7616 37874
rect 7564 37810 7616 37816
rect 7472 36848 7524 36854
rect 7472 36790 7524 36796
rect 7472 36712 7524 36718
rect 7472 36654 7524 36660
rect 7484 36242 7512 36654
rect 7472 36236 7524 36242
rect 7472 36178 7524 36184
rect 7380 36168 7432 36174
rect 7378 36136 7380 36145
rect 7432 36136 7434 36145
rect 7378 36071 7434 36080
rect 7380 36032 7432 36038
rect 7380 35974 7432 35980
rect 7392 35222 7420 35974
rect 7380 35216 7432 35222
rect 7380 35158 7432 35164
rect 7380 34400 7432 34406
rect 7380 34342 7432 34348
rect 7472 34400 7524 34406
rect 7472 34342 7524 34348
rect 7392 34134 7420 34342
rect 7380 34128 7432 34134
rect 7380 34070 7432 34076
rect 7392 33386 7420 34070
rect 7380 33380 7432 33386
rect 7380 33322 7432 33328
rect 7484 31754 7512 34342
rect 7576 32570 7604 37810
rect 7668 35290 7696 38286
rect 7932 38276 7984 38282
rect 7932 38218 7984 38224
rect 7840 37936 7892 37942
rect 7840 37878 7892 37884
rect 7746 36816 7802 36825
rect 7746 36751 7748 36760
rect 7800 36751 7802 36760
rect 7748 36722 7800 36728
rect 7852 36378 7880 37878
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7656 35284 7708 35290
rect 7656 35226 7708 35232
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7564 32564 7616 32570
rect 7564 32506 7616 32512
rect 7668 31890 7696 34342
rect 7760 32774 7788 35974
rect 7840 35488 7892 35494
rect 7840 35430 7892 35436
rect 7852 35290 7880 35430
rect 7840 35284 7892 35290
rect 7840 35226 7892 35232
rect 7838 34912 7894 34921
rect 7838 34847 7894 34856
rect 7852 33862 7880 34847
rect 7840 33856 7892 33862
rect 7840 33798 7892 33804
rect 7838 33688 7894 33697
rect 7838 33623 7894 33632
rect 7748 32768 7800 32774
rect 7748 32710 7800 32716
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7656 31884 7708 31890
rect 7656 31826 7708 31832
rect 7300 31726 7420 31754
rect 7116 31640 7328 31668
rect 6748 31278 6776 31622
rect 6822 31464 6850 31640
rect 6884 31580 7192 31589
rect 6884 31578 6890 31580
rect 6946 31578 6970 31580
rect 7026 31578 7050 31580
rect 7106 31578 7130 31580
rect 7186 31578 7192 31580
rect 6946 31526 6948 31578
rect 7128 31526 7130 31578
rect 6884 31524 6890 31526
rect 6946 31524 6970 31526
rect 7026 31524 7050 31526
rect 7106 31524 7130 31526
rect 7186 31524 7192 31526
rect 6884 31515 7192 31524
rect 7196 31476 7248 31482
rect 6822 31436 6868 31464
rect 6736 31272 6788 31278
rect 6736 31214 6788 31220
rect 6840 30666 6868 31436
rect 7196 31418 7248 31424
rect 7208 30938 7236 31418
rect 7300 31346 7328 31640
rect 7288 31340 7340 31346
rect 7288 31282 7340 31288
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 6828 30660 6880 30666
rect 6748 30620 6828 30648
rect 6748 29345 6776 30620
rect 6828 30602 6880 30608
rect 6884 30492 7192 30501
rect 6884 30490 6890 30492
rect 6946 30490 6970 30492
rect 7026 30490 7050 30492
rect 7106 30490 7130 30492
rect 7186 30490 7192 30492
rect 6946 30438 6948 30490
rect 7128 30438 7130 30490
rect 6884 30436 6890 30438
rect 6946 30436 6970 30438
rect 7026 30436 7050 30438
rect 7106 30436 7130 30438
rect 7186 30436 7192 30438
rect 6884 30427 7192 30436
rect 7196 30252 7248 30258
rect 7248 30212 7328 30240
rect 7196 30194 7248 30200
rect 7104 29640 7156 29646
rect 7102 29608 7104 29617
rect 7156 29608 7158 29617
rect 7102 29543 7158 29552
rect 6884 29404 7192 29413
rect 6884 29402 6890 29404
rect 6946 29402 6970 29404
rect 7026 29402 7050 29404
rect 7106 29402 7130 29404
rect 7186 29402 7192 29404
rect 6946 29350 6948 29402
rect 7128 29350 7130 29402
rect 6884 29348 6890 29350
rect 6946 29348 6970 29350
rect 7026 29348 7050 29350
rect 7106 29348 7130 29350
rect 7186 29348 7192 29350
rect 6734 29336 6790 29345
rect 6884 29339 7192 29348
rect 6734 29271 6790 29280
rect 6748 28098 6776 29271
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7102 29064 7158 29073
rect 7102 28999 7104 29008
rect 7156 28999 7158 29008
rect 7104 28970 7156 28976
rect 7208 28558 7236 29106
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7300 28422 7328 30212
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 6884 28316 7192 28325
rect 6884 28314 6890 28316
rect 6946 28314 6970 28316
rect 7026 28314 7050 28316
rect 7106 28314 7130 28316
rect 7186 28314 7192 28316
rect 6946 28262 6948 28314
rect 7128 28262 7130 28314
rect 6884 28260 6890 28262
rect 6946 28260 6970 28262
rect 7026 28260 7050 28262
rect 7106 28260 7130 28262
rect 7186 28260 7192 28262
rect 6884 28251 7192 28260
rect 6826 28112 6882 28121
rect 6748 28070 6826 28098
rect 6826 28047 6882 28056
rect 7196 28008 7248 28014
rect 7196 27950 7248 27956
rect 6828 27872 6880 27878
rect 7208 27849 7236 27950
rect 7300 27946 7328 28358
rect 7288 27940 7340 27946
rect 7288 27882 7340 27888
rect 6828 27814 6880 27820
rect 7194 27840 7250 27849
rect 6840 27470 6868 27814
rect 7194 27775 7250 27784
rect 7102 27568 7158 27577
rect 7102 27503 7158 27512
rect 7116 27470 7144 27503
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6828 27328 6880 27334
rect 6748 27305 6828 27316
rect 6734 27296 6828 27305
rect 6790 27288 6828 27296
rect 6828 27270 6880 27276
rect 6734 27231 6790 27240
rect 6884 27228 7192 27237
rect 6884 27226 6890 27228
rect 6946 27226 6970 27228
rect 7026 27226 7050 27228
rect 7106 27226 7130 27228
rect 7186 27226 7192 27228
rect 6946 27174 6948 27226
rect 7128 27174 7130 27226
rect 6884 27172 6890 27174
rect 6946 27172 6970 27174
rect 7026 27172 7050 27174
rect 7106 27172 7130 27174
rect 7186 27172 7192 27174
rect 6884 27163 7192 27172
rect 7286 26888 7342 26897
rect 7286 26823 7342 26832
rect 6734 26480 6790 26489
rect 6734 26415 6790 26424
rect 6748 26382 6776 26415
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6552 22772 6604 22778
rect 6552 22714 6604 22720
rect 6748 22658 6776 26318
rect 6884 26140 7192 26149
rect 6884 26138 6890 26140
rect 6946 26138 6970 26140
rect 7026 26138 7050 26140
rect 7106 26138 7130 26140
rect 7186 26138 7192 26140
rect 6946 26086 6948 26138
rect 7128 26086 7130 26138
rect 6884 26084 6890 26086
rect 6946 26084 6970 26086
rect 7026 26084 7050 26086
rect 7106 26084 7130 26086
rect 7186 26084 7192 26086
rect 6884 26075 7192 26084
rect 7300 25974 7328 26823
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 6826 25528 6882 25537
rect 6826 25463 6882 25472
rect 6840 25265 6868 25463
rect 7012 25288 7064 25294
rect 6826 25256 6882 25265
rect 6826 25191 6882 25200
rect 7010 25256 7012 25265
rect 7064 25256 7066 25265
rect 7010 25191 7066 25200
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 6884 25052 7192 25061
rect 6884 25050 6890 25052
rect 6946 25050 6970 25052
rect 7026 25050 7050 25052
rect 7106 25050 7130 25052
rect 7186 25050 7192 25052
rect 6946 24998 6948 25050
rect 7128 24998 7130 25050
rect 6884 24996 6890 24998
rect 6946 24996 6970 24998
rect 7026 24996 7050 24998
rect 7106 24996 7130 24998
rect 7186 24996 7192 24998
rect 6884 24987 7192 24996
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 6932 24410 6960 24754
rect 6920 24404 6972 24410
rect 6920 24346 6972 24352
rect 6884 23964 7192 23973
rect 6884 23962 6890 23964
rect 6946 23962 6970 23964
rect 7026 23962 7050 23964
rect 7106 23962 7130 23964
rect 7186 23962 7192 23964
rect 6946 23910 6948 23962
rect 7128 23910 7130 23962
rect 6884 23908 6890 23910
rect 6946 23908 6970 23910
rect 7026 23908 7050 23910
rect 7106 23908 7130 23910
rect 7186 23908 7192 23910
rect 6884 23899 7192 23908
rect 7300 23798 7328 25094
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 6884 22876 7192 22885
rect 6884 22874 6890 22876
rect 6946 22874 6970 22876
rect 7026 22874 7050 22876
rect 7106 22874 7130 22876
rect 7186 22874 7192 22876
rect 6946 22822 6948 22874
rect 7128 22822 7130 22874
rect 6884 22820 6890 22822
rect 6946 22820 6970 22822
rect 7026 22820 7050 22822
rect 7106 22820 7130 22822
rect 7186 22820 7192 22822
rect 6884 22811 7192 22820
rect 6748 22630 6868 22658
rect 6736 22432 6788 22438
rect 6736 22374 6788 22380
rect 6552 22160 6604 22166
rect 6604 22108 6684 22114
rect 6552 22102 6684 22108
rect 6564 22086 6684 22102
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 20466 6592 21966
rect 6656 21622 6684 22086
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 6748 21486 6776 22374
rect 6840 22137 6868 22630
rect 7300 22506 7328 23734
rect 7288 22500 7340 22506
rect 7288 22442 7340 22448
rect 6826 22128 6882 22137
rect 6826 22063 6882 22072
rect 7392 21978 7420 31726
rect 7472 31748 7524 31754
rect 7472 31690 7524 31696
rect 7564 31476 7616 31482
rect 7564 31418 7616 31424
rect 7472 31408 7524 31414
rect 7472 31350 7524 31356
rect 7484 28529 7512 31350
rect 7576 29560 7604 31418
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7668 29714 7696 30126
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7576 29532 7696 29560
rect 7562 29472 7618 29481
rect 7562 29407 7618 29416
rect 7470 28520 7526 28529
rect 7470 28455 7526 28464
rect 7470 28248 7526 28257
rect 7470 28183 7526 28192
rect 7484 27441 7512 28183
rect 7470 27432 7526 27441
rect 7470 27367 7526 27376
rect 7472 27328 7524 27334
rect 7472 27270 7524 27276
rect 7484 27033 7512 27270
rect 7470 27024 7526 27033
rect 7470 26959 7526 26968
rect 7484 26382 7512 26959
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7576 26228 7604 29407
rect 7668 29209 7696 29532
rect 7654 29200 7710 29209
rect 7654 29135 7656 29144
rect 7708 29135 7710 29144
rect 7656 29106 7708 29112
rect 7668 28082 7696 29106
rect 7760 28778 7788 32506
rect 7852 31482 7880 33623
rect 7840 31476 7892 31482
rect 7840 31418 7892 31424
rect 7838 31240 7894 31249
rect 7838 31175 7840 31184
rect 7892 31175 7894 31184
rect 7840 31146 7892 31152
rect 7944 30190 7972 38218
rect 8128 37942 8156 39986
rect 8116 37936 8168 37942
rect 8116 37878 8168 37884
rect 8116 37392 8168 37398
rect 8220 37369 8248 42162
rect 8300 42084 8352 42090
rect 8300 42026 8352 42032
rect 8312 41993 8340 42026
rect 8298 41984 8354 41993
rect 8298 41919 8354 41928
rect 8496 41818 8524 42706
rect 8588 42362 8616 43318
rect 8772 42770 8800 44463
rect 9048 43450 9076 44463
rect 9036 43444 9088 43450
rect 9036 43386 9088 43392
rect 9128 43172 9180 43178
rect 9128 43114 9180 43120
rect 9140 42906 9168 43114
rect 9128 42900 9180 42906
rect 9128 42842 9180 42848
rect 9220 42832 9272 42838
rect 9220 42774 9272 42780
rect 8760 42764 8812 42770
rect 8760 42706 8812 42712
rect 9036 42696 9088 42702
rect 9036 42638 9088 42644
rect 9126 42664 9182 42673
rect 8576 42356 8628 42362
rect 8576 42298 8628 42304
rect 8484 41812 8536 41818
rect 8484 41754 8536 41760
rect 8852 41608 8904 41614
rect 8852 41550 8904 41556
rect 8576 41064 8628 41070
rect 8576 41006 8628 41012
rect 8392 40112 8444 40118
rect 8392 40054 8444 40060
rect 8404 39642 8432 40054
rect 8392 39636 8444 39642
rect 8392 39578 8444 39584
rect 8588 39438 8616 41006
rect 8668 39840 8720 39846
rect 8668 39782 8720 39788
rect 8680 39574 8708 39782
rect 8668 39568 8720 39574
rect 8668 39510 8720 39516
rect 8576 39432 8628 39438
rect 8576 39374 8628 39380
rect 8666 39400 8722 39409
rect 8300 39024 8352 39030
rect 8300 38966 8352 38972
rect 8312 38418 8340 38966
rect 8392 38956 8444 38962
rect 8392 38898 8444 38904
rect 8300 38412 8352 38418
rect 8300 38354 8352 38360
rect 8300 38004 8352 38010
rect 8300 37946 8352 37952
rect 8116 37334 8168 37340
rect 8206 37360 8262 37369
rect 8024 37256 8076 37262
rect 8024 37198 8076 37204
rect 8036 36922 8064 37198
rect 8024 36916 8076 36922
rect 8024 36858 8076 36864
rect 8024 36372 8076 36378
rect 8024 36314 8076 36320
rect 8036 34082 8064 36314
rect 8128 34406 8156 37334
rect 8206 37295 8262 37304
rect 8208 36916 8260 36922
rect 8208 36858 8260 36864
rect 8220 36718 8248 36858
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 8312 36564 8340 37946
rect 8404 36802 8432 38898
rect 8588 38758 8616 39374
rect 8666 39335 8722 39344
rect 8680 39030 8708 39335
rect 8668 39024 8720 39030
rect 8668 38966 8720 38972
rect 8576 38752 8628 38758
rect 8576 38694 8628 38700
rect 8484 37256 8536 37262
rect 8484 37198 8536 37204
rect 8496 36922 8524 37198
rect 8484 36916 8536 36922
rect 8484 36858 8536 36864
rect 8404 36774 8524 36802
rect 8220 36536 8340 36564
rect 8392 36576 8444 36582
rect 8220 35766 8248 36536
rect 8392 36518 8444 36524
rect 8208 35760 8260 35766
rect 8208 35702 8260 35708
rect 8220 34524 8248 35702
rect 8404 35630 8432 36518
rect 8392 35624 8444 35630
rect 8392 35566 8444 35572
rect 8496 35476 8524 36774
rect 8404 35448 8524 35476
rect 8404 35170 8432 35448
rect 8588 35170 8616 38694
rect 8668 38412 8720 38418
rect 8668 38354 8720 38360
rect 8680 37670 8708 38354
rect 8760 37936 8812 37942
rect 8760 37878 8812 37884
rect 8668 37664 8720 37670
rect 8668 37606 8720 37612
rect 8668 36168 8720 36174
rect 8668 36110 8720 36116
rect 8312 35142 8432 35170
rect 8496 35142 8616 35170
rect 8312 34649 8340 35142
rect 8496 34762 8524 35142
rect 8576 35080 8628 35086
rect 8576 35022 8628 35028
rect 8404 34734 8524 34762
rect 8298 34640 8354 34649
rect 8298 34575 8354 34584
rect 8220 34496 8340 34524
rect 8116 34400 8168 34406
rect 8116 34342 8168 34348
rect 8036 34054 8156 34082
rect 8024 33992 8076 33998
rect 8024 33934 8076 33940
rect 8036 33504 8064 33934
rect 8128 33697 8156 34054
rect 8114 33688 8170 33697
rect 8114 33623 8170 33632
rect 8208 33652 8260 33658
rect 8208 33594 8260 33600
rect 8116 33516 8168 33522
rect 8036 33476 8116 33504
rect 8116 33458 8168 33464
rect 8128 33114 8156 33458
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8024 32904 8076 32910
rect 8024 32846 8076 32852
rect 8036 31385 8064 32846
rect 8220 32473 8248 33594
rect 8206 32464 8262 32473
rect 8206 32399 8262 32408
rect 8312 32348 8340 34496
rect 8220 32320 8340 32348
rect 8116 31884 8168 31890
rect 8116 31826 8168 31832
rect 8022 31376 8078 31385
rect 8022 31311 8078 31320
rect 8036 30977 8064 31311
rect 8022 30968 8078 30977
rect 8022 30903 8078 30912
rect 8128 30258 8156 31826
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7852 29850 7880 29990
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 7840 29708 7892 29714
rect 7944 29696 7972 29990
rect 8116 29844 8168 29850
rect 7892 29668 7972 29696
rect 8036 29804 8116 29832
rect 7840 29650 7892 29656
rect 8036 29594 8064 29804
rect 8116 29786 8168 29792
rect 7944 29566 8064 29594
rect 8116 29640 8168 29646
rect 8116 29582 8168 29588
rect 7944 29510 7972 29566
rect 7932 29504 7984 29510
rect 7932 29446 7984 29452
rect 7760 28750 7880 28778
rect 7748 28552 7800 28558
rect 7748 28494 7800 28500
rect 7656 28076 7708 28082
rect 7656 28018 7708 28024
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26353 7696 27270
rect 7760 26926 7788 28494
rect 7852 27606 7880 28750
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7654 26344 7710 26353
rect 7654 26279 7710 26288
rect 7760 26246 7788 26862
rect 7484 26200 7604 26228
rect 7656 26240 7708 26246
rect 7484 23118 7512 26200
rect 7656 26182 7708 26188
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7668 26058 7696 26182
rect 7576 26030 7696 26058
rect 7576 25838 7604 26030
rect 7852 25974 7880 27406
rect 7656 25968 7708 25974
rect 7654 25936 7656 25945
rect 7840 25968 7892 25974
rect 7708 25936 7710 25945
rect 7840 25910 7892 25916
rect 7654 25871 7710 25880
rect 7748 25900 7800 25906
rect 7564 25832 7616 25838
rect 7564 25774 7616 25780
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7576 23118 7604 24006
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7564 23112 7616 23118
rect 7564 23054 7616 23060
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7300 21950 7420 21978
rect 6884 21788 7192 21797
rect 6884 21786 6890 21788
rect 6946 21786 6970 21788
rect 7026 21786 7050 21788
rect 7106 21786 7130 21788
rect 7186 21786 7192 21788
rect 6946 21734 6948 21786
rect 7128 21734 7130 21786
rect 6884 21732 6890 21734
rect 6946 21732 6970 21734
rect 7026 21732 7050 21734
rect 7106 21732 7130 21734
rect 7186 21732 7192 21734
rect 6884 21723 7192 21732
rect 7196 21548 7248 21554
rect 7196 21490 7248 21496
rect 6736 21480 6788 21486
rect 6736 21422 6788 21428
rect 7208 20913 7236 21490
rect 7194 20904 7250 20913
rect 7194 20839 7250 20848
rect 6884 20700 7192 20709
rect 6884 20698 6890 20700
rect 6946 20698 6970 20700
rect 7026 20698 7050 20700
rect 7106 20698 7130 20700
rect 7186 20698 7192 20700
rect 6946 20646 6948 20698
rect 7128 20646 7130 20698
rect 6884 20644 6890 20646
rect 6946 20644 6970 20646
rect 7026 20644 7050 20646
rect 7106 20644 7130 20646
rect 7186 20644 7192 20646
rect 6884 20635 7192 20644
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 19922 6592 20402
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6564 19334 6592 19858
rect 6656 19514 6684 20198
rect 6826 19816 6882 19825
rect 6826 19751 6882 19760
rect 6840 19718 6868 19751
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6564 19306 6684 19334
rect 6656 18834 6684 19306
rect 6644 18828 6696 18834
rect 6644 18770 6696 18776
rect 6748 18329 6776 19654
rect 6884 19612 7192 19621
rect 6884 19610 6890 19612
rect 6946 19610 6970 19612
rect 7026 19610 7050 19612
rect 7106 19610 7130 19612
rect 7186 19610 7192 19612
rect 6946 19558 6948 19610
rect 7128 19558 7130 19610
rect 6884 19556 6890 19558
rect 6946 19556 6970 19558
rect 7026 19556 7050 19558
rect 7106 19556 7130 19558
rect 7186 19556 7192 19558
rect 6884 19547 7192 19556
rect 7300 19334 7328 21950
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21622 7420 21830
rect 7484 21622 7512 22918
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 7472 21616 7524 21622
rect 7472 21558 7524 21564
rect 7576 19904 7604 22714
rect 7668 22166 7696 25871
rect 7748 25842 7800 25848
rect 7760 25498 7788 25842
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7944 24682 7972 29446
rect 8128 29306 8156 29582
rect 8116 29300 8168 29306
rect 8116 29242 8168 29248
rect 8116 28960 8168 28966
rect 8116 28902 8168 28908
rect 8128 28626 8156 28902
rect 8116 28620 8168 28626
rect 8116 28562 8168 28568
rect 8024 27600 8076 27606
rect 8024 27542 8076 27548
rect 8036 26790 8064 27542
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 8128 26994 8156 27066
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8024 26784 8076 26790
rect 8024 26726 8076 26732
rect 8036 25294 8064 26726
rect 8024 25288 8076 25294
rect 8128 25265 8156 26930
rect 8220 26908 8248 32320
rect 8404 32230 8432 34734
rect 8484 34672 8536 34678
rect 8484 34614 8536 34620
rect 8496 33862 8524 34614
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8392 32224 8444 32230
rect 8312 32184 8392 32212
rect 8312 30802 8340 32184
rect 8392 32166 8444 32172
rect 8392 31884 8444 31890
rect 8392 31826 8444 31832
rect 8404 30870 8432 31826
rect 8496 31822 8524 33798
rect 8484 31816 8536 31822
rect 8484 31758 8536 31764
rect 8392 30864 8444 30870
rect 8392 30806 8444 30812
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 8300 29708 8352 29714
rect 8300 29650 8352 29656
rect 8312 29492 8340 29650
rect 8392 29504 8444 29510
rect 8312 29464 8392 29492
rect 8312 29073 8340 29464
rect 8392 29446 8444 29452
rect 8298 29064 8354 29073
rect 8298 28999 8354 29008
rect 8496 27130 8524 31758
rect 8588 31754 8616 35022
rect 8680 33946 8708 36110
rect 8772 35698 8800 37878
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8772 35465 8800 35634
rect 8758 35456 8814 35465
rect 8758 35391 8814 35400
rect 8758 34096 8814 34105
rect 8758 34031 8760 34040
rect 8812 34031 8814 34040
rect 8760 34002 8812 34008
rect 8680 33918 8800 33946
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8680 33658 8708 33798
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8772 32910 8800 33918
rect 8760 32904 8812 32910
rect 8760 32846 8812 32852
rect 8760 32428 8812 32434
rect 8760 32370 8812 32376
rect 8588 31726 8708 31754
rect 8574 31512 8630 31521
rect 8574 31447 8630 31456
rect 8588 29306 8616 31447
rect 8576 29300 8628 29306
rect 8576 29242 8628 29248
rect 8588 29102 8616 29242
rect 8576 29096 8628 29102
rect 8576 29038 8628 29044
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 8220 26880 8616 26908
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8220 25974 8248 26318
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 8024 25230 8076 25236
rect 8114 25256 8170 25265
rect 7932 24676 7984 24682
rect 7932 24618 7984 24624
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7760 23798 7788 24006
rect 7748 23792 7800 23798
rect 7748 23734 7800 23740
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7944 23186 7972 23462
rect 7932 23180 7984 23186
rect 7932 23122 7984 23128
rect 7656 22160 7708 22166
rect 7656 22102 7708 22108
rect 8036 22094 8064 25230
rect 8114 25191 8170 25200
rect 8128 24970 8156 25191
rect 8206 24984 8262 24993
rect 8128 24942 8206 24970
rect 8206 24919 8262 24928
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8128 23526 8156 23666
rect 8116 23520 8168 23526
rect 8116 23462 8168 23468
rect 8114 23080 8170 23089
rect 8114 23015 8116 23024
rect 8168 23015 8170 23024
rect 8116 22986 8168 22992
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 7760 22066 8064 22094
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7668 21865 7696 21966
rect 7654 21856 7710 21865
rect 7654 21791 7710 21800
rect 7668 20806 7696 21791
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 7484 19876 7604 19904
rect 7656 19916 7708 19922
rect 7484 19514 7512 19876
rect 7656 19858 7708 19864
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7472 19372 7524 19378
rect 7300 19306 7420 19334
rect 7472 19314 7524 19320
rect 6884 18524 7192 18533
rect 6884 18522 6890 18524
rect 6946 18522 6970 18524
rect 7026 18522 7050 18524
rect 7106 18522 7130 18524
rect 7186 18522 7192 18524
rect 6946 18470 6948 18522
rect 7128 18470 7130 18522
rect 6884 18468 6890 18470
rect 6946 18468 6970 18470
rect 7026 18468 7050 18470
rect 7106 18468 7130 18470
rect 7186 18468 7192 18470
rect 6884 18459 7192 18468
rect 6734 18320 6790 18329
rect 6734 18255 6790 18264
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7300 17678 7328 18022
rect 6736 17672 6788 17678
rect 6736 17614 6788 17620
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 6460 17264 6512 17270
rect 6552 17264 6604 17270
rect 6460 17206 6512 17212
rect 6550 17232 6552 17241
rect 6604 17232 6606 17241
rect 6550 17167 6606 17176
rect 6288 17088 6500 17116
rect 6196 16510 6316 16538
rect 6182 16144 6238 16153
rect 6182 16079 6238 16088
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6104 14074 6132 14350
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6090 13424 6146 13433
rect 6090 13359 6146 13368
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6104 12714 6132 13359
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 5920 12566 6132 12594
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 5906 12336 5962 12345
rect 5828 12280 5906 12288
rect 5828 12260 5908 12280
rect 5960 12271 5962 12280
rect 5908 12242 5960 12248
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5828 10674 5856 10746
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5592 10152 5672 10180
rect 5540 10134 5592 10140
rect 5356 10124 5408 10130
rect 5356 10066 5408 10072
rect 5368 8090 5396 10066
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5552 7834 5580 10134
rect 5828 9926 5856 10610
rect 5920 10130 5948 12038
rect 6012 11898 6040 12378
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5998 10704 6054 10713
rect 5998 10639 6054 10648
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5276 7806 5580 7834
rect 5276 7410 5304 7806
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 5370 5304 7346
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5552 7002 5580 7278
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6458 5672 9862
rect 6012 9602 6040 10639
rect 5736 9574 6040 9602
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 6338 5764 9574
rect 5998 9480 6054 9489
rect 5998 9415 6054 9424
rect 6012 9382 6040 9415
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5828 6440 5856 7482
rect 5920 7002 5948 7754
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5828 6412 5948 6440
rect 5644 6310 5764 6338
rect 5816 6316 5868 6322
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 5914 5396 6054
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5276 5234 5304 5306
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5368 3738 5396 5578
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5552 4826 5580 5170
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5092 2746 5212 2774
rect 5092 2582 5120 2746
rect 5644 2650 5672 6310
rect 5816 6258 5868 6264
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 2774 5764 5510
rect 5828 5370 5856 6258
rect 5920 6254 5948 6412
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5914 5948 6054
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6012 5794 6040 8502
rect 6104 6322 6132 12566
rect 6196 10810 6224 16079
rect 6288 12889 6316 16510
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6380 15366 6408 15506
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6380 14074 6408 14894
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6274 12880 6330 12889
rect 6274 12815 6276 12824
rect 6328 12815 6330 12824
rect 6276 12786 6328 12792
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6196 6798 6224 10746
rect 6288 7954 6316 12582
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6288 6322 6316 7890
rect 6380 7886 6408 8842
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 5920 5766 6040 5794
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5920 5250 5948 5766
rect 5828 5222 5948 5250
rect 5828 3210 5856 5222
rect 5906 5128 5962 5137
rect 5906 5063 5962 5072
rect 5920 3398 5948 5063
rect 6000 5024 6052 5030
rect 5998 4992 6000 5001
rect 6052 4992 6054 5001
rect 5998 4927 6054 4936
rect 6196 4146 6224 6190
rect 6380 5914 6408 7142
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6380 5234 6408 5850
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6380 4690 6408 5170
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 5828 3182 5948 3210
rect 5736 2746 5856 2774
rect 5828 2650 5856 2746
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 4896 2440 4948 2446
rect 5724 2440 5776 2446
rect 4896 2382 4948 2388
rect 5644 2400 5724 2428
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 4342 54 4476 82
rect 4540 82 4568 1226
rect 4816 1000 4844 1906
rect 4908 1562 4936 2382
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5460 2106 5488 2246
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 5538 1864 5594 1873
rect 5538 1799 5594 1808
rect 5552 1766 5580 1799
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 4896 1556 4948 1562
rect 4896 1498 4948 1504
rect 5644 1442 5672 2400
rect 5724 2382 5776 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5828 2310 5856 2382
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5920 1970 5948 3182
rect 6012 2774 6040 3402
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6104 2990 6132 3334
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6012 2746 6132 2774
rect 6104 2310 6132 2746
rect 6182 2408 6238 2417
rect 6182 2343 6238 2352
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5460 1414 5672 1442
rect 5264 1352 5316 1358
rect 5264 1294 5316 1300
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 4816 972 4936 1000
rect 4908 160 4936 972
rect 5184 882 5212 1158
rect 5172 876 5224 882
rect 5172 818 5224 824
rect 4618 82 4674 160
rect 4540 54 4674 82
rect 4342 0 4398 54
rect 4618 0 4674 54
rect 4894 0 4950 160
rect 5170 82 5226 160
rect 5276 82 5304 1294
rect 5460 160 5488 1414
rect 5540 1352 5592 1358
rect 5538 1320 5540 1329
rect 5736 1340 5764 1906
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 5828 1494 5856 1838
rect 6104 1766 6132 2246
rect 6196 2038 6224 2343
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6184 2032 6236 2038
rect 6184 1974 6236 1980
rect 6092 1760 6144 1766
rect 6092 1702 6144 1708
rect 5816 1488 5868 1494
rect 5816 1430 5868 1436
rect 5592 1320 5594 1329
rect 5736 1312 6040 1340
rect 5538 1255 5594 1264
rect 5632 1284 5684 1290
rect 5684 1244 5764 1272
rect 5632 1226 5684 1232
rect 5736 160 5764 1244
rect 6012 160 6040 1312
rect 6288 1018 6316 2246
rect 6472 1902 6500 17088
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 15065 6592 15302
rect 6550 15056 6606 15065
rect 6550 14991 6606 15000
rect 6552 14544 6604 14550
rect 6552 14486 6604 14492
rect 6564 14006 6592 14486
rect 6656 14396 6684 15914
rect 6748 14634 6776 17614
rect 6884 17436 7192 17445
rect 6884 17434 6890 17436
rect 6946 17434 6970 17436
rect 7026 17434 7050 17436
rect 7106 17434 7130 17436
rect 7186 17434 7192 17436
rect 6946 17382 6948 17434
rect 7128 17382 7130 17434
rect 6884 17380 6890 17382
rect 6946 17380 6970 17382
rect 7026 17380 7050 17382
rect 7106 17380 7130 17382
rect 7186 17380 7192 17382
rect 6884 17371 7192 17380
rect 6918 17096 6974 17105
rect 6918 17031 6974 17040
rect 6932 16658 6960 17031
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 7288 16584 7340 16590
rect 7392 16561 7420 19306
rect 7484 18970 7512 19314
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7576 18873 7604 19722
rect 7668 19310 7696 19858
rect 7760 19825 7788 22066
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7838 21448 7894 21457
rect 7838 21383 7840 21392
rect 7892 21383 7894 21392
rect 7840 21354 7892 21360
rect 7838 21312 7894 21321
rect 7838 21247 7894 21256
rect 7852 20942 7880 21247
rect 7840 20936 7892 20942
rect 7838 20904 7840 20913
rect 7892 20904 7894 20913
rect 7838 20839 7894 20848
rect 7840 20596 7892 20602
rect 7840 20538 7892 20544
rect 7746 19816 7802 19825
rect 7746 19751 7802 19760
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7562 18864 7618 18873
rect 7562 18799 7618 18808
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17270 7512 17478
rect 7576 17338 7696 17354
rect 7576 17332 7708 17338
rect 7576 17326 7656 17332
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7470 16960 7526 16969
rect 7576 16946 7604 17326
rect 7656 17274 7708 17280
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7526 16918 7604 16946
rect 7470 16895 7526 16904
rect 7472 16652 7524 16658
rect 7472 16594 7524 16600
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7288 16526 7340 16532
rect 7378 16552 7434 16561
rect 6884 16348 7192 16357
rect 6884 16346 6890 16348
rect 6946 16346 6970 16348
rect 7026 16346 7050 16348
rect 7106 16346 7130 16348
rect 7186 16346 7192 16348
rect 6946 16294 6948 16346
rect 7128 16294 7130 16346
rect 6884 16292 6890 16294
rect 6946 16292 6970 16294
rect 7026 16292 7050 16294
rect 7106 16292 7130 16294
rect 7186 16292 7192 16294
rect 6884 16283 7192 16292
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6840 15570 6868 15914
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 7024 15502 7052 15982
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6884 15260 7192 15269
rect 6884 15258 6890 15260
rect 6946 15258 6970 15260
rect 7026 15258 7050 15260
rect 7106 15258 7130 15260
rect 7186 15258 7192 15260
rect 6946 15206 6948 15258
rect 7128 15206 7130 15258
rect 6884 15204 6890 15206
rect 6946 15204 6970 15206
rect 7026 15204 7050 15206
rect 7106 15204 7130 15206
rect 7186 15204 7192 15206
rect 6884 15195 7192 15204
rect 7300 15162 7328 16526
rect 7378 16487 7434 16496
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 6826 15056 6882 15065
rect 6826 14991 6882 15000
rect 6840 14940 6868 14991
rect 6920 14952 6972 14958
rect 6840 14912 6920 14940
rect 6920 14894 6972 14900
rect 6748 14606 7052 14634
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6736 14408 6788 14414
rect 6656 14368 6736 14396
rect 6840 14385 6868 14486
rect 7024 14414 7052 14606
rect 7012 14408 7064 14414
rect 6736 14350 6788 14356
rect 6826 14376 6882 14385
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6748 13938 6776 14350
rect 7012 14350 7064 14356
rect 6826 14311 6882 14320
rect 6884 14172 7192 14181
rect 6884 14170 6890 14172
rect 6946 14170 6970 14172
rect 7026 14170 7050 14172
rect 7106 14170 7130 14172
rect 7186 14170 7192 14172
rect 6946 14118 6948 14170
rect 7128 14118 7130 14170
rect 6884 14116 6890 14118
rect 6946 14116 6970 14118
rect 7026 14116 7050 14118
rect 7106 14116 7130 14118
rect 7186 14116 7192 14118
rect 6884 14107 7192 14116
rect 6736 13932 6788 13938
rect 6656 13892 6736 13920
rect 6656 13433 6684 13892
rect 6736 13874 6788 13880
rect 6642 13424 6698 13433
rect 6642 13359 6698 13368
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 6884 13084 7192 13093
rect 6884 13082 6890 13084
rect 6946 13082 6970 13084
rect 7026 13082 7050 13084
rect 7106 13082 7130 13084
rect 7186 13082 7192 13084
rect 6946 13030 6948 13082
rect 7128 13030 7130 13082
rect 6884 13028 6890 13030
rect 6946 13028 6970 13030
rect 7026 13028 7050 13030
rect 7106 13028 7130 13030
rect 7186 13028 7192 13030
rect 6884 13019 7192 13028
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 6840 12306 6868 12922
rect 7104 12708 7156 12714
rect 7104 12650 7156 12656
rect 6828 12300 6880 12306
rect 6656 12260 6828 12288
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 10674 6592 10746
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6656 10112 6684 12260
rect 6828 12242 6880 12248
rect 6920 12300 6972 12306
rect 7116 12288 7144 12650
rect 6972 12260 7144 12288
rect 6920 12242 6972 12248
rect 7208 12238 7236 12922
rect 7300 12850 7328 13330
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11354 6776 12038
rect 6884 11996 7192 12005
rect 6884 11994 6890 11996
rect 6946 11994 6970 11996
rect 7026 11994 7050 11996
rect 7106 11994 7130 11996
rect 7186 11994 7192 11996
rect 6946 11942 6948 11994
rect 7128 11942 7130 11994
rect 6884 11940 6890 11942
rect 6946 11940 6970 11942
rect 7026 11940 7050 11942
rect 7106 11940 7130 11942
rect 7186 11940 7192 11942
rect 6884 11931 7192 11940
rect 7300 11830 7328 12786
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11150 6868 11698
rect 7010 11248 7066 11257
rect 7010 11183 7066 11192
rect 7024 11150 7052 11183
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 6884 10908 7192 10917
rect 6884 10906 6890 10908
rect 6946 10906 6970 10908
rect 7026 10906 7050 10908
rect 7106 10906 7130 10908
rect 7186 10906 7192 10908
rect 6946 10854 6948 10906
rect 7128 10854 7130 10906
rect 6884 10852 6890 10854
rect 6946 10852 6970 10854
rect 7026 10852 7050 10854
rect 7106 10852 7130 10854
rect 7186 10852 7192 10854
rect 6884 10843 7192 10852
rect 6826 10568 6882 10577
rect 6826 10503 6882 10512
rect 6736 10124 6788 10130
rect 6656 10084 6736 10112
rect 6736 10066 6788 10072
rect 6840 10010 6868 10503
rect 6656 9982 6868 10010
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6564 7954 6592 9454
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6564 6322 6592 7890
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6564 5574 6592 5850
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6550 3632 6606 3641
rect 6550 3567 6606 3576
rect 6564 3126 6592 3567
rect 6656 3176 6684 9982
rect 6884 9820 7192 9829
rect 6884 9818 6890 9820
rect 6946 9818 6970 9820
rect 7026 9818 7050 9820
rect 7106 9818 7130 9820
rect 7186 9818 7192 9820
rect 6946 9766 6948 9818
rect 7128 9766 7130 9818
rect 6884 9764 6890 9766
rect 6946 9764 6970 9766
rect 7026 9764 7050 9766
rect 7106 9764 7130 9766
rect 7186 9764 7192 9766
rect 6884 9755 7192 9764
rect 7300 8906 7328 10950
rect 7392 10810 7420 15370
rect 7484 15026 7512 16594
rect 7576 15706 7604 16594
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7576 14618 7604 14894
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 14006 7512 14350
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7484 11354 7512 12310
rect 7576 11914 7604 14418
rect 7668 12084 7696 17138
rect 7760 15434 7788 19751
rect 7852 19378 7880 20538
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7852 16590 7880 17002
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7838 16144 7894 16153
rect 7838 16079 7840 16088
rect 7892 16079 7894 16088
rect 7840 16050 7892 16056
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7760 12152 7788 14894
rect 7840 13728 7892 13734
rect 7840 13670 7892 13676
rect 7852 12782 7880 13670
rect 7944 12986 7972 19450
rect 8036 19145 8064 21966
rect 8128 20890 8156 22442
rect 8220 21078 8248 24686
rect 8312 24206 8340 26182
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8404 24886 8432 25638
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8496 24750 8524 25230
rect 8484 24744 8536 24750
rect 8484 24686 8536 24692
rect 8392 24336 8444 24342
rect 8392 24278 8444 24284
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8312 22574 8340 24142
rect 8404 23662 8432 24278
rect 8392 23656 8444 23662
rect 8392 23598 8444 23604
rect 8392 23520 8444 23526
rect 8392 23462 8444 23468
rect 8404 23118 8432 23462
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8300 22568 8352 22574
rect 8300 22510 8352 22516
rect 8312 21185 8340 22510
rect 8496 22273 8524 24686
rect 8482 22264 8538 22273
rect 8482 22199 8538 22208
rect 8392 21616 8444 21622
rect 8392 21558 8444 21564
rect 8298 21176 8354 21185
rect 8404 21146 8432 21558
rect 8484 21480 8536 21486
rect 8484 21422 8536 21428
rect 8496 21146 8524 21422
rect 8298 21111 8354 21120
rect 8392 21140 8444 21146
rect 8208 21072 8260 21078
rect 8208 21014 8260 21020
rect 8128 20862 8248 20890
rect 8312 20874 8340 21111
rect 8392 21082 8444 21088
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8484 21004 8536 21010
rect 8484 20946 8536 20952
rect 8116 20800 8168 20806
rect 8114 20768 8116 20777
rect 8168 20768 8170 20777
rect 8114 20703 8170 20712
rect 8022 19136 8078 19145
rect 8022 19071 8078 19080
rect 8036 18766 8064 19071
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 8128 18442 8156 20703
rect 8220 20618 8248 20862
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8220 20590 8432 20618
rect 8404 19854 8432 20590
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8312 19514 8340 19790
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8208 19440 8260 19446
rect 8206 19408 8208 19417
rect 8260 19408 8262 19417
rect 8404 19378 8432 19790
rect 8206 19343 8262 19352
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8312 18698 8340 19314
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8128 18414 8248 18442
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 8128 13938 8156 18294
rect 8220 14482 8248 18414
rect 8300 18420 8352 18426
rect 8404 18408 8432 19314
rect 8352 18380 8432 18408
rect 8300 18362 8352 18368
rect 8312 18057 8340 18362
rect 8496 18290 8524 20946
rect 8588 19446 8616 26880
rect 8680 26586 8708 31726
rect 8772 30297 8800 32370
rect 8758 30288 8814 30297
rect 8758 30223 8814 30232
rect 8760 30116 8812 30122
rect 8760 30058 8812 30064
rect 8772 29510 8800 30058
rect 8864 29850 8892 41550
rect 8942 40216 8998 40225
rect 8942 40151 8998 40160
rect 8956 38010 8984 40151
rect 8944 38004 8996 38010
rect 8944 37946 8996 37952
rect 8944 37664 8996 37670
rect 8944 37606 8996 37612
rect 8956 36582 8984 37606
rect 9048 37262 9076 42638
rect 9126 42599 9182 42608
rect 9140 42566 9168 42599
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 9128 42356 9180 42362
rect 9128 42298 9180 42304
rect 9140 42226 9168 42298
rect 9128 42220 9180 42226
rect 9128 42162 9180 42168
rect 9128 40384 9180 40390
rect 9128 40326 9180 40332
rect 9140 40225 9168 40326
rect 9126 40216 9182 40225
rect 9126 40151 9182 40160
rect 9140 40118 9168 40151
rect 9232 40118 9260 42774
rect 9324 42770 9352 44463
rect 9600 43450 9628 44463
rect 9876 43450 9904 44463
rect 9588 43444 9640 43450
rect 9588 43386 9640 43392
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9404 43376 9456 43382
rect 9404 43318 9456 43324
rect 9416 43110 9444 43318
rect 9956 43308 10008 43314
rect 10152 43296 10180 44463
rect 10008 43268 10180 43296
rect 10324 43308 10376 43314
rect 9956 43250 10008 43256
rect 10428 43296 10456 44463
rect 10508 43648 10560 43654
rect 10508 43590 10560 43596
rect 10520 43450 10548 43590
rect 10508 43444 10560 43450
rect 10508 43386 10560 43392
rect 10704 43314 10732 44463
rect 10376 43268 10456 43296
rect 10692 43308 10744 43314
rect 10324 43250 10376 43256
rect 10980 43296 11008 44463
rect 11256 43314 11284 44463
rect 11532 43602 11560 44463
rect 11808 44146 11836 44463
rect 11808 44118 11928 44146
rect 11532 43574 11652 43602
rect 11060 43308 11112 43314
rect 10980 43268 11060 43296
rect 10692 43250 10744 43256
rect 11060 43250 11112 43256
rect 11244 43308 11296 43314
rect 11244 43250 11296 43256
rect 9680 43240 9732 43246
rect 9680 43182 9732 43188
rect 9404 43104 9456 43110
rect 9404 43046 9456 43052
rect 9692 42906 9720 43182
rect 10600 43104 10652 43110
rect 10600 43046 10652 43052
rect 10876 43104 10928 43110
rect 10876 43046 10928 43052
rect 11244 43104 11296 43110
rect 11244 43046 11296 43052
rect 9851 43004 10159 43013
rect 9851 43002 9857 43004
rect 9913 43002 9937 43004
rect 9993 43002 10017 43004
rect 10073 43002 10097 43004
rect 10153 43002 10159 43004
rect 9913 42950 9915 43002
rect 10095 42950 10097 43002
rect 9851 42948 9857 42950
rect 9913 42948 9937 42950
rect 9993 42948 10017 42950
rect 10073 42948 10097 42950
rect 10153 42948 10159 42950
rect 9851 42939 10159 42948
rect 10612 42906 10640 43046
rect 9680 42900 9732 42906
rect 9680 42842 9732 42848
rect 10600 42900 10652 42906
rect 10600 42842 10652 42848
rect 9402 42800 9458 42809
rect 9312 42764 9364 42770
rect 9402 42735 9458 42744
rect 9312 42706 9364 42712
rect 9416 42702 9444 42735
rect 9404 42696 9456 42702
rect 9404 42638 9456 42644
rect 9956 42696 10008 42702
rect 9956 42638 10008 42644
rect 9588 42628 9640 42634
rect 9588 42570 9640 42576
rect 9496 42356 9548 42362
rect 9496 42298 9548 42304
rect 9404 42220 9456 42226
rect 9404 42162 9456 42168
rect 9416 41857 9444 42162
rect 9508 42158 9536 42298
rect 9496 42152 9548 42158
rect 9496 42094 9548 42100
rect 9402 41848 9458 41857
rect 9402 41783 9458 41792
rect 9600 41414 9628 42570
rect 9968 42362 9996 42638
rect 10416 42628 10468 42634
rect 10416 42570 10468 42576
rect 9956 42356 10008 42362
rect 9956 42298 10008 42304
rect 9864 42220 9916 42226
rect 9864 42162 9916 42168
rect 9876 42129 9904 42162
rect 9862 42120 9918 42129
rect 9862 42055 9918 42064
rect 9851 41916 10159 41925
rect 9851 41914 9857 41916
rect 9913 41914 9937 41916
rect 9993 41914 10017 41916
rect 10073 41914 10097 41916
rect 10153 41914 10159 41916
rect 9913 41862 9915 41914
rect 10095 41862 10097 41914
rect 9851 41860 9857 41862
rect 9913 41860 9937 41862
rect 9993 41860 10017 41862
rect 10073 41860 10097 41862
rect 10153 41860 10159 41862
rect 9851 41851 10159 41860
rect 10048 41812 10100 41818
rect 10048 41754 10100 41760
rect 9508 41386 9628 41414
rect 9312 40588 9364 40594
rect 9312 40530 9364 40536
rect 9324 40186 9352 40530
rect 9508 40202 9536 41386
rect 10060 41070 10088 41754
rect 10324 41608 10376 41614
rect 10324 41550 10376 41556
rect 10048 41064 10100 41070
rect 10048 41006 10100 41012
rect 9588 40928 9640 40934
rect 9588 40870 9640 40876
rect 9680 40928 9732 40934
rect 9680 40870 9732 40876
rect 9312 40180 9364 40186
rect 9312 40122 9364 40128
rect 9416 40174 9536 40202
rect 9128 40112 9180 40118
rect 9128 40054 9180 40060
rect 9220 40112 9272 40118
rect 9220 40054 9272 40060
rect 9128 38752 9180 38758
rect 9128 38694 9180 38700
rect 9140 37806 9168 38694
rect 9232 38554 9260 40054
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 9232 37942 9260 38490
rect 9220 37936 9272 37942
rect 9220 37878 9272 37884
rect 9128 37800 9180 37806
rect 9128 37742 9180 37748
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 8944 36576 8996 36582
rect 8944 36518 8996 36524
rect 8956 36242 8984 36518
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8942 36136 8998 36145
rect 8942 36071 8998 36080
rect 8956 34898 8984 36071
rect 8956 34870 9076 34898
rect 9048 34746 9076 34870
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 9036 34740 9088 34746
rect 9036 34682 9088 34688
rect 8956 34626 8984 34682
rect 9034 34640 9090 34649
rect 8956 34598 9034 34626
rect 9140 34626 9168 36722
rect 9232 35766 9260 37878
rect 9312 36780 9364 36786
rect 9312 36722 9364 36728
rect 9324 36174 9352 36722
rect 9312 36168 9364 36174
rect 9416 36145 9444 40174
rect 9496 40112 9548 40118
rect 9496 40054 9548 40060
rect 9508 39642 9536 40054
rect 9600 39982 9628 40870
rect 9692 40730 9720 40870
rect 9851 40828 10159 40837
rect 9851 40826 9857 40828
rect 9913 40826 9937 40828
rect 9993 40826 10017 40828
rect 10073 40826 10097 40828
rect 10153 40826 10159 40828
rect 9913 40774 9915 40826
rect 10095 40774 10097 40826
rect 9851 40772 9857 40774
rect 9913 40772 9937 40774
rect 9993 40772 10017 40774
rect 10073 40772 10097 40774
rect 10153 40772 10159 40774
rect 9851 40763 10159 40772
rect 9680 40724 9732 40730
rect 9680 40666 9732 40672
rect 9772 40724 9824 40730
rect 9772 40666 9824 40672
rect 9784 40526 9812 40666
rect 10336 40662 10364 41550
rect 10324 40656 10376 40662
rect 10324 40598 10376 40604
rect 10048 40588 10100 40594
rect 10048 40530 10100 40536
rect 9772 40520 9824 40526
rect 9772 40462 9824 40468
rect 9956 40520 10008 40526
rect 9956 40462 10008 40468
rect 9772 40384 9824 40390
rect 9968 40372 9996 40462
rect 9824 40344 9996 40372
rect 9772 40326 9824 40332
rect 10060 40118 10088 40530
rect 10336 40118 10364 40598
rect 9772 40112 9824 40118
rect 9772 40054 9824 40060
rect 10048 40112 10100 40118
rect 10048 40054 10100 40060
rect 10324 40112 10376 40118
rect 10324 40054 10376 40060
rect 9680 40044 9732 40050
rect 9680 39986 9732 39992
rect 9588 39976 9640 39982
rect 9588 39918 9640 39924
rect 9496 39636 9548 39642
rect 9496 39578 9548 39584
rect 9496 38344 9548 38350
rect 9496 38286 9548 38292
rect 9508 37942 9536 38286
rect 9496 37936 9548 37942
rect 9496 37878 9548 37884
rect 9692 37874 9720 39986
rect 9784 37874 9812 40054
rect 10324 39840 10376 39846
rect 10324 39782 10376 39788
rect 9851 39740 10159 39749
rect 9851 39738 9857 39740
rect 9913 39738 9937 39740
rect 9993 39738 10017 39740
rect 10073 39738 10097 39740
rect 10153 39738 10159 39740
rect 9913 39686 9915 39738
rect 10095 39686 10097 39738
rect 9851 39684 9857 39686
rect 9913 39684 9937 39686
rect 9993 39684 10017 39686
rect 10073 39684 10097 39686
rect 10153 39684 10159 39686
rect 9851 39675 10159 39684
rect 10232 39432 10284 39438
rect 10232 39374 10284 39380
rect 10244 39250 10272 39374
rect 10336 39370 10364 39782
rect 10324 39364 10376 39370
rect 10324 39306 10376 39312
rect 10244 39222 10364 39250
rect 9851 38652 10159 38661
rect 9851 38650 9857 38652
rect 9913 38650 9937 38652
rect 9993 38650 10017 38652
rect 10073 38650 10097 38652
rect 10153 38650 10159 38652
rect 9913 38598 9915 38650
rect 10095 38598 10097 38650
rect 9851 38596 9857 38598
rect 9913 38596 9937 38598
rect 9993 38596 10017 38598
rect 10073 38596 10097 38598
rect 10153 38596 10159 38598
rect 9851 38587 10159 38596
rect 10140 38208 10192 38214
rect 10140 38150 10192 38156
rect 10152 38010 10180 38150
rect 10140 38004 10192 38010
rect 10140 37946 10192 37952
rect 9680 37868 9732 37874
rect 9680 37810 9732 37816
rect 9772 37868 9824 37874
rect 9772 37810 9824 37816
rect 9784 37754 9812 37810
rect 9692 37726 9812 37754
rect 9692 37210 9720 37726
rect 9851 37564 10159 37573
rect 9851 37562 9857 37564
rect 9913 37562 9937 37564
rect 9993 37562 10017 37564
rect 10073 37562 10097 37564
rect 10153 37562 10159 37564
rect 9913 37510 9915 37562
rect 10095 37510 10097 37562
rect 9851 37508 9857 37510
rect 9913 37508 9937 37510
rect 9993 37508 10017 37510
rect 10073 37508 10097 37510
rect 10153 37508 10159 37510
rect 9851 37499 10159 37508
rect 9600 37182 9720 37210
rect 10048 37256 10100 37262
rect 10048 37198 10100 37204
rect 9772 37188 9824 37194
rect 9312 36110 9364 36116
rect 9402 36136 9458 36145
rect 9402 36071 9458 36080
rect 9220 35760 9272 35766
rect 9220 35702 9272 35708
rect 9600 35698 9628 37182
rect 9772 37130 9824 37136
rect 9784 36854 9812 37130
rect 9772 36848 9824 36854
rect 9772 36790 9824 36796
rect 10060 36718 10088 37198
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 9851 36476 10159 36485
rect 9851 36474 9857 36476
rect 9913 36474 9937 36476
rect 9993 36474 10017 36476
rect 10073 36474 10097 36476
rect 10153 36474 10159 36476
rect 9913 36422 9915 36474
rect 10095 36422 10097 36474
rect 9851 36420 9857 36422
rect 9913 36420 9937 36422
rect 9993 36420 10017 36422
rect 10073 36420 10097 36422
rect 10153 36420 10159 36422
rect 9851 36411 10159 36420
rect 9864 36236 9916 36242
rect 9864 36178 9916 36184
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9588 35692 9640 35698
rect 9588 35634 9640 35640
rect 9312 35624 9364 35630
rect 9232 35584 9312 35612
rect 9232 34921 9260 35584
rect 9312 35566 9364 35572
rect 9600 35290 9628 35634
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 9600 34921 9628 35226
rect 9692 35086 9720 36110
rect 9876 36038 9904 36178
rect 10140 36100 10192 36106
rect 10140 36042 10192 36048
rect 9864 36032 9916 36038
rect 9864 35974 9916 35980
rect 9956 36032 10008 36038
rect 9956 35974 10008 35980
rect 9968 35834 9996 35974
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 9772 35488 9824 35494
rect 10152 35476 10180 36042
rect 10152 35448 10272 35476
rect 9772 35430 9824 35436
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9218 34912 9274 34921
rect 9218 34847 9274 34856
rect 9586 34912 9642 34921
rect 9586 34847 9642 34856
rect 9232 34746 9260 34847
rect 9220 34740 9272 34746
rect 9220 34682 9272 34688
rect 9680 34672 9732 34678
rect 9140 34598 9352 34626
rect 9680 34614 9732 34620
rect 9034 34575 9090 34584
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 9036 34400 9088 34406
rect 9088 34377 9168 34388
rect 9088 34368 9182 34377
rect 9088 34360 9126 34368
rect 9036 34342 9088 34348
rect 9126 34303 9182 34312
rect 8944 33992 8996 33998
rect 8942 33960 8944 33969
rect 8996 33960 8998 33969
rect 8942 33895 8998 33904
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8956 31414 8984 33798
rect 9232 33590 9260 34478
rect 9220 33584 9272 33590
rect 9220 33526 9272 33532
rect 9036 32972 9088 32978
rect 9036 32914 9088 32920
rect 9048 32314 9076 32914
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9048 32286 9168 32314
rect 9036 32224 9088 32230
rect 9036 32166 9088 32172
rect 9048 31686 9076 32166
rect 9140 31890 9168 32286
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 9232 31754 9260 32846
rect 9324 32366 9352 34598
rect 9588 34604 9640 34610
rect 9588 34546 9640 34552
rect 9496 34400 9548 34406
rect 9494 34368 9496 34377
rect 9548 34368 9550 34377
rect 9494 34303 9550 34312
rect 9496 33652 9548 33658
rect 9600 33640 9628 34546
rect 9692 34202 9720 34614
rect 9784 34542 9812 35430
rect 9851 35388 10159 35397
rect 9851 35386 9857 35388
rect 9913 35386 9937 35388
rect 9993 35386 10017 35388
rect 10073 35386 10097 35388
rect 10153 35386 10159 35388
rect 9913 35334 9915 35386
rect 10095 35334 10097 35386
rect 9851 35332 9857 35334
rect 9913 35332 9937 35334
rect 9993 35332 10017 35334
rect 10073 35332 10097 35334
rect 10153 35332 10159 35334
rect 9851 35323 10159 35332
rect 10244 35272 10272 35448
rect 10152 35244 10272 35272
rect 10046 35184 10102 35193
rect 10152 35154 10180 35244
rect 10046 35119 10102 35128
rect 10140 35148 10192 35154
rect 10060 35034 10088 35119
rect 10336 35136 10364 39222
rect 10428 35873 10456 42570
rect 10692 41472 10744 41478
rect 10692 41414 10744 41420
rect 10520 41386 10732 41414
rect 10520 40662 10548 41386
rect 10508 40656 10560 40662
rect 10508 40598 10560 40604
rect 10888 40594 10916 43046
rect 11060 40928 11112 40934
rect 11060 40870 11112 40876
rect 11072 40594 11100 40870
rect 10876 40588 10928 40594
rect 10876 40530 10928 40536
rect 11060 40588 11112 40594
rect 11060 40530 11112 40536
rect 10784 40520 10836 40526
rect 10784 40462 10836 40468
rect 10796 40118 10824 40462
rect 10692 40112 10744 40118
rect 10692 40054 10744 40060
rect 10784 40112 10836 40118
rect 10784 40054 10836 40060
rect 10600 37664 10652 37670
rect 10600 37606 10652 37612
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 10414 35864 10470 35873
rect 10414 35799 10470 35808
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10428 35329 10456 35634
rect 10414 35320 10470 35329
rect 10414 35255 10470 35264
rect 10416 35216 10468 35222
rect 10416 35158 10468 35164
rect 10140 35090 10192 35096
rect 10244 35108 10364 35136
rect 10244 35034 10272 35108
rect 10428 35068 10456 35158
rect 9956 35012 10008 35018
rect 9956 34954 10008 34960
rect 10060 35006 10272 35034
rect 10336 35040 10456 35068
rect 9968 34746 9996 34954
rect 9864 34740 9916 34746
rect 9864 34682 9916 34688
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9876 34406 9904 34682
rect 10060 34678 10088 35006
rect 10048 34672 10100 34678
rect 10048 34614 10100 34620
rect 10048 34536 10100 34542
rect 10048 34478 10100 34484
rect 9864 34400 9916 34406
rect 10060 34388 10088 34478
rect 10060 34360 10272 34388
rect 9864 34342 9916 34348
rect 9851 34300 10159 34309
rect 9851 34298 9857 34300
rect 9913 34298 9937 34300
rect 9993 34298 10017 34300
rect 10073 34298 10097 34300
rect 10153 34298 10159 34300
rect 9913 34246 9915 34298
rect 10095 34246 10097 34298
rect 9851 34244 9857 34246
rect 9913 34244 9937 34246
rect 9993 34244 10017 34246
rect 10073 34244 10097 34246
rect 10153 34244 10159 34246
rect 9851 34235 10159 34244
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9680 34060 9732 34066
rect 9680 34002 9732 34008
rect 9692 33658 9720 34002
rect 10244 33998 10272 34360
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 9548 33612 9628 33640
rect 9680 33652 9732 33658
rect 9496 33594 9548 33600
rect 9680 33594 9732 33600
rect 9416 33510 9720 33538
rect 9416 33289 9444 33510
rect 9402 33280 9458 33289
rect 9402 33215 9458 33224
rect 9312 32360 9364 32366
rect 9312 32302 9364 32308
rect 9140 31726 9260 31754
rect 9036 31680 9088 31686
rect 9036 31622 9088 31628
rect 8944 31408 8996 31414
rect 8944 31350 8996 31356
rect 9036 31408 9088 31414
rect 9036 31350 9088 31356
rect 9048 30938 9076 31350
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 8944 30796 8996 30802
rect 8944 30738 8996 30744
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 8760 29504 8812 29510
rect 8760 29446 8812 29452
rect 8772 29170 8800 29446
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 8760 27532 8812 27538
rect 8760 27474 8812 27480
rect 8772 27130 8800 27474
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8668 26580 8720 26586
rect 8668 26522 8720 26528
rect 8666 26208 8722 26217
rect 8666 26143 8722 26152
rect 8680 24818 8708 26143
rect 8760 25832 8812 25838
rect 8758 25800 8760 25809
rect 8812 25800 8814 25809
rect 8758 25735 8814 25744
rect 8758 25528 8814 25537
rect 8758 25463 8814 25472
rect 8772 25226 8800 25463
rect 8760 25220 8812 25226
rect 8760 25162 8812 25168
rect 8864 24818 8892 29242
rect 8956 29073 8984 30738
rect 9140 30734 9168 31726
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9232 31278 9260 31622
rect 9220 31272 9272 31278
rect 9220 31214 9272 31220
rect 9128 30728 9180 30734
rect 9128 30670 9180 30676
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 8942 29064 8998 29073
rect 8942 28999 8998 29008
rect 9048 28506 9076 29786
rect 8956 28478 9076 28506
rect 8956 25945 8984 28478
rect 9036 28416 9088 28422
rect 9036 28358 9088 28364
rect 8942 25936 8998 25945
rect 8942 25871 8998 25880
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8852 24812 8904 24818
rect 8852 24754 8904 24760
rect 8680 21010 8708 24754
rect 8864 23798 8892 24754
rect 9048 24410 9076 28358
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 9140 22234 9168 30670
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9232 28422 9260 28494
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9232 26926 9260 27270
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9324 26874 9352 32302
rect 9508 31498 9536 33510
rect 9692 33114 9720 33510
rect 9864 33516 9916 33522
rect 9864 33458 9916 33464
rect 9876 33425 9904 33458
rect 9862 33416 9918 33425
rect 9862 33351 9918 33360
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9680 33108 9732 33114
rect 9680 33050 9732 33056
rect 9784 32434 9812 33254
rect 9851 33212 10159 33221
rect 9851 33210 9857 33212
rect 9913 33210 9937 33212
rect 9993 33210 10017 33212
rect 10073 33210 10097 33212
rect 10153 33210 10159 33212
rect 9913 33158 9915 33210
rect 10095 33158 10097 33210
rect 9851 33156 9857 33158
rect 9913 33156 9937 33158
rect 9993 33156 10017 33158
rect 10073 33156 10097 33158
rect 10153 33156 10159 33158
rect 9851 33147 10159 33156
rect 10140 32496 10192 32502
rect 10140 32438 10192 32444
rect 9772 32428 9824 32434
rect 9772 32370 9824 32376
rect 10152 32337 10180 32438
rect 10138 32328 10194 32337
rect 10138 32263 10194 32272
rect 9851 32124 10159 32133
rect 9851 32122 9857 32124
rect 9913 32122 9937 32124
rect 9993 32122 10017 32124
rect 10073 32122 10097 32124
rect 10153 32122 10159 32124
rect 9913 32070 9915 32122
rect 10095 32070 10097 32122
rect 9851 32068 9857 32070
rect 9913 32068 9937 32070
rect 9993 32068 10017 32070
rect 10073 32068 10097 32070
rect 10153 32068 10159 32070
rect 9851 32059 10159 32068
rect 9588 32020 9640 32026
rect 9588 31962 9640 31968
rect 9600 31668 9628 31962
rect 9600 31640 9674 31668
rect 9646 31634 9674 31640
rect 9646 31606 9904 31634
rect 9508 31470 9628 31498
rect 9404 31340 9456 31346
rect 9456 31300 9536 31328
rect 9404 31282 9456 31288
rect 9404 30320 9456 30326
rect 9404 30262 9456 30268
rect 9416 29714 9444 30262
rect 9404 29708 9456 29714
rect 9404 29650 9456 29656
rect 9508 29220 9536 31300
rect 9600 29424 9628 31470
rect 9772 31408 9824 31414
rect 9692 31356 9772 31362
rect 9692 31350 9824 31356
rect 9692 31334 9812 31350
rect 9692 31113 9720 31334
rect 9876 31260 9904 31606
rect 9784 31232 9904 31260
rect 9678 31104 9734 31113
rect 9678 31039 9734 31048
rect 9784 29832 9812 31232
rect 9851 31036 10159 31045
rect 9851 31034 9857 31036
rect 9913 31034 9937 31036
rect 9993 31034 10017 31036
rect 10073 31034 10097 31036
rect 10153 31034 10159 31036
rect 9913 30982 9915 31034
rect 10095 30982 10097 31034
rect 9851 30980 9857 30982
rect 9913 30980 9937 30982
rect 9993 30980 10017 30982
rect 10073 30980 10097 30982
rect 10153 30980 10159 30982
rect 9851 30971 10159 30980
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10152 30705 10180 30874
rect 10138 30696 10194 30705
rect 10336 30666 10364 35040
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10428 34610 10456 34682
rect 10416 34604 10468 34610
rect 10416 34546 10468 34552
rect 10520 33980 10548 36518
rect 10612 36242 10640 37606
rect 10600 36236 10652 36242
rect 10600 36178 10652 36184
rect 10600 35488 10652 35494
rect 10600 35430 10652 35436
rect 10612 35222 10640 35430
rect 10600 35216 10652 35222
rect 10600 35158 10652 35164
rect 10704 35068 10732 40054
rect 11256 37126 11284 43046
rect 11624 42702 11652 43574
rect 11704 43104 11756 43110
rect 11704 43046 11756 43052
rect 11716 42945 11744 43046
rect 11702 42936 11758 42945
rect 11702 42871 11758 42880
rect 11900 42702 11928 44118
rect 12084 43314 12112 44463
rect 12360 43364 12388 44463
rect 12440 43376 12492 43382
rect 12360 43336 12440 43364
rect 12636 43364 12664 44463
rect 12912 43738 12940 44463
rect 13188 43874 13216 44463
rect 13188 43846 13400 43874
rect 12912 43710 13216 43738
rect 12818 43548 13126 43557
rect 12818 43546 12824 43548
rect 12880 43546 12904 43548
rect 12960 43546 12984 43548
rect 13040 43546 13064 43548
rect 13120 43546 13126 43548
rect 12880 43494 12882 43546
rect 13062 43494 13064 43546
rect 12818 43492 12824 43494
rect 12880 43492 12904 43494
rect 12960 43492 12984 43494
rect 13040 43492 13064 43494
rect 13120 43492 13126 43494
rect 12818 43483 13126 43492
rect 12808 43376 12860 43382
rect 12636 43336 12808 43364
rect 12440 43318 12492 43324
rect 13188 43364 13216 43710
rect 13372 43450 13400 43846
rect 13360 43444 13412 43450
rect 13360 43386 13412 43392
rect 13464 43382 13492 44463
rect 12808 43318 12860 43324
rect 13004 43336 13216 43364
rect 13452 43376 13504 43382
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 12256 43104 12308 43110
rect 12256 43046 12308 43052
rect 12532 43104 12584 43110
rect 12532 43046 12584 43052
rect 12624 43104 12676 43110
rect 12624 43046 12676 43052
rect 12268 42945 12296 43046
rect 12544 42945 12572 43046
rect 12254 42936 12310 42945
rect 12254 42871 12310 42880
rect 12530 42936 12586 42945
rect 12530 42871 12586 42880
rect 12256 42764 12308 42770
rect 12256 42706 12308 42712
rect 12440 42764 12492 42770
rect 12440 42706 12492 42712
rect 11612 42696 11664 42702
rect 11612 42638 11664 42644
rect 11888 42696 11940 42702
rect 11888 42638 11940 42644
rect 11336 42628 11388 42634
rect 11336 42570 11388 42576
rect 11348 38486 11376 42570
rect 11796 42560 11848 42566
rect 11796 42502 11848 42508
rect 12164 42560 12216 42566
rect 12164 42502 12216 42508
rect 11808 42265 11836 42502
rect 11794 42256 11850 42265
rect 12176 42226 12204 42502
rect 11794 42191 11850 42200
rect 12164 42220 12216 42226
rect 12164 42162 12216 42168
rect 11796 40724 11848 40730
rect 11796 40666 11848 40672
rect 11704 40520 11756 40526
rect 11704 40462 11756 40468
rect 11520 40384 11572 40390
rect 11440 40344 11520 40372
rect 11440 39982 11468 40344
rect 11520 40326 11572 40332
rect 11428 39976 11480 39982
rect 11428 39918 11480 39924
rect 11336 38480 11388 38486
rect 11336 38422 11388 38428
rect 11336 38344 11388 38350
rect 11336 38286 11388 38292
rect 11060 37120 11112 37126
rect 11060 37062 11112 37068
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 10784 36712 10836 36718
rect 10784 36654 10836 36660
rect 10612 35040 10732 35068
rect 10612 34524 10640 35040
rect 10692 34672 10744 34678
rect 10690 34640 10692 34649
rect 10744 34640 10746 34649
rect 10690 34575 10746 34584
rect 10612 34496 10732 34524
rect 10520 33952 10640 33980
rect 10508 33312 10560 33318
rect 10508 33254 10560 33260
rect 10520 33046 10548 33254
rect 10508 33040 10560 33046
rect 10508 32982 10560 32988
rect 10612 32858 10640 33952
rect 10704 33658 10732 34496
rect 10692 33652 10744 33658
rect 10692 33594 10744 33600
rect 10692 33516 10744 33522
rect 10692 33458 10744 33464
rect 10704 32978 10732 33458
rect 10796 33318 10824 36654
rect 11072 36310 11100 37062
rect 11060 36304 11112 36310
rect 11060 36246 11112 36252
rect 11244 36168 11296 36174
rect 11244 36110 11296 36116
rect 11256 35766 11284 36110
rect 11244 35760 11296 35766
rect 11244 35702 11296 35708
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 10980 35086 11008 35634
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 11060 35080 11112 35086
rect 11060 35022 11112 35028
rect 10876 34400 10928 34406
rect 10876 34342 10928 34348
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10692 32972 10744 32978
rect 10692 32914 10744 32920
rect 10888 32910 10916 34342
rect 10980 34134 11008 35022
rect 11072 34746 11100 35022
rect 11060 34740 11112 34746
rect 11060 34682 11112 34688
rect 10968 34128 11020 34134
rect 10968 34070 11020 34076
rect 11256 33969 11284 35090
rect 11242 33960 11298 33969
rect 11242 33895 11298 33904
rect 11060 33584 11112 33590
rect 11060 33526 11112 33532
rect 10876 32904 10928 32910
rect 10612 32830 10732 32858
rect 10928 32864 11008 32892
rect 10876 32846 10928 32852
rect 10416 32768 10468 32774
rect 10416 32710 10468 32716
rect 10428 30802 10456 32710
rect 10600 32496 10652 32502
rect 10600 32438 10652 32444
rect 10612 31346 10640 32438
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10416 30796 10468 30802
rect 10416 30738 10468 30744
rect 10138 30631 10194 30640
rect 10324 30660 10376 30666
rect 10152 30258 10180 30631
rect 10324 30602 10376 30608
rect 10428 30546 10456 30738
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10704 30682 10732 32830
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10888 32042 10916 32370
rect 10796 32014 10916 32042
rect 10796 30802 10824 32014
rect 10874 31920 10930 31929
rect 10874 31855 10930 31864
rect 10888 31822 10916 31855
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 10876 31204 10928 31210
rect 10876 31146 10928 31152
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10508 30660 10560 30666
rect 10508 30602 10560 30608
rect 10336 30518 10456 30546
rect 10336 30376 10364 30518
rect 10336 30348 10456 30376
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 9851 29948 10159 29957
rect 9851 29946 9857 29948
rect 9913 29946 9937 29948
rect 9993 29946 10017 29948
rect 10073 29946 10097 29948
rect 10153 29946 10159 29948
rect 9913 29894 9915 29946
rect 10095 29894 10097 29946
rect 9851 29892 9857 29894
rect 9913 29892 9937 29894
rect 9993 29892 10017 29894
rect 10073 29892 10097 29894
rect 10153 29892 10159 29894
rect 9851 29883 10159 29892
rect 9784 29804 9904 29832
rect 9772 29572 9824 29578
rect 9772 29514 9824 29520
rect 9600 29396 9720 29424
rect 9506 29192 9536 29220
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9416 28801 9444 29106
rect 9506 29084 9534 29192
rect 9506 29056 9536 29084
rect 9402 28792 9458 28801
rect 9402 28727 9458 28736
rect 9416 28529 9444 28727
rect 9402 28520 9458 28529
rect 9402 28455 9458 28464
rect 9404 27396 9456 27402
rect 9404 27338 9456 27344
rect 9416 27130 9444 27338
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9324 26846 9444 26874
rect 9312 26784 9364 26790
rect 9312 26726 9364 26732
rect 9324 26382 9352 26726
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 9220 23792 9272 23798
rect 9220 23734 9272 23740
rect 9232 22778 9260 23734
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9036 22228 9088 22234
rect 9036 22170 9088 22176
rect 9128 22228 9180 22234
rect 9128 22170 9180 22176
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8956 21554 8984 21626
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8944 21548 8996 21554
rect 8944 21490 8996 21496
rect 8668 21004 8720 21010
rect 8668 20946 8720 20952
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8680 20398 8708 20742
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8680 19334 8708 20334
rect 8588 19306 8708 19334
rect 8484 18284 8536 18290
rect 8404 18244 8484 18272
rect 8298 18048 8354 18057
rect 8298 17983 8354 17992
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 8036 12850 8064 13262
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7838 12336 7894 12345
rect 7838 12271 7840 12280
rect 7892 12271 7894 12280
rect 7840 12242 7892 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7760 12124 7880 12152
rect 7668 12056 7788 12084
rect 7576 11886 7696 11914
rect 7562 11792 7618 11801
rect 7562 11727 7618 11736
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7576 10985 7604 11727
rect 7562 10976 7618 10985
rect 7562 10911 7618 10920
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7392 10266 7420 10406
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 6884 8732 7192 8741
rect 6884 8730 6890 8732
rect 6946 8730 6970 8732
rect 7026 8730 7050 8732
rect 7106 8730 7130 8732
rect 7186 8730 7192 8732
rect 6946 8678 6948 8730
rect 7128 8678 7130 8730
rect 6884 8676 6890 8678
rect 6946 8676 6970 8678
rect 7026 8676 7050 8678
rect 7106 8676 7130 8678
rect 7186 8676 7192 8678
rect 6884 8667 7192 8676
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 7546 6776 8366
rect 7194 8120 7250 8129
rect 7300 8090 7328 8434
rect 7392 8430 7420 8842
rect 7484 8480 7512 10406
rect 7576 10266 7604 10474
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9178 7604 9522
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7668 8906 7696 11886
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7564 8492 7616 8498
rect 7484 8452 7564 8480
rect 7564 8434 7616 8440
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7194 8055 7196 8064
rect 7248 8055 7250 8064
rect 7288 8084 7340 8090
rect 7196 8026 7248 8032
rect 7288 8026 7340 8032
rect 7208 7732 7236 8026
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7208 7704 7328 7732
rect 6884 7644 7192 7653
rect 6884 7642 6890 7644
rect 6946 7642 6970 7644
rect 7026 7642 7050 7644
rect 7106 7642 7130 7644
rect 7186 7642 7192 7644
rect 6946 7590 6948 7642
rect 7128 7590 7130 7642
rect 6884 7588 6890 7590
rect 6946 7588 6970 7590
rect 7026 7588 7050 7590
rect 7106 7588 7130 7590
rect 7186 7588 7192 7590
rect 6884 7579 7192 7588
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6748 5234 6776 6802
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 7300 6322 7328 7704
rect 7392 6322 7420 7890
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 7546 7512 7822
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7576 6866 7604 8434
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 7012 6180 7064 6186
rect 7012 6122 7064 6128
rect 6840 5778 6868 6122
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6932 5681 6960 6054
rect 6918 5672 6974 5681
rect 7024 5642 7052 6122
rect 7300 5794 7328 6258
rect 7472 5908 7524 5914
rect 7576 5896 7604 6258
rect 7524 5868 7604 5896
rect 7472 5850 7524 5856
rect 7470 5808 7526 5817
rect 7300 5766 7470 5794
rect 7470 5743 7526 5752
rect 7286 5672 7342 5681
rect 6918 5607 6974 5616
rect 7012 5636 7064 5642
rect 7286 5607 7342 5616
rect 7380 5636 7432 5642
rect 7012 5578 7064 5584
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6826 4584 6882 4593
rect 6826 4519 6828 4528
rect 6880 4519 6882 4528
rect 6828 4490 6880 4496
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6748 3602 6776 4082
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 7300 3534 7328 5607
rect 7380 5578 7432 5584
rect 7392 5370 7420 5578
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 7300 3194 7328 3334
rect 7484 3194 7512 5743
rect 7668 5574 7696 8842
rect 7760 8566 7788 12056
rect 7852 11898 7880 12124
rect 8036 11898 8064 12174
rect 7840 11892 7892 11898
rect 7840 11834 7892 11840
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7852 6984 7880 11086
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 7930 10024 7986 10033
rect 7930 9959 7986 9968
rect 7760 6956 7880 6984
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7760 4282 7788 6956
rect 7838 6896 7894 6905
rect 7838 6831 7894 6840
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7852 3534 7880 6831
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7288 3188 7340 3194
rect 6656 3148 6868 3176
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6840 3058 6868 3148
rect 7288 3130 7340 3136
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 6932 2650 6960 2994
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6550 2544 6606 2553
rect 6550 2479 6606 2488
rect 6564 2106 6592 2479
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6748 1494 6776 2382
rect 7024 2310 7052 2994
rect 7668 2990 7696 3470
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7194 2408 7250 2417
rect 7194 2343 7250 2352
rect 7208 2310 7236 2343
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 7300 1834 7328 2586
rect 7760 2514 7788 3062
rect 7944 2650 7972 9959
rect 8036 4486 8064 11018
rect 8128 11014 8156 13874
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8220 12850 8248 13398
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 8312 12646 8340 17983
rect 8404 16250 8432 18244
rect 8484 18226 8536 18232
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16250 8524 16594
rect 8392 16244 8444 16250
rect 8392 16186 8444 16192
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8404 13190 8432 13398
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8404 12186 8432 12718
rect 8588 12434 8616 19306
rect 8668 18624 8720 18630
rect 8666 18592 8668 18601
rect 8720 18592 8722 18601
rect 8666 18527 8722 18536
rect 8772 18358 8800 21490
rect 8864 21146 8892 21490
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 8852 21004 8904 21010
rect 8852 20946 8904 20952
rect 8864 20602 8892 20946
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8850 20224 8906 20233
rect 8850 20159 8906 20168
rect 8760 18352 8812 18358
rect 8760 18294 8812 18300
rect 8864 17490 8892 20159
rect 8956 19786 8984 21490
rect 8944 19780 8996 19786
rect 8944 19722 8996 19728
rect 8944 18828 8996 18834
rect 8944 18770 8996 18776
rect 8956 18426 8984 18770
rect 8944 18420 8996 18426
rect 8944 18362 8996 18368
rect 8772 17462 8892 17490
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 16114 8708 17138
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8680 15026 8708 16050
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8220 12158 8432 12186
rect 8496 12406 8616 12434
rect 8220 11370 8248 12158
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8312 11558 8340 12038
rect 8496 11762 8524 12406
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8496 11642 8524 11698
rect 8404 11614 8524 11642
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8220 11342 8340 11370
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8208 9512 8260 9518
rect 8312 9466 8340 11342
rect 8260 9460 8340 9466
rect 8208 9454 8340 9460
rect 8128 8634 8156 9454
rect 8220 9438 8340 9454
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8312 8129 8340 9438
rect 8298 8120 8354 8129
rect 8298 8055 8354 8064
rect 8298 7848 8354 7857
rect 8404 7834 8432 11614
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 10674 8616 11494
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8484 9920 8536 9926
rect 8680 9908 8708 14758
rect 8772 12782 8800 17462
rect 9048 16182 9076 22170
rect 9128 21684 9180 21690
rect 9128 21626 9180 21632
rect 9140 20097 9168 21626
rect 9220 20596 9272 20602
rect 9220 20538 9272 20544
rect 9126 20088 9182 20097
rect 9126 20023 9182 20032
rect 9140 19514 9168 20023
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 8864 13938 8892 15098
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8772 11558 8800 12582
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8680 9880 8800 9908
rect 8484 9862 8536 9868
rect 8496 8974 8524 9862
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8680 9178 8708 9522
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8496 8514 8524 8910
rect 8496 8486 8616 8514
rect 8588 8430 8616 8486
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8354 7806 8432 7834
rect 8298 7783 8354 7792
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8206 6216 8262 6225
rect 8206 6151 8262 6160
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8128 3534 8156 4014
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8220 3466 8248 6151
rect 8404 5642 8432 6666
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8496 4146 8524 8298
rect 8668 7404 8720 7410
rect 8772 7392 8800 9880
rect 8864 9602 8892 13874
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8956 13394 8984 13738
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 9048 12850 9076 15506
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9140 13530 9168 15438
rect 9232 15076 9260 20538
rect 9324 17542 9352 26318
rect 9416 22982 9444 26846
rect 9508 24857 9536 29056
rect 9692 28994 9720 29396
rect 9600 28966 9720 28994
rect 9600 28558 9628 28966
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9680 28416 9732 28422
rect 9586 28384 9642 28393
rect 9680 28358 9732 28364
rect 9586 28319 9642 28328
rect 9600 28082 9628 28319
rect 9588 28076 9640 28082
rect 9588 28018 9640 28024
rect 9692 27470 9720 28358
rect 9680 27464 9732 27470
rect 9680 27406 9732 27412
rect 9784 27418 9812 29514
rect 9876 28994 9904 29804
rect 9876 28966 10364 28994
rect 9851 28860 10159 28869
rect 9851 28858 9857 28860
rect 9913 28858 9937 28860
rect 9993 28858 10017 28860
rect 10073 28858 10097 28860
rect 10153 28858 10159 28860
rect 9913 28806 9915 28858
rect 10095 28806 10097 28858
rect 9851 28804 9857 28806
rect 9913 28804 9937 28806
rect 9993 28804 10017 28806
rect 10073 28804 10097 28806
rect 10153 28804 10159 28806
rect 9851 28795 10159 28804
rect 10048 28416 10100 28422
rect 9876 28376 10048 28404
rect 9876 28014 9904 28376
rect 10048 28358 10100 28364
rect 10336 28370 10364 28966
rect 10428 28490 10456 30348
rect 10520 29646 10548 30602
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10336 28342 10456 28370
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9968 27962 9996 28154
rect 10428 28082 10456 28342
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 9968 27934 10272 27962
rect 9851 27772 10159 27781
rect 9851 27770 9857 27772
rect 9913 27770 9937 27772
rect 9993 27770 10017 27772
rect 10073 27770 10097 27772
rect 10153 27770 10159 27772
rect 9913 27718 9915 27770
rect 10095 27718 10097 27770
rect 9851 27716 9857 27718
rect 9913 27716 9937 27718
rect 9993 27716 10017 27718
rect 10073 27716 10097 27718
rect 10153 27716 10159 27718
rect 9851 27707 10159 27716
rect 10244 27656 10272 27934
rect 10428 27860 10456 28018
rect 10520 27985 10548 29582
rect 10506 27976 10562 27985
rect 10506 27911 10562 27920
rect 10428 27832 10548 27860
rect 10324 27668 10376 27674
rect 10244 27628 10324 27656
rect 10324 27610 10376 27616
rect 10416 27600 10468 27606
rect 10414 27568 10416 27577
rect 10468 27568 10470 27577
rect 10414 27503 10470 27512
rect 10520 27452 10548 27832
rect 10244 27424 10548 27452
rect 9784 27402 9904 27418
rect 9588 27396 9640 27402
rect 9784 27396 9916 27402
rect 9784 27390 9864 27396
rect 9588 27338 9640 27344
rect 9864 27338 9916 27344
rect 9600 25838 9628 27338
rect 9876 26926 9904 27338
rect 9772 26920 9824 26926
rect 9772 26862 9824 26868
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9692 25770 9720 26454
rect 9784 26432 9812 26862
rect 9851 26684 10159 26693
rect 9851 26682 9857 26684
rect 9913 26682 9937 26684
rect 9993 26682 10017 26684
rect 10073 26682 10097 26684
rect 10153 26682 10159 26684
rect 9913 26630 9915 26682
rect 10095 26630 10097 26682
rect 9851 26628 9857 26630
rect 9913 26628 9937 26630
rect 9993 26628 10017 26630
rect 10073 26628 10097 26630
rect 10153 26628 10159 26630
rect 9851 26619 10159 26628
rect 9956 26444 10008 26450
rect 9784 26404 9956 26432
rect 9956 26386 10008 26392
rect 9968 26058 9996 26386
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10244 26330 10272 27424
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10416 26376 10468 26382
rect 10322 26344 10378 26353
rect 10046 26072 10102 26081
rect 9968 26030 10046 26058
rect 10046 26007 10102 26016
rect 9772 25832 9824 25838
rect 10048 25832 10100 25838
rect 9772 25774 9824 25780
rect 9862 25800 9918 25809
rect 9680 25764 9732 25770
rect 9680 25706 9732 25712
rect 9494 24848 9550 24857
rect 9494 24783 9550 24792
rect 9692 24682 9720 25706
rect 9784 25158 9812 25774
rect 9918 25780 10048 25786
rect 9918 25774 10100 25780
rect 9918 25758 10088 25774
rect 9862 25735 9918 25744
rect 10152 25684 10180 26318
rect 10244 26302 10322 26330
rect 10416 26318 10468 26324
rect 10322 26279 10378 26288
rect 10428 25838 10456 26318
rect 10416 25832 10468 25838
rect 10416 25774 10468 25780
rect 10152 25656 10272 25684
rect 9851 25596 10159 25605
rect 9851 25594 9857 25596
rect 9913 25594 9937 25596
rect 9993 25594 10017 25596
rect 10073 25594 10097 25596
rect 10153 25594 10159 25596
rect 9913 25542 9915 25594
rect 10095 25542 10097 25594
rect 9851 25540 9857 25542
rect 9913 25540 9937 25542
rect 9993 25540 10017 25542
rect 10073 25540 10097 25542
rect 10153 25540 10159 25542
rect 9851 25531 10159 25540
rect 9772 25152 9824 25158
rect 9772 25094 9824 25100
rect 9680 24676 9732 24682
rect 9680 24618 9732 24624
rect 9784 24274 9812 25094
rect 9851 24508 10159 24517
rect 9851 24506 9857 24508
rect 9913 24506 9937 24508
rect 9993 24506 10017 24508
rect 10073 24506 10097 24508
rect 10153 24506 10159 24508
rect 9913 24454 9915 24506
rect 10095 24454 10097 24506
rect 9851 24452 9857 24454
rect 9913 24452 9937 24454
rect 9993 24452 10017 24454
rect 10073 24452 10097 24454
rect 10153 24452 10159 24454
rect 9851 24443 10159 24452
rect 10244 24392 10272 25656
rect 10428 25498 10456 25774
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10322 25392 10378 25401
rect 10322 25327 10378 25336
rect 10336 25294 10364 25327
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10336 24410 10364 24618
rect 10152 24364 10272 24392
rect 10324 24404 10376 24410
rect 9772 24268 9824 24274
rect 9772 24210 9824 24216
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9600 24041 9628 24142
rect 9680 24064 9732 24070
rect 9586 24032 9642 24041
rect 9680 24006 9732 24012
rect 9586 23967 9642 23976
rect 9586 23760 9642 23769
rect 9586 23695 9588 23704
rect 9640 23695 9642 23704
rect 9588 23666 9640 23672
rect 9692 23662 9720 24006
rect 9770 23896 9826 23905
rect 9770 23831 9772 23840
rect 9824 23831 9826 23840
rect 9864 23860 9916 23866
rect 9772 23802 9824 23808
rect 9864 23802 9916 23808
rect 9770 23760 9826 23769
rect 9770 23695 9772 23704
rect 9824 23695 9826 23704
rect 9772 23666 9824 23672
rect 9680 23656 9732 23662
rect 9876 23610 9904 23802
rect 10152 23798 10180 24364
rect 10324 24346 10376 24352
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9680 23598 9732 23604
rect 9784 23582 9904 23610
rect 10138 23624 10194 23633
rect 9678 23488 9734 23497
rect 9678 23423 9734 23432
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9416 20874 9444 22918
rect 9586 22264 9642 22273
rect 9496 22228 9548 22234
rect 9586 22199 9642 22208
rect 9496 22170 9548 22176
rect 9508 21468 9536 22170
rect 9600 22030 9628 22199
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9692 21690 9720 23423
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9784 21570 9812 23582
rect 10138 23559 10140 23568
rect 10192 23559 10194 23568
rect 10140 23530 10192 23536
rect 9851 23420 10159 23429
rect 9851 23418 9857 23420
rect 9913 23418 9937 23420
rect 9993 23418 10017 23420
rect 10073 23418 10097 23420
rect 10153 23418 10159 23420
rect 9913 23366 9915 23418
rect 10095 23366 10097 23418
rect 9851 23364 9857 23366
rect 9913 23364 9937 23366
rect 9993 23364 10017 23366
rect 10073 23364 10097 23366
rect 10153 23364 10159 23366
rect 9851 23355 10159 23364
rect 10138 23216 10194 23225
rect 10138 23151 10194 23160
rect 10152 23050 10180 23151
rect 10140 23044 10192 23050
rect 10140 22986 10192 22992
rect 9851 22332 10159 22341
rect 9851 22330 9857 22332
rect 9913 22330 9937 22332
rect 9993 22330 10017 22332
rect 10073 22330 10097 22332
rect 10153 22330 10159 22332
rect 9913 22278 9915 22330
rect 10095 22278 10097 22330
rect 9851 22276 9857 22278
rect 9913 22276 9937 22278
rect 9993 22276 10017 22278
rect 10073 22276 10097 22278
rect 10153 22276 10159 22278
rect 9851 22267 10159 22276
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9862 21584 9918 21593
rect 9784 21542 9862 21570
rect 9862 21519 9918 21528
rect 9876 21486 9904 21519
rect 9588 21480 9640 21486
rect 9508 21440 9588 21468
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 9508 20618 9536 21440
rect 9588 21422 9640 21428
rect 9864 21480 9916 21486
rect 9864 21422 9916 21428
rect 9968 21332 9996 22170
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21418 10088 21966
rect 10048 21412 10100 21418
rect 10048 21354 10100 21360
rect 9784 21304 9996 21332
rect 9586 21176 9642 21185
rect 9586 21111 9642 21120
rect 9600 20942 9628 21111
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9784 20641 9812 21304
rect 9851 21244 10159 21253
rect 9851 21242 9857 21244
rect 9913 21242 9937 21244
rect 9993 21242 10017 21244
rect 10073 21242 10097 21244
rect 10153 21242 10159 21244
rect 9913 21190 9915 21242
rect 10095 21190 10097 21242
rect 9851 21188 9857 21190
rect 9913 21188 9937 21190
rect 9993 21188 10017 21190
rect 10073 21188 10097 21190
rect 10153 21188 10159 21190
rect 9851 21179 10159 21188
rect 9416 20590 9536 20618
rect 9770 20632 9826 20641
rect 9416 20262 9444 20590
rect 9770 20567 9826 20576
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9324 15570 9352 17478
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9312 15088 9364 15094
rect 9232 15048 9312 15076
rect 9312 15030 9364 15036
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9232 12850 9260 13670
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8942 12744 8998 12753
rect 8942 12679 8998 12688
rect 8956 11830 8984 12679
rect 9048 12170 9076 12786
rect 9324 12646 9352 13806
rect 9312 12640 9364 12646
rect 9312 12582 9364 12588
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 9048 11121 9076 11222
rect 9140 11150 9168 11562
rect 9416 11234 9444 20198
rect 9784 20040 9812 20567
rect 9851 20156 10159 20165
rect 9851 20154 9857 20156
rect 9913 20154 9937 20156
rect 9993 20154 10017 20156
rect 10073 20154 10097 20156
rect 10153 20154 10159 20156
rect 9913 20102 9915 20154
rect 10095 20102 10097 20154
rect 9851 20100 9857 20102
rect 9913 20100 9937 20102
rect 9993 20100 10017 20102
rect 10073 20100 10097 20102
rect 10153 20100 10159 20102
rect 9851 20091 10159 20100
rect 9784 20012 9996 20040
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9692 18714 9720 19110
rect 9508 18698 9720 18714
rect 9496 18692 9720 18698
rect 9548 18686 9720 18692
rect 9496 18634 9548 18640
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9508 18329 9536 18362
rect 9600 18358 9628 18566
rect 9588 18352 9640 18358
rect 9494 18320 9550 18329
rect 9588 18294 9640 18300
rect 9494 18255 9550 18264
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17270 9628 18158
rect 9784 18136 9812 19382
rect 9968 19174 9996 20012
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 19446 10088 19790
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9851 19068 10159 19077
rect 9851 19066 9857 19068
rect 9913 19066 9937 19068
rect 9993 19066 10017 19068
rect 10073 19066 10097 19068
rect 10153 19066 10159 19068
rect 9913 19014 9915 19066
rect 10095 19014 10097 19066
rect 9851 19012 9857 19014
rect 9913 19012 9937 19014
rect 9993 19012 10017 19014
rect 10073 19012 10097 19014
rect 10153 19012 10159 19014
rect 9851 19003 10159 19012
rect 9862 18864 9918 18873
rect 9862 18799 9918 18808
rect 9876 18698 9904 18799
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 10060 18601 10088 18634
rect 10046 18592 10102 18601
rect 10046 18527 10102 18536
rect 9692 18108 9812 18136
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9692 15994 9720 18108
rect 10244 18068 10272 24210
rect 10324 24132 10376 24138
rect 10324 24074 10376 24080
rect 10336 23866 10364 24074
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10336 21350 10364 22578
rect 10428 22030 10456 22918
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10416 21412 10468 21418
rect 10416 21354 10468 21360
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10324 21004 10376 21010
rect 10428 20992 10456 21354
rect 10376 20964 10456 20992
rect 10324 20946 10376 20952
rect 10336 19854 10364 20946
rect 10520 20618 10548 27066
rect 10612 22964 10640 30670
rect 10704 30654 10824 30682
rect 10692 30184 10744 30190
rect 10692 30126 10744 30132
rect 10704 29714 10732 30126
rect 10692 29708 10744 29714
rect 10692 29650 10744 29656
rect 10690 29336 10746 29345
rect 10690 29271 10692 29280
rect 10744 29271 10746 29280
rect 10692 29242 10744 29248
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 10704 25770 10732 28494
rect 10692 25764 10744 25770
rect 10692 25706 10744 25712
rect 10690 24712 10746 24721
rect 10690 24647 10746 24656
rect 10704 23118 10732 24647
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10612 22936 10732 22964
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10612 21486 10640 21830
rect 10704 21690 10732 22936
rect 10692 21684 10744 21690
rect 10692 21626 10744 21632
rect 10600 21480 10652 21486
rect 10600 21422 10652 21428
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10598 21040 10654 21049
rect 10598 20975 10654 20984
rect 10612 20942 10640 20975
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10428 20602 10548 20618
rect 10416 20596 10548 20602
rect 10468 20590 10548 20596
rect 10416 20538 10468 20544
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10322 19408 10378 19417
rect 10322 19343 10324 19352
rect 10376 19343 10378 19352
rect 10324 19314 10376 19320
rect 10324 19168 10376 19174
rect 10428 19156 10456 20538
rect 10508 20528 10560 20534
rect 10508 20470 10560 20476
rect 10520 19938 10548 20470
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10612 20058 10640 20402
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10520 19910 10640 19938
rect 10428 19128 10548 19156
rect 10324 19110 10376 19116
rect 9784 18040 10272 18068
rect 9784 17746 9812 18040
rect 9851 17980 10159 17989
rect 9851 17978 9857 17980
rect 9913 17978 9937 17980
rect 9993 17978 10017 17980
rect 10073 17978 10097 17980
rect 10153 17978 10159 17980
rect 9913 17926 9915 17978
rect 10095 17926 10097 17978
rect 9851 17924 9857 17926
rect 9913 17924 9937 17926
rect 9993 17924 10017 17926
rect 10073 17924 10097 17926
rect 10153 17924 10159 17926
rect 9851 17915 10159 17924
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9864 17740 9916 17746
rect 9864 17682 9916 17688
rect 9784 16726 9812 17682
rect 9876 17542 9904 17682
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 9864 17536 9916 17542
rect 10152 17524 10180 17614
rect 10336 17592 10364 19110
rect 10520 18970 10548 19128
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10612 18737 10640 19910
rect 10598 18728 10654 18737
rect 10598 18663 10654 18672
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 17814 10548 18022
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10612 17660 10640 18566
rect 10704 18358 10732 21286
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10692 17672 10744 17678
rect 10612 17632 10692 17660
rect 10692 17614 10744 17620
rect 10336 17564 10456 17592
rect 10152 17496 10364 17524
rect 9864 17478 9916 17484
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 9851 16892 10159 16901
rect 9851 16890 9857 16892
rect 9913 16890 9937 16892
rect 9993 16890 10017 16892
rect 10073 16890 10097 16892
rect 10153 16890 10159 16892
rect 9913 16838 9915 16890
rect 10095 16838 10097 16890
rect 9851 16836 9857 16838
rect 9913 16836 9937 16838
rect 9993 16836 10017 16838
rect 10073 16836 10097 16838
rect 10153 16836 10159 16838
rect 9851 16827 10159 16836
rect 9772 16720 9824 16726
rect 9772 16662 9824 16668
rect 9770 16552 9826 16561
rect 9770 16487 9826 16496
rect 9784 16114 9812 16487
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9600 15966 9720 15994
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12986 9536 13262
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9232 11206 9444 11234
rect 9128 11144 9180 11150
rect 9034 11112 9090 11121
rect 9128 11086 9180 11092
rect 9034 11047 9090 11056
rect 9232 10690 9260 11206
rect 9312 11144 9364 11150
rect 9600 11132 9628 15966
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15706 9720 15846
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15094 9720 15506
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9784 14600 9812 16050
rect 9851 15804 10159 15813
rect 9851 15802 9857 15804
rect 9913 15802 9937 15804
rect 9993 15802 10017 15804
rect 10073 15802 10097 15804
rect 10153 15802 10159 15804
rect 9913 15750 9915 15802
rect 10095 15750 10097 15802
rect 9851 15748 9857 15750
rect 9913 15748 9937 15750
rect 9993 15748 10017 15750
rect 10073 15748 10097 15750
rect 10153 15748 10159 15750
rect 9851 15739 10159 15748
rect 10244 15620 10272 17138
rect 9862 15600 9918 15609
rect 9862 15535 9918 15544
rect 9968 15592 10272 15620
rect 9876 15502 9904 15535
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9968 15162 9996 15592
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10152 15162 10180 15438
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 9851 14716 10159 14725
rect 9851 14714 9857 14716
rect 9913 14714 9937 14716
rect 9993 14714 10017 14716
rect 10073 14714 10097 14716
rect 10153 14714 10159 14716
rect 9913 14662 9915 14714
rect 10095 14662 10097 14714
rect 9851 14660 9857 14662
rect 9913 14660 9937 14662
rect 9993 14660 10017 14662
rect 10073 14660 10097 14662
rect 10153 14660 10159 14662
rect 9851 14651 10159 14660
rect 9784 14572 9904 14600
rect 9876 13938 9904 14572
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9851 13628 10159 13637
rect 9851 13626 9857 13628
rect 9913 13626 9937 13628
rect 9993 13626 10017 13628
rect 10073 13626 10097 13628
rect 10153 13626 10159 13628
rect 9913 13574 9915 13626
rect 10095 13574 10097 13626
rect 9851 13572 9857 13574
rect 9913 13572 9937 13574
rect 9993 13572 10017 13574
rect 10073 13572 10097 13574
rect 10153 13572 10159 13574
rect 9851 13563 10159 13572
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9968 12986 9996 13194
rect 10152 13172 10180 13330
rect 10244 13240 10272 14962
rect 10336 13410 10364 17496
rect 10428 17202 10456 17564
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17338 10548 17478
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10414 17096 10470 17105
rect 10414 17031 10470 17040
rect 10428 13734 10456 17031
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10520 14618 10548 16934
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 15706 10640 16050
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 10508 13728 10560 13734
rect 10508 13670 10560 13676
rect 10598 13696 10654 13705
rect 10416 13524 10468 13530
rect 10520 13512 10548 13670
rect 10598 13631 10654 13640
rect 10468 13484 10548 13512
rect 10416 13466 10468 13472
rect 10336 13382 10548 13410
rect 10244 13212 10456 13240
rect 10152 13144 10364 13172
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10232 12980 10284 12986
rect 10232 12922 10284 12928
rect 9851 12540 10159 12549
rect 9851 12538 9857 12540
rect 9913 12538 9937 12540
rect 9993 12538 10017 12540
rect 10073 12538 10097 12540
rect 10153 12538 10159 12540
rect 9913 12486 9915 12538
rect 10095 12486 10097 12538
rect 9851 12484 9857 12486
rect 9913 12484 9937 12486
rect 9993 12484 10017 12486
rect 10073 12484 10097 12486
rect 10153 12484 10159 12486
rect 9851 12475 10159 12484
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9692 11218 9720 11494
rect 9680 11212 9732 11218
rect 9784 11200 9812 12378
rect 9851 11452 10159 11461
rect 9851 11450 9857 11452
rect 9913 11450 9937 11452
rect 9993 11450 10017 11452
rect 10073 11450 10097 11452
rect 10153 11450 10159 11452
rect 9913 11398 9915 11450
rect 10095 11398 10097 11450
rect 9851 11396 9857 11398
rect 9913 11396 9937 11398
rect 9993 11396 10017 11398
rect 10073 11396 10097 11398
rect 10153 11396 10159 11398
rect 9851 11387 10159 11396
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 9864 11212 9916 11218
rect 9784 11172 9864 11200
rect 9680 11154 9732 11160
rect 9864 11154 9916 11160
rect 9364 11104 9628 11132
rect 9956 11144 10008 11150
rect 9312 11086 9364 11092
rect 10060 11121 10088 11290
rect 10140 11144 10192 11150
rect 9956 11086 10008 11092
rect 10046 11112 10102 11121
rect 9494 10976 9550 10985
rect 9550 10934 9628 10962
rect 9494 10911 9550 10920
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9232 10674 9444 10690
rect 9232 10668 9456 10674
rect 9232 10662 9404 10668
rect 9404 10610 9456 10616
rect 8864 9574 9352 9602
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9048 9178 9076 9454
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9140 8974 9168 9386
rect 9324 8974 9352 9574
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8720 7364 8800 7392
rect 8668 7346 8720 7352
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6934 9076 7142
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9140 6780 9168 8910
rect 9324 7546 9352 8910
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9048 6752 9168 6780
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8956 6254 8984 6666
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8024 2576 8076 2582
rect 7852 2524 8024 2530
rect 7852 2518 8076 2524
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7852 2502 8064 2518
rect 8588 2514 8616 5578
rect 8944 5160 8996 5166
rect 8944 5102 8996 5108
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8680 4078 8708 4422
rect 8956 4282 8984 5102
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8956 2854 8984 4218
rect 9048 3534 9076 6752
rect 9232 5778 9260 7278
rect 9310 6760 9366 6769
rect 9416 6746 9444 10610
rect 9508 7478 9536 10746
rect 9600 10742 9628 10934
rect 9588 10736 9640 10742
rect 9588 10678 9640 10684
rect 9968 10452 9996 11086
rect 10140 11086 10192 11092
rect 10046 11047 10102 11056
rect 10152 10810 10180 11086
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9784 10424 9996 10452
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 6866 9536 7142
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9366 6718 9444 6746
rect 9310 6695 9366 6704
rect 9508 6458 9536 6802
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9310 5944 9366 5953
rect 9310 5879 9366 5888
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9324 5545 9352 5879
rect 9416 5642 9444 6122
rect 9508 5914 9536 6122
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5710 9628 9862
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9692 8537 9720 9454
rect 9678 8528 9734 8537
rect 9678 8463 9734 8472
rect 9692 7546 9720 8463
rect 9784 7546 9812 10424
rect 9851 10364 10159 10373
rect 9851 10362 9857 10364
rect 9913 10362 9937 10364
rect 9993 10362 10017 10364
rect 10073 10362 10097 10364
rect 10153 10362 10159 10364
rect 9913 10310 9915 10362
rect 10095 10310 10097 10362
rect 9851 10308 9857 10310
rect 9913 10308 9937 10310
rect 9993 10308 10017 10310
rect 10073 10308 10097 10310
rect 10153 10308 10159 10310
rect 9851 10299 10159 10308
rect 10244 9674 10272 12922
rect 10152 9646 10272 9674
rect 10152 9518 10180 9646
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 10336 9466 10364 13144
rect 10428 12850 10456 13212
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10428 12753 10456 12786
rect 10414 12744 10470 12753
rect 10414 12679 10470 12688
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10428 9586 10456 9930
rect 10520 9722 10548 13382
rect 10612 11626 10640 13631
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10704 9722 10732 17614
rect 10796 16114 10824 30654
rect 10888 29850 10916 31146
rect 10980 30190 11008 32864
rect 11072 30870 11100 33526
rect 11242 33008 11298 33017
rect 11348 32978 11376 38286
rect 11440 36174 11468 39918
rect 11716 39506 11744 40462
rect 11704 39500 11756 39506
rect 11704 39442 11756 39448
rect 11716 39098 11744 39442
rect 11704 39092 11756 39098
rect 11704 39034 11756 39040
rect 11520 38888 11572 38894
rect 11520 38830 11572 38836
rect 11532 37874 11560 38830
rect 11704 38548 11756 38554
rect 11704 38490 11756 38496
rect 11520 37868 11572 37874
rect 11520 37810 11572 37816
rect 11428 36168 11480 36174
rect 11480 36116 11560 36122
rect 11428 36110 11560 36116
rect 11440 36094 11560 36110
rect 11428 35760 11480 35766
rect 11428 35702 11480 35708
rect 11242 32943 11298 32952
rect 11336 32972 11388 32978
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 11164 32570 11192 32846
rect 11152 32564 11204 32570
rect 11152 32506 11204 32512
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11164 30920 11192 32166
rect 11256 31754 11284 32943
rect 11336 32914 11388 32920
rect 11348 32366 11376 32914
rect 11336 32360 11388 32366
rect 11336 32302 11388 32308
rect 11256 31726 11376 31754
rect 11244 31680 11296 31686
rect 11244 31622 11296 31628
rect 11256 31113 11284 31622
rect 11242 31104 11298 31113
rect 11242 31039 11298 31048
rect 11164 30892 11284 30920
rect 11060 30864 11112 30870
rect 11060 30806 11112 30812
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11164 30394 11192 30738
rect 11152 30388 11204 30394
rect 11152 30330 11204 30336
rect 10968 30184 11020 30190
rect 10968 30126 11020 30132
rect 10876 29844 10928 29850
rect 10928 29804 11100 29832
rect 10876 29786 10928 29792
rect 11072 29714 11100 29804
rect 11164 29782 11192 30330
rect 11256 30122 11284 30892
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 11152 29776 11204 29782
rect 11152 29718 11204 29724
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 11058 29472 11114 29481
rect 11058 29407 11114 29416
rect 11072 29073 11100 29407
rect 11348 29322 11376 31726
rect 11440 30802 11468 35702
rect 11532 32745 11560 36094
rect 11716 35834 11744 38490
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11610 35320 11666 35329
rect 11610 35255 11612 35264
rect 11664 35255 11666 35264
rect 11612 35226 11664 35232
rect 11610 34504 11666 34513
rect 11610 34439 11666 34448
rect 11624 33046 11652 34439
rect 11716 34105 11744 35770
rect 11808 35601 11836 40666
rect 11888 39976 11940 39982
rect 11888 39918 11940 39924
rect 11900 38486 11928 39918
rect 11980 39364 12032 39370
rect 11980 39306 12032 39312
rect 11888 38480 11940 38486
rect 11888 38422 11940 38428
rect 11794 35592 11850 35601
rect 11794 35527 11850 35536
rect 11808 35290 11836 35527
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 11794 34912 11850 34921
rect 11794 34847 11850 34856
rect 11702 34096 11758 34105
rect 11702 34031 11758 34040
rect 11716 33386 11744 34031
rect 11704 33380 11756 33386
rect 11704 33322 11756 33328
rect 11612 33040 11664 33046
rect 11612 32982 11664 32988
rect 11518 32736 11574 32745
rect 11518 32671 11574 32680
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11532 30802 11560 32302
rect 11716 31754 11744 33322
rect 11624 31726 11744 31754
rect 11428 30796 11480 30802
rect 11428 30738 11480 30744
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11532 30394 11560 30738
rect 11520 30388 11572 30394
rect 11520 30330 11572 30336
rect 11624 29714 11652 31726
rect 11704 31136 11756 31142
rect 11704 31078 11756 31084
rect 11716 30394 11744 31078
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11244 29300 11296 29306
rect 11348 29294 11560 29322
rect 11244 29242 11296 29248
rect 10874 29064 10930 29073
rect 10874 28999 10930 29008
rect 11058 29064 11114 29073
rect 11058 28999 11114 29008
rect 11152 29028 11204 29034
rect 10888 24970 10916 28999
rect 11152 28970 11204 28976
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10980 26586 11008 28494
rect 11072 28082 11100 28902
rect 11164 28762 11192 28970
rect 11152 28756 11204 28762
rect 11152 28698 11204 28704
rect 11150 28384 11206 28393
rect 11150 28319 11206 28328
rect 11164 28150 11192 28319
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11072 26450 11100 27814
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25945 11008 26182
rect 10966 25936 11022 25945
rect 10966 25871 11022 25880
rect 11164 25498 11192 28086
rect 11152 25492 11204 25498
rect 11152 25434 11204 25440
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11072 25158 11100 25230
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 10888 24942 11008 24970
rect 10980 24410 11008 24942
rect 11164 24750 11192 25434
rect 11152 24744 11204 24750
rect 11152 24686 11204 24692
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10874 24304 10930 24313
rect 10874 24239 10930 24248
rect 10888 24206 10916 24239
rect 10876 24200 10928 24206
rect 10876 24142 10928 24148
rect 10888 22234 10916 24142
rect 10980 22574 11008 24346
rect 11256 24154 11284 29242
rect 11336 29164 11388 29170
rect 11336 29106 11388 29112
rect 11348 28558 11376 29106
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11440 28762 11468 28902
rect 11428 28756 11480 28762
rect 11428 28698 11480 28704
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11532 28257 11560 29294
rect 11612 28756 11664 28762
rect 11612 28698 11664 28704
rect 11518 28248 11574 28257
rect 11518 28183 11574 28192
rect 11336 28076 11388 28082
rect 11336 28018 11388 28024
rect 11348 25158 11376 28018
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11440 27470 11468 27814
rect 11518 27704 11574 27713
rect 11518 27639 11574 27648
rect 11532 27470 11560 27639
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11428 26240 11480 26246
rect 11428 26182 11480 26188
rect 11336 25152 11388 25158
rect 11336 25094 11388 25100
rect 11164 24126 11284 24154
rect 11060 23180 11112 23186
rect 11060 23122 11112 23128
rect 11072 22778 11100 23122
rect 11060 22772 11112 22778
rect 11164 22760 11192 24126
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 23118 11284 24006
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11164 22732 11284 22760
rect 11060 22714 11112 22720
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 11060 22568 11112 22574
rect 11256 22556 11284 22732
rect 11348 22574 11376 25094
rect 11060 22510 11112 22516
rect 11164 22528 11284 22556
rect 11336 22568 11388 22574
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10968 21684 11020 21690
rect 10968 21626 11020 21632
rect 10874 21584 10930 21593
rect 10874 21519 10930 21528
rect 10888 19854 10916 21519
rect 10980 21468 11008 21626
rect 11072 21622 11100 22510
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 10980 21440 11100 21468
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10980 20398 11008 20742
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10876 19848 10928 19854
rect 10876 19790 10928 19796
rect 11072 19334 11100 21440
rect 10888 19306 11100 19334
rect 10888 18698 10916 19306
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10888 15994 10916 17478
rect 10980 17338 11008 17614
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 10796 15966 10916 15994
rect 10796 13530 10824 15966
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 10888 14929 10916 14962
rect 10874 14920 10930 14929
rect 10874 14855 10930 14864
rect 10980 14657 11008 15302
rect 10966 14648 11022 14657
rect 10966 14583 11022 14592
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10416 9580 10468 9586
rect 10416 9522 10468 9528
rect 10336 9438 10456 9466
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 9851 9276 10159 9285
rect 9851 9274 9857 9276
rect 9913 9274 9937 9276
rect 9993 9274 10017 9276
rect 10073 9274 10097 9276
rect 10153 9274 10159 9276
rect 9913 9222 9915 9274
rect 10095 9222 10097 9274
rect 9851 9220 9857 9222
rect 9913 9220 9937 9222
rect 9993 9220 10017 9222
rect 10073 9220 10097 9222
rect 10153 9220 10159 9222
rect 9851 9211 10159 9220
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8362 10088 8910
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9851 8188 10159 8197
rect 9851 8186 9857 8188
rect 9913 8186 9937 8188
rect 9993 8186 10017 8188
rect 10073 8186 10097 8188
rect 10153 8186 10159 8188
rect 9913 8134 9915 8186
rect 10095 8134 10097 8186
rect 9851 8132 9857 8134
rect 9913 8132 9937 8134
rect 9993 8132 10017 8134
rect 10073 8132 10097 8134
rect 10153 8132 10159 8134
rect 9851 8123 10159 8132
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9784 7206 9812 7482
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9851 7100 10159 7109
rect 9851 7098 9857 7100
rect 9913 7098 9937 7100
rect 9993 7098 10017 7100
rect 10073 7098 10097 7100
rect 10153 7098 10159 7100
rect 9913 7046 9915 7098
rect 10095 7046 10097 7098
rect 9851 7044 9857 7046
rect 9913 7044 9937 7046
rect 9993 7044 10017 7046
rect 10073 7044 10097 7046
rect 10153 7044 10159 7046
rect 9851 7035 10159 7044
rect 10244 6882 10272 8842
rect 10336 8634 10364 9318
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 9864 6860 9916 6866
rect 9968 6854 10272 6882
rect 10336 6866 10364 7142
rect 9968 6848 9996 6854
rect 9916 6820 9996 6848
rect 9864 6802 9916 6808
rect 9876 6610 9904 6802
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9784 6582 9904 6610
rect 9784 6322 9812 6582
rect 10060 6458 10088 6734
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9876 6322 9904 6394
rect 10244 6338 10272 6854
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9864 6316 9916 6322
rect 10244 6310 10364 6338
rect 9864 6258 9916 6264
rect 9876 6100 9904 6258
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 9784 6072 9904 6100
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9310 5536 9366 5545
rect 9310 5471 9366 5480
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 3534 9168 4422
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9048 3346 9076 3470
rect 9126 3360 9182 3369
rect 9048 3318 9126 3346
rect 9126 3295 9182 3304
rect 9324 3194 9352 4082
rect 9680 4072 9732 4078
rect 9784 4060 9812 6072
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 9864 5704 9916 5710
rect 10048 5704 10100 5710
rect 9864 5646 9916 5652
rect 10046 5672 10048 5681
rect 10100 5672 10102 5681
rect 9876 5234 9904 5646
rect 10046 5607 10102 5616
rect 10244 5370 10272 6190
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10336 5250 10364 6310
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10244 5222 10364 5250
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 10244 4185 10272 5222
rect 10428 4486 10456 9438
rect 10520 9042 10548 9658
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10612 9178 10640 9522
rect 10796 9518 10824 13466
rect 10888 12986 10916 14350
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10980 12986 11008 13262
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12434 11008 12582
rect 10888 12406 11008 12434
rect 10784 9512 10836 9518
rect 10704 9472 10784 9500
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10520 5234 10548 8298
rect 10704 6458 10732 9472
rect 10784 9454 10836 9460
rect 10888 8362 10916 12406
rect 11072 12356 11100 16662
rect 10980 12328 11100 12356
rect 10980 9994 11008 12328
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10980 8072 11008 9454
rect 11058 8936 11114 8945
rect 11058 8871 11114 8880
rect 10888 8044 11008 8072
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10796 6934 10824 7890
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10600 6248 10652 6254
rect 10796 6202 10824 6870
rect 10600 6190 10652 6196
rect 10612 5914 10640 6190
rect 10704 6174 10824 6202
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10612 4214 10640 5238
rect 10416 4208 10468 4214
rect 10230 4176 10286 4185
rect 10416 4150 10468 4156
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10230 4111 10286 4120
rect 9732 4032 9812 4060
rect 10048 4072 10100 4078
rect 9680 4014 9732 4020
rect 10138 4040 10194 4049
rect 10100 4020 10138 4026
rect 10048 4014 10138 4020
rect 10060 3998 10138 4014
rect 10138 3975 10194 3984
rect 9680 3936 9732 3942
rect 9956 3936 10008 3942
rect 9680 3878 9732 3884
rect 9784 3896 9956 3924
rect 9494 3768 9550 3777
rect 9404 3732 9456 3738
rect 9494 3703 9496 3712
rect 9404 3674 9456 3680
rect 9548 3703 9550 3712
rect 9496 3674 9548 3680
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 8576 2508 8628 2514
rect 7852 2446 7880 2502
rect 8576 2450 8628 2456
rect 7656 2440 7708 2446
rect 7392 2400 7656 2428
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 6644 1488 6696 1494
rect 6644 1430 6696 1436
rect 6736 1488 6788 1494
rect 6736 1430 6788 1436
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6550 1320 6606 1329
rect 6276 1012 6328 1018
rect 6276 954 6328 960
rect 5170 54 5304 82
rect 5170 0 5226 54
rect 5446 0 5502 160
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 82 6330 160
rect 6380 82 6408 1294
rect 6460 1284 6512 1290
rect 6550 1255 6606 1264
rect 6460 1226 6512 1232
rect 6274 54 6408 82
rect 6472 82 6500 1226
rect 6564 1222 6592 1255
rect 6552 1216 6604 1222
rect 6552 1158 6604 1164
rect 6550 82 6606 160
rect 6472 54 6606 82
rect 6656 82 6684 1430
rect 6736 1216 6788 1222
rect 6734 1184 6736 1193
rect 6788 1184 6790 1193
rect 6734 1119 6790 1128
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 7300 1000 7328 1498
rect 7116 972 7328 1000
rect 7116 160 7144 972
rect 7392 160 7420 2400
rect 7656 2382 7708 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7932 2440 7984 2446
rect 8208 2440 8260 2446
rect 7932 2382 7984 2388
rect 8036 2400 8208 2428
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7564 2304 7616 2310
rect 7840 2304 7892 2310
rect 7564 2246 7616 2252
rect 7746 2272 7802 2281
rect 7484 1358 7512 2246
rect 7576 2106 7604 2246
rect 7840 2246 7892 2252
rect 7746 2207 7802 2216
rect 7654 2136 7710 2145
rect 7564 2100 7616 2106
rect 7760 2106 7788 2207
rect 7852 2106 7880 2246
rect 7654 2071 7710 2080
rect 7748 2100 7800 2106
rect 7564 2042 7616 2048
rect 7668 1834 7696 2071
rect 7748 2042 7800 2048
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7656 1828 7708 1834
rect 7656 1770 7708 1776
rect 7944 1442 7972 2382
rect 7668 1414 7972 1442
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7472 1216 7524 1222
rect 7472 1158 7524 1164
rect 7484 814 7512 1158
rect 7472 808 7524 814
rect 7472 750 7524 756
rect 7668 160 7696 1414
rect 7932 1352 7984 1358
rect 7930 1320 7932 1329
rect 7984 1320 7986 1329
rect 7930 1255 7986 1264
rect 8036 1170 8064 2400
rect 8760 2440 8812 2446
rect 8208 2382 8260 2388
rect 8482 2408 8538 2417
rect 8538 2366 8708 2394
rect 8760 2382 8812 2388
rect 8482 2343 8538 2352
rect 8208 2304 8260 2310
rect 8114 2272 8170 2281
rect 8208 2246 8260 2252
rect 8300 2304 8352 2310
rect 8484 2304 8536 2310
rect 8300 2246 8352 2252
rect 8390 2272 8446 2281
rect 8114 2207 8170 2216
rect 8128 2106 8156 2207
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 7944 1142 8064 1170
rect 7944 160 7972 1142
rect 8220 160 8248 2246
rect 8312 1358 8340 2246
rect 8484 2246 8536 2252
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8390 2207 8446 2216
rect 8404 2106 8432 2207
rect 8496 2106 8524 2246
rect 8588 2106 8616 2246
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 8484 2100 8536 2106
rect 8484 2042 8536 2048
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8680 2038 8708 2366
rect 8668 2032 8720 2038
rect 8668 1974 8720 1980
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8496 1834 8524 1906
rect 8484 1828 8536 1834
rect 8484 1770 8536 1776
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 8392 1352 8444 1358
rect 8680 1329 8708 1498
rect 8392 1294 8444 1300
rect 8666 1320 8722 1329
rect 6826 82 6882 160
rect 6656 54 6882 82
rect 6274 0 6330 54
rect 6550 0 6606 54
rect 6826 0 6882 54
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8404 134 8432 1294
rect 8666 1255 8722 1264
rect 8772 354 8800 2382
rect 8850 2272 8906 2281
rect 8850 2207 8906 2216
rect 8864 2106 8892 2207
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8956 1970 8984 2790
rect 9232 2530 9260 2790
rect 9048 2502 9260 2530
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 9048 1850 9076 2502
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9218 2408 9274 2417
rect 8864 1834 9076 1850
rect 8852 1828 9076 1834
rect 8904 1822 9076 1828
rect 8852 1770 8904 1776
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 8864 1290 8892 1498
rect 8852 1284 8904 1290
rect 8852 1226 8904 1232
rect 8496 326 8800 354
rect 8496 160 8524 326
rect 9140 218 9168 2382
rect 9218 2343 9274 2352
rect 9232 2038 9260 2343
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9324 490 9352 2994
rect 9416 2038 9444 3674
rect 9692 3670 9720 3878
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9784 3505 9812 3896
rect 9956 3878 10008 3884
rect 10140 3936 10192 3942
rect 10244 3924 10272 4111
rect 10192 3896 10272 3924
rect 10324 3936 10376 3942
rect 10140 3878 10192 3884
rect 10324 3878 10376 3884
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9770 3496 9826 3505
rect 9968 3482 9996 3538
rect 10140 3528 10192 3534
rect 9968 3454 10088 3482
rect 10192 3488 10272 3516
rect 10140 3470 10192 3476
rect 9770 3431 9826 3440
rect 9954 3224 10010 3233
rect 9954 3159 10010 3168
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9494 2680 9550 2689
rect 9494 2615 9496 2624
rect 9548 2615 9550 2624
rect 9496 2586 9548 2592
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9508 1562 9536 2382
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 8772 190 9168 218
rect 9232 462 9352 490
rect 8772 160 8800 190
rect 8392 128 8444 134
rect 8392 70 8444 76
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 82 9090 160
rect 9232 82 9260 462
rect 9600 218 9628 3062
rect 9968 2854 9996 3159
rect 10060 3058 10088 3454
rect 10138 3360 10194 3369
rect 10138 3295 10194 3304
rect 10152 3126 10180 3295
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9876 2310 9904 2382
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9680 1896 9732 1902
rect 9678 1864 9680 1873
rect 9732 1864 9734 1873
rect 9678 1799 9734 1808
rect 9876 1766 9904 2246
rect 10244 2106 10272 3488
rect 10336 3126 10364 3878
rect 10428 3126 10456 4150
rect 10704 4146 10732 6174
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10796 5710 10824 6054
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10888 5370 10916 8044
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 10980 7818 11008 7919
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 11072 5896 11100 8871
rect 11164 7562 11192 22528
rect 11336 22510 11388 22516
rect 11440 21978 11468 26182
rect 11532 25906 11560 27406
rect 11624 27130 11652 28698
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 11716 28150 11744 28494
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11704 27940 11756 27946
rect 11704 27882 11756 27888
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11624 25226 11652 25978
rect 11716 25294 11744 27882
rect 11808 27402 11836 34847
rect 11900 34746 11928 38422
rect 11992 38418 12020 39306
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 11980 38004 12032 38010
rect 11980 37946 12032 37952
rect 11992 35766 12020 37946
rect 11980 35760 12032 35766
rect 11980 35702 12032 35708
rect 12072 35284 12124 35290
rect 12072 35226 12124 35232
rect 11980 35080 12032 35086
rect 12084 35068 12112 35226
rect 12032 35040 12112 35068
rect 11980 35022 12032 35028
rect 11888 34740 11940 34746
rect 11940 34700 12020 34728
rect 11888 34682 11940 34688
rect 11888 33992 11940 33998
rect 11888 33934 11940 33940
rect 11900 32978 11928 33934
rect 11992 33522 12020 34700
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 11900 32026 11928 32914
rect 11992 32434 12020 33458
rect 11980 32428 12032 32434
rect 11980 32370 12032 32376
rect 12084 32314 12112 35040
rect 12164 32904 12216 32910
rect 12162 32872 12164 32881
rect 12216 32872 12218 32881
rect 12162 32807 12218 32816
rect 11992 32286 12112 32314
rect 11888 32020 11940 32026
rect 11888 31962 11940 31968
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11900 29714 11928 30738
rect 11888 29708 11940 29714
rect 11888 29650 11940 29656
rect 11992 28994 12020 32286
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 12084 30802 12112 31622
rect 12176 31414 12204 32807
rect 12164 31408 12216 31414
rect 12164 31350 12216 31356
rect 12164 31136 12216 31142
rect 12164 31078 12216 31084
rect 12072 30796 12124 30802
rect 12072 30738 12124 30744
rect 12070 30696 12126 30705
rect 12070 30631 12126 30640
rect 12084 29170 12112 30631
rect 12176 30598 12204 31078
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 12176 29510 12204 30126
rect 12164 29504 12216 29510
rect 12164 29446 12216 29452
rect 12072 29164 12124 29170
rect 12072 29106 12124 29112
rect 11992 28966 12204 28994
rect 11886 28792 11942 28801
rect 11886 28727 11942 28736
rect 11900 28558 11928 28727
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11900 26382 11928 28358
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11808 26042 11836 26318
rect 11796 26036 11848 26042
rect 11796 25978 11848 25984
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11900 25158 11928 25978
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11610 24984 11666 24993
rect 11610 24919 11666 24928
rect 11624 24818 11652 24919
rect 11520 24812 11572 24818
rect 11520 24754 11572 24760
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11532 24410 11560 24754
rect 11888 24676 11940 24682
rect 11888 24618 11940 24624
rect 11520 24404 11572 24410
rect 11520 24346 11572 24352
rect 11900 24206 11928 24618
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11796 23792 11848 23798
rect 11702 23760 11758 23769
rect 11612 23724 11664 23730
rect 11848 23752 11928 23780
rect 11796 23734 11848 23740
rect 11702 23695 11758 23704
rect 11612 23666 11664 23672
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11256 21950 11468 21978
rect 11256 21894 11284 21950
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 20602 11284 21830
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 11426 20496 11482 20505
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11256 20097 11284 20198
rect 11242 20088 11298 20097
rect 11242 20023 11298 20032
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19310 11284 19790
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11256 18766 11284 19246
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 17270 11284 18702
rect 11348 18154 11376 20470
rect 11426 20431 11428 20440
rect 11480 20431 11482 20440
rect 11428 20402 11480 20408
rect 11336 18148 11388 18154
rect 11336 18090 11388 18096
rect 11348 17746 11376 18090
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11244 17264 11296 17270
rect 11532 17218 11560 23462
rect 11624 22982 11652 23666
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11716 22574 11744 23695
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11704 22568 11756 22574
rect 11808 22545 11836 23054
rect 11704 22510 11756 22516
rect 11794 22536 11850 22545
rect 11794 22471 11850 22480
rect 11612 22432 11664 22438
rect 11612 22374 11664 22380
rect 11624 19854 11652 22374
rect 11702 22128 11758 22137
rect 11702 22063 11758 22072
rect 11716 20942 11744 22063
rect 11900 21962 11928 23752
rect 11992 23662 12020 27814
rect 12072 27396 12124 27402
rect 12072 27338 12124 27344
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12084 22710 12112 27338
rect 12176 26772 12204 28966
rect 12268 27577 12296 42706
rect 12348 40384 12400 40390
rect 12348 40326 12400 40332
rect 12360 39982 12388 40326
rect 12348 39976 12400 39982
rect 12348 39918 12400 39924
rect 12360 38350 12388 39918
rect 12348 38344 12400 38350
rect 12348 38286 12400 38292
rect 12360 38010 12388 38286
rect 12348 38004 12400 38010
rect 12348 37946 12400 37952
rect 12346 37224 12402 37233
rect 12346 37159 12402 37168
rect 12360 35766 12388 37159
rect 12348 35760 12400 35766
rect 12348 35702 12400 35708
rect 12360 34921 12388 35702
rect 12346 34912 12402 34921
rect 12346 34847 12402 34856
rect 12452 33862 12480 42706
rect 12532 41200 12584 41206
rect 12532 41142 12584 41148
rect 12544 40526 12572 41142
rect 12532 40520 12584 40526
rect 12532 40462 12584 40468
rect 12532 40384 12584 40390
rect 12532 40326 12584 40332
rect 12544 39914 12572 40326
rect 12532 39908 12584 39914
rect 12532 39850 12584 39856
rect 12532 38752 12584 38758
rect 12532 38694 12584 38700
rect 12544 38554 12572 38694
rect 12532 38548 12584 38554
rect 12532 38490 12584 38496
rect 12636 38434 12664 43046
rect 13004 42702 13032 43336
rect 13452 43318 13504 43324
rect 13636 43308 13688 43314
rect 13636 43250 13688 43256
rect 12992 42696 13044 42702
rect 12992 42638 13044 42644
rect 13268 42628 13320 42634
rect 13268 42570 13320 42576
rect 12818 42460 13126 42469
rect 12818 42458 12824 42460
rect 12880 42458 12904 42460
rect 12960 42458 12984 42460
rect 13040 42458 13064 42460
rect 13120 42458 13126 42460
rect 12880 42406 12882 42458
rect 13062 42406 13064 42458
rect 12818 42404 12824 42406
rect 12880 42404 12904 42406
rect 12960 42404 12984 42406
rect 13040 42404 13064 42406
rect 13120 42404 13126 42406
rect 12818 42395 13126 42404
rect 12818 41372 13126 41381
rect 12818 41370 12824 41372
rect 12880 41370 12904 41372
rect 12960 41370 12984 41372
rect 13040 41370 13064 41372
rect 13120 41370 13126 41372
rect 12880 41318 12882 41370
rect 13062 41318 13064 41370
rect 12818 41316 12824 41318
rect 12880 41316 12904 41318
rect 12960 41316 12984 41318
rect 13040 41316 13064 41318
rect 13120 41316 13126 41318
rect 12818 41307 13126 41316
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12728 40050 12756 40462
rect 12818 40284 13126 40293
rect 12818 40282 12824 40284
rect 12880 40282 12904 40284
rect 12960 40282 12984 40284
rect 13040 40282 13064 40284
rect 13120 40282 13126 40284
rect 12880 40230 12882 40282
rect 13062 40230 13064 40282
rect 12818 40228 12824 40230
rect 12880 40228 12904 40230
rect 12960 40228 12984 40230
rect 13040 40228 13064 40230
rect 13120 40228 13126 40230
rect 12818 40219 13126 40228
rect 12716 40044 12768 40050
rect 12716 39986 12768 39992
rect 12818 39196 13126 39205
rect 12818 39194 12824 39196
rect 12880 39194 12904 39196
rect 12960 39194 12984 39196
rect 13040 39194 13064 39196
rect 13120 39194 13126 39196
rect 12880 39142 12882 39194
rect 13062 39142 13064 39194
rect 12818 39140 12824 39142
rect 12880 39140 12904 39142
rect 12960 39140 12984 39142
rect 13040 39140 13064 39142
rect 13120 39140 13126 39142
rect 12818 39131 13126 39140
rect 13280 38554 13308 42570
rect 13452 42560 13504 42566
rect 13452 42502 13504 42508
rect 13360 39976 13412 39982
rect 13360 39918 13412 39924
rect 13372 39642 13400 39918
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 12636 38406 12756 38434
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12636 38010 12664 38286
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 12532 36576 12584 36582
rect 12532 36518 12584 36524
rect 12544 36310 12572 36518
rect 12532 36304 12584 36310
rect 12532 36246 12584 36252
rect 12624 35760 12676 35766
rect 12624 35702 12676 35708
rect 12636 34746 12664 35702
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 12440 33856 12492 33862
rect 12440 33798 12492 33804
rect 12532 33448 12584 33454
rect 12622 33416 12678 33425
rect 12584 33396 12622 33402
rect 12532 33390 12622 33396
rect 12544 33374 12622 33390
rect 12622 33351 12678 33360
rect 12530 33280 12586 33289
rect 12360 33238 12530 33266
rect 12360 31822 12388 33238
rect 12530 33215 12586 33224
rect 12532 32904 12584 32910
rect 12452 32864 12532 32892
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12360 31278 12388 31758
rect 12452 31521 12480 32864
rect 12532 32846 12584 32852
rect 12728 31906 12756 38406
rect 12818 38108 13126 38117
rect 12818 38106 12824 38108
rect 12880 38106 12904 38108
rect 12960 38106 12984 38108
rect 13040 38106 13064 38108
rect 13120 38106 13126 38108
rect 12880 38054 12882 38106
rect 13062 38054 13064 38106
rect 12818 38052 12824 38054
rect 12880 38052 12904 38054
rect 12960 38052 12984 38054
rect 13040 38052 13064 38054
rect 13120 38052 13126 38054
rect 12818 38043 13126 38052
rect 12818 37020 13126 37029
rect 12818 37018 12824 37020
rect 12880 37018 12904 37020
rect 12960 37018 12984 37020
rect 13040 37018 13064 37020
rect 13120 37018 13126 37020
rect 12880 36966 12882 37018
rect 13062 36966 13064 37018
rect 12818 36964 12824 36966
rect 12880 36964 12904 36966
rect 12960 36964 12984 36966
rect 13040 36964 13064 36966
rect 13120 36964 13126 36966
rect 12818 36955 13126 36964
rect 13464 36530 13492 42502
rect 13648 42294 13676 43250
rect 13740 42752 13768 44463
rect 14016 43602 14044 44463
rect 14292 43602 14320 44463
rect 14016 43574 14136 43602
rect 14292 43574 14412 43602
rect 13820 43104 13872 43110
rect 13820 43046 13872 43052
rect 13832 42945 13860 43046
rect 13818 42936 13874 42945
rect 13818 42871 13874 42880
rect 13820 42764 13872 42770
rect 13740 42724 13820 42752
rect 13820 42706 13872 42712
rect 14108 42702 14136 43574
rect 14280 43104 14332 43110
rect 14280 43046 14332 43052
rect 14292 42945 14320 43046
rect 14278 42936 14334 42945
rect 14278 42871 14334 42880
rect 14384 42702 14412 43574
rect 14568 43364 14596 44463
rect 14844 43382 14872 44463
rect 14740 43376 14792 43382
rect 14568 43336 14740 43364
rect 14740 43318 14792 43324
rect 14832 43376 14884 43382
rect 14832 43318 14884 43324
rect 14924 43172 14976 43178
rect 14924 43114 14976 43120
rect 14740 43104 14792 43110
rect 14740 43046 14792 43052
rect 14752 42838 14780 43046
rect 14936 42945 14964 43114
rect 14922 42936 14978 42945
rect 14922 42871 14978 42880
rect 14740 42832 14792 42838
rect 14740 42774 14792 42780
rect 15120 42752 15148 44463
rect 15292 43716 15344 43722
rect 15292 43658 15344 43664
rect 15304 43450 15332 43658
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15396 43364 15424 44463
rect 15568 43376 15620 43382
rect 15396 43336 15568 43364
rect 15568 43318 15620 43324
rect 15672 43296 15700 44463
rect 15948 43382 15976 44463
rect 15936 43376 15988 43382
rect 16224 43364 16252 44463
rect 16396 43376 16448 43382
rect 16224 43336 16396 43364
rect 15936 43318 15988 43324
rect 16396 43318 16448 43324
rect 15844 43308 15896 43314
rect 15672 43268 15844 43296
rect 15844 43250 15896 43256
rect 15568 43172 15620 43178
rect 15568 43114 15620 43120
rect 16304 43172 16356 43178
rect 16304 43114 16356 43120
rect 15200 42764 15252 42770
rect 15120 42724 15200 42752
rect 15200 42706 15252 42712
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 14372 42696 14424 42702
rect 14372 42638 14424 42644
rect 15292 42696 15344 42702
rect 15292 42638 15344 42644
rect 14740 42628 14792 42634
rect 14740 42570 14792 42576
rect 14556 42560 14608 42566
rect 14556 42502 14608 42508
rect 13636 42288 13688 42294
rect 13636 42230 13688 42236
rect 14094 40624 14150 40633
rect 14150 40582 14228 40610
rect 14094 40559 14150 40568
rect 13544 40452 13596 40458
rect 13544 40394 13596 40400
rect 13372 36502 13492 36530
rect 12818 35932 13126 35941
rect 12818 35930 12824 35932
rect 12880 35930 12904 35932
rect 12960 35930 12984 35932
rect 13040 35930 13064 35932
rect 13120 35930 13126 35932
rect 12880 35878 12882 35930
rect 13062 35878 13064 35930
rect 12818 35876 12824 35878
rect 12880 35876 12904 35878
rect 12960 35876 12984 35878
rect 13040 35876 13064 35878
rect 13120 35876 13126 35878
rect 12818 35867 13126 35876
rect 12808 35624 12860 35630
rect 12808 35566 12860 35572
rect 12900 35624 12952 35630
rect 12900 35566 12952 35572
rect 12820 35290 12848 35566
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 12912 35086 12940 35566
rect 12992 35488 13044 35494
rect 12992 35430 13044 35436
rect 12900 35080 12952 35086
rect 13004 35057 13032 35430
rect 13174 35184 13230 35193
rect 13174 35119 13230 35128
rect 12900 35022 12952 35028
rect 12990 35048 13046 35057
rect 12912 34950 12940 35022
rect 12990 34983 13046 34992
rect 12900 34944 12952 34950
rect 12900 34886 12952 34892
rect 12818 34844 13126 34853
rect 12818 34842 12824 34844
rect 12880 34842 12904 34844
rect 12960 34842 12984 34844
rect 13040 34842 13064 34844
rect 13120 34842 13126 34844
rect 12880 34790 12882 34842
rect 13062 34790 13064 34842
rect 12818 34788 12824 34790
rect 12880 34788 12904 34790
rect 12960 34788 12984 34790
rect 13040 34788 13064 34790
rect 13120 34788 13126 34790
rect 12818 34779 13126 34788
rect 13188 33862 13216 35119
rect 13266 34640 13322 34649
rect 13266 34575 13322 34584
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 12818 33756 13126 33765
rect 12818 33754 12824 33756
rect 12880 33754 12904 33756
rect 12960 33754 12984 33756
rect 13040 33754 13064 33756
rect 13120 33754 13126 33756
rect 12880 33702 12882 33754
rect 13062 33702 13064 33754
rect 12818 33700 12824 33702
rect 12880 33700 12904 33702
rect 12960 33700 12984 33702
rect 13040 33700 13064 33702
rect 13120 33700 13126 33702
rect 12818 33691 13126 33700
rect 12808 33448 12860 33454
rect 12808 33390 12860 33396
rect 12820 32774 12848 33390
rect 12900 33312 12952 33318
rect 12900 33254 12952 33260
rect 12912 33114 12940 33254
rect 12900 33108 12952 33114
rect 12900 33050 12952 33056
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12818 32668 13126 32677
rect 12818 32666 12824 32668
rect 12880 32666 12904 32668
rect 12960 32666 12984 32668
rect 13040 32666 13064 32668
rect 13120 32666 13126 32668
rect 12880 32614 12882 32666
rect 13062 32614 13064 32666
rect 12818 32612 12824 32614
rect 12880 32612 12904 32614
rect 12960 32612 12984 32614
rect 13040 32612 13064 32614
rect 13120 32612 13126 32614
rect 12818 32603 13126 32612
rect 12636 31878 12756 31906
rect 12532 31816 12584 31822
rect 12636 31793 12664 31878
rect 12532 31758 12584 31764
rect 12622 31784 12678 31793
rect 12438 31512 12494 31521
rect 12438 31447 12494 31456
rect 12348 31272 12400 31278
rect 12348 31214 12400 31220
rect 12360 30938 12388 31214
rect 12440 31204 12492 31210
rect 12440 31146 12492 31152
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 12348 30592 12400 30598
rect 12348 30534 12400 30540
rect 12360 29850 12388 30534
rect 12348 29844 12400 29850
rect 12348 29786 12400 29792
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 12360 27713 12388 29582
rect 12346 27704 12402 27713
rect 12346 27639 12402 27648
rect 12254 27568 12310 27577
rect 12360 27538 12388 27639
rect 12254 27503 12310 27512
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 12256 27328 12308 27334
rect 12256 27270 12308 27276
rect 12268 26926 12296 27270
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12176 26744 12296 26772
rect 12164 26308 12216 26314
rect 12164 26250 12216 26256
rect 12176 25226 12204 26250
rect 12268 25906 12296 26744
rect 12256 25900 12308 25906
rect 12256 25842 12308 25848
rect 12164 25220 12216 25226
rect 12164 25162 12216 25168
rect 12164 24744 12216 24750
rect 12164 24686 12216 24692
rect 12268 24698 12296 25842
rect 12176 24274 12204 24686
rect 12268 24670 12388 24698
rect 12164 24268 12216 24274
rect 12164 24210 12216 24216
rect 12176 23186 12204 24210
rect 12256 24132 12308 24138
rect 12256 24074 12308 24080
rect 12268 23798 12296 24074
rect 12360 24041 12388 24670
rect 12346 24032 12402 24041
rect 12346 23967 12402 23976
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12254 23488 12310 23497
rect 12254 23423 12310 23432
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 11888 21956 11940 21962
rect 11888 21898 11940 21904
rect 11980 21956 12032 21962
rect 11980 21898 12032 21904
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11808 20942 11836 21422
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11716 19718 11744 20402
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11610 19000 11666 19009
rect 11610 18935 11666 18944
rect 11624 18766 11652 18935
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11244 17206 11296 17212
rect 11256 16658 11284 17206
rect 11348 17190 11560 17218
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15434 11284 16050
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 14482 11284 15370
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11256 12889 11284 14418
rect 11242 12880 11298 12889
rect 11242 12815 11298 12824
rect 11256 12714 11284 12815
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11256 11762 11284 12650
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 9722 11284 10610
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11164 7534 11284 7562
rect 11072 5868 11192 5896
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10704 4049 10732 4082
rect 10690 4040 10746 4049
rect 10612 3998 10690 4026
rect 10506 3768 10562 3777
rect 10506 3703 10562 3712
rect 10520 3505 10548 3703
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 9864 1760 9916 1766
rect 9864 1702 9916 1708
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10048 1420 10100 1426
rect 10048 1362 10100 1368
rect 9680 1352 9732 1358
rect 9956 1352 10008 1358
rect 9732 1312 9904 1340
rect 9680 1294 9732 1300
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9784 950 9812 1158
rect 9772 944 9824 950
rect 9772 886 9824 892
rect 9324 190 9628 218
rect 9324 160 9352 190
rect 9876 160 9904 1312
rect 9956 1294 10008 1300
rect 9968 1018 9996 1294
rect 9956 1012 10008 1018
rect 9956 954 10008 960
rect 10060 626 10088 1362
rect 10428 1358 10456 2246
rect 10520 1902 10548 2994
rect 10612 2774 10640 3998
rect 10690 3975 10746 3984
rect 10888 3233 10916 5170
rect 10980 5166 11008 5646
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11072 5545 11100 5578
rect 11058 5536 11114 5545
rect 11058 5471 11114 5480
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10874 3224 10930 3233
rect 10874 3159 10930 3168
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 10784 2984 10836 2990
rect 11072 2961 11100 3062
rect 10784 2926 10836 2932
rect 11058 2952 11114 2961
rect 10612 2746 10732 2774
rect 10704 2514 10732 2746
rect 10796 2650 10824 2926
rect 11058 2887 11114 2896
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11060 2576 11112 2582
rect 11060 2518 11112 2524
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10336 746 10364 1158
rect 10324 740 10376 746
rect 10324 682 10376 688
rect 10060 598 10180 626
rect 10152 160 10180 598
rect 9034 54 9260 82
rect 9034 0 9090 54
rect 9310 0 9366 160
rect 9404 128 9456 134
rect 9586 82 9642 160
rect 9456 76 9642 82
rect 9404 70 9642 76
rect 9416 54 9642 70
rect 9586 0 9642 54
rect 9862 0 9918 160
rect 10138 0 10194 160
rect 10414 82 10470 160
rect 10520 82 10548 1702
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10704 160 10732 1158
rect 10980 160 11008 1702
rect 11072 950 11100 2518
rect 11164 2446 11192 5868
rect 11256 2514 11284 7534
rect 11244 2508 11296 2514
rect 11244 2450 11296 2456
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11060 944 11112 950
rect 11060 886 11112 892
rect 10414 54 10548 82
rect 10414 0 10470 54
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11164 82 11192 1362
rect 11348 1340 11376 17190
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11428 15428 11480 15434
rect 11428 15370 11480 15376
rect 11440 14822 11468 15370
rect 11518 15192 11574 15201
rect 11518 15127 11574 15136
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11532 14414 11560 15127
rect 11624 14464 11652 15438
rect 11716 15434 11744 19314
rect 11900 18873 11928 21898
rect 11992 21690 12020 21898
rect 11980 21684 12032 21690
rect 11980 21626 12032 21632
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11992 20058 12020 20878
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11980 19712 12032 19718
rect 12084 19700 12112 22646
rect 12164 22568 12216 22574
rect 12164 22510 12216 22516
rect 12176 21962 12204 22510
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12032 19672 12112 19700
rect 11980 19654 12032 19660
rect 11886 18864 11942 18873
rect 11886 18799 11942 18808
rect 11796 18352 11848 18358
rect 11794 18320 11796 18329
rect 11848 18320 11850 18329
rect 11794 18255 11850 18264
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11808 15094 11836 18255
rect 11900 17678 11928 18799
rect 11888 17672 11940 17678
rect 11888 17614 11940 17620
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 17066 11928 17478
rect 11888 17060 11940 17066
rect 11888 17002 11940 17008
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11624 14436 11744 14464
rect 11520 14408 11572 14414
rect 11572 14368 11652 14396
rect 11520 14350 11572 14356
rect 11624 13977 11652 14368
rect 11716 14006 11744 14436
rect 11704 14000 11756 14006
rect 11610 13968 11666 13977
rect 11704 13942 11756 13948
rect 11610 13903 11666 13912
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11440 7818 11468 13466
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11612 12096 11664 12102
rect 11808 12084 11836 15030
rect 11900 14958 11928 15302
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11886 14376 11942 14385
rect 11886 14311 11888 14320
rect 11940 14311 11942 14320
rect 11888 14282 11940 14288
rect 11888 12844 11940 12850
rect 11992 12832 12020 19654
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12084 18630 12112 18770
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12176 18290 12204 21558
rect 12268 19378 12296 23423
rect 12360 22574 12388 23967
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 12348 20936 12400 20942
rect 12348 20878 12400 20884
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12268 18358 12296 18566
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12176 17678 12204 18226
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12254 17232 12310 17241
rect 12176 16182 12204 17206
rect 12254 17167 12256 17176
rect 12308 17167 12310 17176
rect 12256 17138 12308 17144
rect 12256 16516 12308 16522
rect 12256 16458 12308 16464
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12268 16028 12296 16458
rect 12176 16000 12296 16028
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12084 14618 12112 14962
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 14272 12124 14278
rect 12176 14260 12204 16000
rect 12360 15706 12388 20878
rect 12452 17921 12480 31146
rect 12544 30938 12572 31758
rect 12622 31719 12678 31728
rect 12818 31580 13126 31589
rect 12818 31578 12824 31580
rect 12880 31578 12904 31580
rect 12960 31578 12984 31580
rect 13040 31578 13064 31580
rect 13120 31578 13126 31580
rect 12880 31526 12882 31578
rect 13062 31526 13064 31578
rect 12818 31524 12824 31526
rect 12880 31524 12904 31526
rect 12960 31524 12984 31526
rect 13040 31524 13064 31526
rect 13120 31524 13126 31526
rect 12818 31515 13126 31524
rect 12532 30932 12584 30938
rect 12532 30874 12584 30880
rect 12532 30796 12584 30802
rect 12532 30738 12584 30744
rect 12544 30258 12572 30738
rect 12818 30492 13126 30501
rect 12818 30490 12824 30492
rect 12880 30490 12904 30492
rect 12960 30490 12984 30492
rect 13040 30490 13064 30492
rect 13120 30490 13126 30492
rect 12880 30438 12882 30490
rect 13062 30438 13064 30490
rect 12818 30436 12824 30438
rect 12880 30436 12904 30438
rect 12960 30436 12984 30438
rect 13040 30436 13064 30438
rect 13120 30436 13126 30438
rect 12818 30427 13126 30436
rect 12532 30252 12584 30258
rect 12532 30194 12584 30200
rect 12544 29102 12572 30194
rect 12624 30116 12676 30122
rect 12624 30058 12676 30064
rect 12636 29578 12664 30058
rect 12716 29640 12768 29646
rect 12714 29608 12716 29617
rect 12768 29608 12770 29617
rect 12624 29572 12676 29578
rect 12714 29543 12770 29552
rect 12624 29514 12676 29520
rect 12818 29404 13126 29413
rect 12818 29402 12824 29404
rect 12880 29402 12904 29404
rect 12960 29402 12984 29404
rect 13040 29402 13064 29404
rect 13120 29402 13126 29404
rect 12880 29350 12882 29402
rect 13062 29350 13064 29402
rect 12818 29348 12824 29350
rect 12880 29348 12904 29350
rect 12960 29348 12984 29350
rect 13040 29348 13064 29350
rect 13120 29348 13126 29350
rect 12818 29339 13126 29348
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 12818 28316 13126 28325
rect 12818 28314 12824 28316
rect 12880 28314 12904 28316
rect 12960 28314 12984 28316
rect 13040 28314 13064 28316
rect 13120 28314 13126 28316
rect 12880 28262 12882 28314
rect 13062 28262 13064 28314
rect 12818 28260 12824 28262
rect 12880 28260 12904 28262
rect 12960 28260 12984 28262
rect 13040 28260 13064 28262
rect 13120 28260 13126 28262
rect 12818 28251 13126 28260
rect 13188 28082 13216 28358
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12624 28008 12676 28014
rect 12624 27950 12676 27956
rect 12992 28008 13044 28014
rect 12992 27950 13044 27956
rect 12532 27532 12584 27538
rect 12532 27474 12584 27480
rect 12544 27130 12572 27474
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12636 27062 12664 27950
rect 13004 27878 13032 27950
rect 12992 27872 13044 27878
rect 12992 27814 13044 27820
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 12624 26240 12676 26246
rect 12624 26182 12676 26188
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25362 12572 25638
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12636 25158 12664 26182
rect 12728 25294 12756 27270
rect 12818 27228 13126 27237
rect 12818 27226 12824 27228
rect 12880 27226 12904 27228
rect 12960 27226 12984 27228
rect 13040 27226 13064 27228
rect 13120 27226 13126 27228
rect 12880 27174 12882 27226
rect 13062 27174 13064 27226
rect 12818 27172 12824 27174
rect 12880 27172 12904 27174
rect 12960 27172 12984 27174
rect 13040 27172 13064 27174
rect 13120 27172 13126 27174
rect 12818 27163 13126 27172
rect 12900 26852 12952 26858
rect 12900 26794 12952 26800
rect 12912 26246 12940 26794
rect 13280 26761 13308 34575
rect 13372 29238 13400 36502
rect 13556 35465 13584 40394
rect 13636 39840 13688 39846
rect 13636 39782 13688 39788
rect 13648 39642 13676 39782
rect 13636 39636 13688 39642
rect 13636 39578 13688 39584
rect 13636 37868 13688 37874
rect 13636 37810 13688 37816
rect 13542 35456 13598 35465
rect 13542 35391 13598 35400
rect 13648 35290 13676 37810
rect 14096 37664 14148 37670
rect 14096 37606 14148 37612
rect 13636 35284 13688 35290
rect 13636 35226 13688 35232
rect 13452 34604 13504 34610
rect 13452 34546 13504 34552
rect 13464 30598 13492 34546
rect 13544 34128 13596 34134
rect 13544 34070 13596 34076
rect 13556 33674 13584 34070
rect 13648 33998 13676 35226
rect 13728 34604 13780 34610
rect 13728 34546 13780 34552
rect 13636 33992 13688 33998
rect 13636 33934 13688 33940
rect 13556 33646 13676 33674
rect 13648 33454 13676 33646
rect 13740 33561 13768 34546
rect 14108 34542 14136 37606
rect 14096 34536 14148 34542
rect 14096 34478 14148 34484
rect 14108 34218 14136 34478
rect 14016 34190 14136 34218
rect 14016 34066 14044 34190
rect 14004 34060 14056 34066
rect 14004 34002 14056 34008
rect 13726 33552 13782 33561
rect 13726 33487 13782 33496
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 13820 33380 13872 33386
rect 13820 33322 13872 33328
rect 13728 32496 13780 32502
rect 13728 32438 13780 32444
rect 13634 31920 13690 31929
rect 13634 31855 13690 31864
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13556 30666 13584 31622
rect 13648 31482 13676 31855
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13544 30660 13596 30666
rect 13544 30602 13596 30608
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13636 29776 13688 29782
rect 13636 29718 13688 29724
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 13360 29232 13412 29238
rect 13360 29174 13412 29180
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13464 26926 13492 29038
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 13266 26752 13322 26761
rect 13266 26687 13322 26696
rect 12900 26240 12952 26246
rect 12900 26182 12952 26188
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 12818 26140 13126 26149
rect 12818 26138 12824 26140
rect 12880 26138 12904 26140
rect 12960 26138 12984 26140
rect 13040 26138 13064 26140
rect 13120 26138 13126 26140
rect 12880 26086 12882 26138
rect 13062 26086 13064 26138
rect 12818 26084 12824 26086
rect 12880 26084 12904 26086
rect 12960 26084 12984 26086
rect 13040 26084 13064 26086
rect 13120 26084 13126 26086
rect 12818 26075 13126 26084
rect 13280 25906 13308 26182
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 12992 25764 13044 25770
rect 12992 25706 13044 25712
rect 13004 25498 13032 25706
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12818 25052 13126 25061
rect 12818 25050 12824 25052
rect 12880 25050 12904 25052
rect 12960 25050 12984 25052
rect 13040 25050 13064 25052
rect 13120 25050 13126 25052
rect 12880 24998 12882 25050
rect 13062 24998 13064 25050
rect 12818 24996 12824 24998
rect 12880 24996 12904 24998
rect 12960 24996 12984 24998
rect 13040 24996 13064 24998
rect 13120 24996 13126 24998
rect 12818 24987 13126 24996
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 12818 23964 13126 23973
rect 12818 23962 12824 23964
rect 12880 23962 12904 23964
rect 12960 23962 12984 23964
rect 13040 23962 13064 23964
rect 13120 23962 13126 23964
rect 12880 23910 12882 23962
rect 13062 23910 13064 23962
rect 12818 23908 12824 23910
rect 12880 23908 12904 23910
rect 12960 23908 12984 23910
rect 13040 23908 13064 23910
rect 13120 23908 13126 23910
rect 12818 23899 13126 23908
rect 13188 23662 13216 24550
rect 13176 23656 13228 23662
rect 13176 23598 13228 23604
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12530 21176 12586 21185
rect 12530 21111 12586 21120
rect 12438 17912 12494 17921
rect 12438 17847 12494 17856
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12452 17202 12480 17478
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12254 15464 12310 15473
rect 12254 15399 12310 15408
rect 12124 14232 12204 14260
rect 12072 14214 12124 14220
rect 11940 12804 12020 12832
rect 11888 12786 11940 12792
rect 11900 12753 11928 12786
rect 11886 12744 11942 12753
rect 11886 12679 11942 12688
rect 12084 12628 12112 14214
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13841 12204 14010
rect 12162 13832 12218 13841
rect 12162 13767 12218 13776
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11664 12056 11836 12084
rect 11900 12600 12112 12628
rect 11612 12038 11664 12044
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10266 11560 10542
rect 11520 10260 11572 10266
rect 11520 10202 11572 10208
rect 11624 9926 11652 12038
rect 11702 10704 11758 10713
rect 11900 10674 11928 12600
rect 12176 12170 12204 13330
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 11702 10639 11758 10648
rect 11888 10668 11940 10674
rect 11716 10062 11744 10639
rect 11888 10610 11940 10616
rect 12084 10606 12112 11766
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11532 8906 11560 9590
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11624 8566 11652 9862
rect 11886 9480 11942 9489
rect 11886 9415 11942 9424
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11532 8090 11560 8366
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11428 7812 11480 7818
rect 11428 7754 11480 7760
rect 11624 6322 11652 8502
rect 11794 8392 11850 8401
rect 11716 8350 11794 8378
rect 11716 8294 11744 8350
rect 11794 8327 11850 8336
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11794 8256 11850 8265
rect 11794 8191 11850 8200
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11518 5944 11574 5953
rect 11518 5879 11574 5888
rect 11532 5710 11560 5879
rect 11520 5704 11572 5710
rect 11440 5664 11520 5692
rect 11440 4593 11468 5664
rect 11520 5646 11572 5652
rect 11426 4584 11482 4593
rect 11426 4519 11482 4528
rect 11440 1494 11468 4519
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11532 3126 11560 4082
rect 11808 3194 11836 8191
rect 11900 7886 11928 9415
rect 11992 8566 12020 9930
rect 12084 9674 12112 10542
rect 12176 9994 12204 12106
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12268 9761 12296 15399
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14618 12388 14962
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12360 13394 12388 14554
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12452 13297 12480 16934
rect 12544 16590 12572 21111
rect 12636 20398 12664 23530
rect 13280 23508 13308 25638
rect 13372 23866 13400 26862
rect 13556 26489 13584 29514
rect 13648 29102 13676 29718
rect 13740 29306 13768 32438
rect 13832 31890 13860 33322
rect 14016 33046 14044 33458
rect 14200 33402 14228 40582
rect 14372 37256 14424 37262
rect 14372 37198 14424 37204
rect 14384 36854 14412 37198
rect 14372 36848 14424 36854
rect 14372 36790 14424 36796
rect 14280 36032 14332 36038
rect 14280 35974 14332 35980
rect 14108 33374 14228 33402
rect 14292 34184 14320 35974
rect 14370 35320 14426 35329
rect 14370 35255 14426 35264
rect 14384 35086 14412 35255
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14372 34196 14424 34202
rect 14292 34156 14372 34184
rect 14004 33040 14056 33046
rect 14004 32982 14056 32988
rect 13912 32972 13964 32978
rect 13912 32914 13964 32920
rect 13924 32570 13952 32914
rect 13912 32564 13964 32570
rect 13912 32506 13964 32512
rect 14108 32008 14136 33374
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14200 32842 14228 33254
rect 14188 32836 14240 32842
rect 14188 32778 14240 32784
rect 14186 32600 14242 32609
rect 14186 32535 14242 32544
rect 14200 32502 14228 32535
rect 14188 32496 14240 32502
rect 14188 32438 14240 32444
rect 14108 31980 14228 32008
rect 13820 31884 13872 31890
rect 13820 31826 13872 31832
rect 13832 30258 13860 31826
rect 14200 31770 14228 31980
rect 14292 31822 14320 34156
rect 14372 34138 14424 34144
rect 14372 33856 14424 33862
rect 14372 33798 14424 33804
rect 14198 31742 14228 31770
rect 14280 31816 14332 31822
rect 14280 31758 14332 31764
rect 14198 31634 14226 31742
rect 14198 31606 14228 31634
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 13924 30802 13952 31282
rect 14004 31136 14056 31142
rect 14004 31078 14056 31084
rect 14016 30802 14044 31078
rect 13912 30796 13964 30802
rect 13912 30738 13964 30744
rect 14004 30796 14056 30802
rect 14004 30738 14056 30744
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 14096 30252 14148 30258
rect 14096 30194 14148 30200
rect 13832 29714 13860 30194
rect 14108 29753 14136 30194
rect 14094 29744 14150 29753
rect 13820 29708 13872 29714
rect 14094 29679 14150 29688
rect 13820 29650 13872 29656
rect 14200 29578 14228 31606
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 13728 28960 13780 28966
rect 13728 28902 13780 28908
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 13634 28112 13690 28121
rect 13634 28047 13690 28056
rect 13648 27334 13676 28047
rect 13740 27878 13768 28902
rect 14108 28558 14136 28902
rect 14384 28558 14412 33798
rect 14476 32502 14504 34886
rect 14464 32496 14516 32502
rect 14464 32438 14516 32444
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14476 31142 14504 31962
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 14096 28552 14148 28558
rect 14096 28494 14148 28500
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 13832 28393 13860 28494
rect 13912 28416 13964 28422
rect 13818 28384 13874 28393
rect 13912 28358 13964 28364
rect 14004 28416 14056 28422
rect 14004 28358 14056 28364
rect 13818 28319 13874 28328
rect 13820 28008 13872 28014
rect 13820 27950 13872 27956
rect 13728 27872 13780 27878
rect 13728 27814 13780 27820
rect 13636 27328 13688 27334
rect 13636 27270 13688 27276
rect 13636 27124 13688 27130
rect 13636 27066 13688 27072
rect 13542 26480 13598 26489
rect 13542 26415 13598 26424
rect 13450 25936 13506 25945
rect 13450 25871 13506 25880
rect 13464 25702 13492 25871
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13648 25650 13676 27066
rect 13740 25838 13768 27814
rect 13832 27402 13860 27950
rect 13924 27878 13952 28358
rect 14016 28082 14044 28358
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 14004 27464 14056 27470
rect 14004 27406 14056 27412
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13832 26994 13860 27338
rect 14016 27130 14044 27406
rect 14004 27124 14056 27130
rect 14004 27066 14056 27072
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 14108 26382 14136 28494
rect 14280 28416 14332 28422
rect 14280 28358 14332 28364
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 14096 26376 14148 26382
rect 14096 26318 14148 26324
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13924 25684 13952 26318
rect 14292 25906 14320 28358
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14004 25900 14056 25906
rect 14280 25900 14332 25906
rect 14056 25860 14136 25888
rect 14004 25842 14056 25848
rect 13924 25656 14044 25684
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13360 23656 13412 23662
rect 13464 23644 13492 25638
rect 13648 25622 13768 25650
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 13412 23616 13492 23644
rect 13360 23598 13412 23604
rect 13188 23480 13308 23508
rect 12818 22876 13126 22885
rect 12818 22874 12824 22876
rect 12880 22874 12904 22876
rect 12960 22874 12984 22876
rect 13040 22874 13064 22876
rect 13120 22874 13126 22876
rect 12880 22822 12882 22874
rect 13062 22822 13064 22874
rect 12818 22820 12824 22822
rect 12880 22820 12904 22822
rect 12960 22820 12984 22822
rect 13040 22820 13064 22822
rect 13120 22820 13126 22822
rect 12818 22811 13126 22820
rect 12818 21788 13126 21797
rect 12818 21786 12824 21788
rect 12880 21786 12904 21788
rect 12960 21786 12984 21788
rect 13040 21786 13064 21788
rect 13120 21786 13126 21788
rect 12880 21734 12882 21786
rect 13062 21734 13064 21786
rect 12818 21732 12824 21734
rect 12880 21732 12904 21734
rect 12960 21732 12984 21734
rect 13040 21732 13064 21734
rect 13120 21732 13126 21734
rect 12818 21723 13126 21732
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12728 20398 12756 20742
rect 12818 20700 13126 20709
rect 12818 20698 12824 20700
rect 12880 20698 12904 20700
rect 12960 20698 12984 20700
rect 13040 20698 13064 20700
rect 13120 20698 13126 20700
rect 12880 20646 12882 20698
rect 13062 20646 13064 20698
rect 12818 20644 12824 20646
rect 12880 20644 12904 20646
rect 12960 20644 12984 20646
rect 13040 20644 13064 20646
rect 13120 20644 13126 20646
rect 12818 20635 13126 20644
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12716 19848 12768 19854
rect 12714 19816 12716 19825
rect 12768 19816 12770 19825
rect 12714 19751 12770 19760
rect 12818 19612 13126 19621
rect 12818 19610 12824 19612
rect 12880 19610 12904 19612
rect 12960 19610 12984 19612
rect 13040 19610 13064 19612
rect 13120 19610 13126 19612
rect 12880 19558 12882 19610
rect 13062 19558 13064 19610
rect 12818 19556 12824 19558
rect 12880 19556 12904 19558
rect 12960 19556 12984 19558
rect 13040 19556 13064 19558
rect 13120 19556 13126 19558
rect 12818 19547 13126 19556
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12624 18352 12676 18358
rect 12624 18294 12676 18300
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12636 15162 12664 18294
rect 12728 18222 12756 19110
rect 12818 18524 13126 18533
rect 12818 18522 12824 18524
rect 12880 18522 12904 18524
rect 12960 18522 12984 18524
rect 13040 18522 13064 18524
rect 13120 18522 13126 18524
rect 12880 18470 12882 18522
rect 13062 18470 13064 18522
rect 12818 18468 12824 18470
rect 12880 18468 12904 18470
rect 12960 18468 12984 18470
rect 13040 18468 13064 18470
rect 13120 18468 13126 18470
rect 12818 18459 13126 18468
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12716 17740 12768 17746
rect 12716 17682 12768 17688
rect 12728 16250 12756 17682
rect 13096 17678 13124 18090
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12818 17436 13126 17445
rect 12818 17434 12824 17436
rect 12880 17434 12904 17436
rect 12960 17434 12984 17436
rect 13040 17434 13064 17436
rect 13120 17434 13126 17436
rect 12880 17382 12882 17434
rect 13062 17382 13064 17434
rect 12818 17380 12824 17382
rect 12880 17380 12904 17382
rect 12960 17380 12984 17382
rect 13040 17380 13064 17382
rect 13120 17380 13126 17382
rect 12818 17371 13126 17380
rect 12818 16348 13126 16357
rect 12818 16346 12824 16348
rect 12880 16346 12904 16348
rect 12960 16346 12984 16348
rect 13040 16346 13064 16348
rect 13120 16346 13126 16348
rect 12880 16294 12882 16346
rect 13062 16294 13064 16346
rect 12818 16292 12824 16294
rect 12880 16292 12904 16294
rect 12960 16292 12984 16294
rect 13040 16292 13064 16294
rect 13120 16292 13126 16294
rect 12818 16283 13126 16292
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12624 15156 12676 15162
rect 12544 15116 12624 15144
rect 12438 13288 12494 13297
rect 12438 13223 12494 13232
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12360 12170 12388 12854
rect 12544 12832 12572 15116
rect 12624 15098 12676 15104
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12636 14074 12664 14350
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12636 12900 12664 13806
rect 12728 13530 12756 16050
rect 12818 15260 13126 15269
rect 12818 15258 12824 15260
rect 12880 15258 12904 15260
rect 12960 15258 12984 15260
rect 13040 15258 13064 15260
rect 13120 15258 13126 15260
rect 12880 15206 12882 15258
rect 13062 15206 13064 15258
rect 12818 15204 12824 15206
rect 12880 15204 12904 15206
rect 12960 15204 12984 15206
rect 13040 15204 13064 15206
rect 13120 15204 13126 15206
rect 12818 15195 13126 15204
rect 13188 15162 13216 23480
rect 13268 23180 13320 23186
rect 13268 23122 13320 23128
rect 13280 21486 13308 23122
rect 13372 22930 13400 23598
rect 13556 23225 13584 24210
rect 13542 23216 13598 23225
rect 13542 23151 13598 23160
rect 13542 22944 13598 22953
rect 13372 22902 13542 22930
rect 13542 22879 13598 22888
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 13372 21010 13400 21966
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13450 21176 13506 21185
rect 13556 21162 13584 21490
rect 13506 21134 13584 21162
rect 13450 21111 13506 21120
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13280 20602 13308 20878
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13372 20466 13400 20946
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13556 20058 13584 20402
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 17762 13308 19790
rect 13372 17921 13400 19994
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13358 17912 13414 17921
rect 13358 17847 13414 17856
rect 13280 17734 13400 17762
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17338 13308 17614
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 16046 13308 16526
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 12818 14172 13126 14181
rect 12818 14170 12824 14172
rect 12880 14170 12904 14172
rect 12960 14170 12984 14172
rect 13040 14170 13064 14172
rect 13120 14170 13126 14172
rect 12880 14118 12882 14170
rect 13062 14118 13064 14170
rect 12818 14116 12824 14118
rect 12880 14116 12904 14118
rect 12960 14116 12984 14118
rect 13040 14116 13064 14118
rect 13120 14116 13126 14118
rect 12818 14107 13126 14116
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12820 13326 12848 14010
rect 13188 13870 13216 14214
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12818 13084 13126 13093
rect 12818 13082 12824 13084
rect 12880 13082 12904 13084
rect 12960 13082 12984 13084
rect 13040 13082 13064 13084
rect 13120 13082 13126 13084
rect 12880 13030 12882 13082
rect 13062 13030 13064 13082
rect 12818 13028 12824 13030
rect 12880 13028 12904 13030
rect 12960 13028 12984 13030
rect 13040 13028 13064 13030
rect 13120 13028 13126 13030
rect 12818 13019 13126 13028
rect 13280 12968 13308 15982
rect 13372 15570 13400 17734
rect 13360 15564 13412 15570
rect 13360 15506 13412 15512
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13372 13938 13400 14486
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13096 12940 13308 12968
rect 12636 12872 12848 12900
rect 12544 12804 12664 12832
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12360 9994 12388 12106
rect 12544 11898 12572 12242
rect 12636 12102 12664 12804
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12238 12756 12582
rect 12820 12238 12848 12872
rect 13096 12434 13124 12940
rect 13096 12406 13216 12434
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12624 12096 12676 12102
rect 12676 12056 12756 12084
rect 12624 12038 12676 12044
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12254 9752 12310 9761
rect 12254 9687 12310 9696
rect 12084 9646 12204 9674
rect 12176 9382 12204 9646
rect 12360 9636 12388 9930
rect 12268 9608 12388 9636
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12084 8090 12112 8434
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7954 12204 9318
rect 12268 8566 12296 9608
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12162 7304 12218 7313
rect 12084 7262 12162 7290
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 4486 11928 6190
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 12084 3641 12112 7262
rect 12162 7239 12218 7248
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5914 12204 6122
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12162 5808 12218 5817
rect 12162 5743 12218 5752
rect 12176 5001 12204 5743
rect 12162 4992 12218 5001
rect 12162 4927 12218 4936
rect 12268 4706 12296 8502
rect 12544 8242 12572 11018
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12636 9722 12664 9998
rect 12728 9926 12756 12056
rect 12818 11996 13126 12005
rect 12818 11994 12824 11996
rect 12880 11994 12904 11996
rect 12960 11994 12984 11996
rect 13040 11994 13064 11996
rect 13120 11994 13126 11996
rect 12880 11942 12882 11994
rect 13062 11942 13064 11994
rect 12818 11940 12824 11942
rect 12880 11940 12904 11942
rect 12960 11940 12984 11942
rect 13040 11940 13064 11942
rect 13120 11940 13126 11942
rect 12818 11931 13126 11940
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12912 11286 12940 11562
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12818 10908 13126 10917
rect 12818 10906 12824 10908
rect 12880 10906 12904 10908
rect 12960 10906 12984 10908
rect 13040 10906 13064 10908
rect 13120 10906 13126 10908
rect 12880 10854 12882 10906
rect 13062 10854 13064 10906
rect 12818 10852 12824 10854
rect 12880 10852 12904 10854
rect 12960 10852 12984 10854
rect 13040 10852 13064 10854
rect 13120 10852 13126 10854
rect 12818 10843 13126 10852
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12624 8492 12676 8498
rect 12728 8480 12756 9862
rect 12818 9820 13126 9829
rect 12818 9818 12824 9820
rect 12880 9818 12904 9820
rect 12960 9818 12984 9820
rect 13040 9818 13064 9820
rect 13120 9818 13126 9820
rect 12880 9766 12882 9818
rect 13062 9766 13064 9818
rect 12818 9764 12824 9766
rect 12880 9764 12904 9766
rect 12960 9764 12984 9766
rect 13040 9764 13064 9766
rect 13120 9764 13126 9766
rect 12818 9755 13126 9764
rect 12818 8732 13126 8741
rect 12818 8730 12824 8732
rect 12880 8730 12904 8732
rect 12960 8730 12984 8732
rect 13040 8730 13064 8732
rect 13120 8730 13126 8732
rect 12880 8678 12882 8730
rect 13062 8678 13064 8730
rect 12818 8676 12824 8678
rect 12880 8676 12904 8678
rect 12960 8676 12984 8678
rect 13040 8676 13064 8678
rect 13120 8676 13126 8678
rect 12818 8667 13126 8676
rect 13188 8650 13216 12406
rect 13372 9110 13400 13874
rect 13464 12434 13492 19790
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13556 17270 13584 19343
rect 13648 19258 13676 24754
rect 13740 23730 13768 25622
rect 13912 24812 13964 24818
rect 13912 24754 13964 24760
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23730 13860 24006
rect 13728 23724 13780 23730
rect 13728 23666 13780 23672
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13726 23352 13782 23361
rect 13726 23287 13782 23296
rect 13740 19378 13768 23287
rect 13832 23186 13860 23462
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13648 19230 13722 19258
rect 13694 18986 13722 19230
rect 13694 18958 13768 18986
rect 13634 18728 13690 18737
rect 13634 18663 13690 18672
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13556 15366 13584 17206
rect 13544 15360 13596 15366
rect 13544 15302 13596 15308
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13556 13904 13584 15098
rect 13648 14550 13676 18663
rect 13740 17202 13768 18958
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13832 18358 13860 18906
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13924 17252 13952 24754
rect 14016 22778 14044 25656
rect 14108 24342 14136 25860
rect 14280 25842 14332 25848
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14096 24336 14148 24342
rect 14096 24278 14148 24284
rect 14292 23526 14320 24686
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14384 23202 14412 27950
rect 14476 24614 14504 30534
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14568 24154 14596 42502
rect 14752 41414 14780 42570
rect 14832 42560 14884 42566
rect 14884 42520 15056 42548
rect 14832 42502 14884 42508
rect 14752 41386 14964 41414
rect 14936 38654 14964 41386
rect 14660 38626 14964 38654
rect 14660 31414 14688 38626
rect 14832 33992 14884 33998
rect 14752 33952 14832 33980
rect 14752 31906 14780 33952
rect 14832 33934 14884 33940
rect 14924 33856 14976 33862
rect 14924 33798 14976 33804
rect 14936 33266 14964 33798
rect 14844 33238 14964 33266
rect 14844 33046 14872 33238
rect 14832 33040 14884 33046
rect 15028 32994 15056 42520
rect 15304 42090 15332 42638
rect 15476 42560 15528 42566
rect 15476 42502 15528 42508
rect 15488 42362 15516 42502
rect 15476 42356 15528 42362
rect 15476 42298 15528 42304
rect 15292 42084 15344 42090
rect 15292 42026 15344 42032
rect 15200 42016 15252 42022
rect 15200 41958 15252 41964
rect 15384 42016 15436 42022
rect 15384 41958 15436 41964
rect 15212 41478 15240 41958
rect 15200 41472 15252 41478
rect 15200 41414 15252 41420
rect 15108 41268 15160 41274
rect 15108 41210 15160 41216
rect 15120 41177 15148 41210
rect 15106 41168 15162 41177
rect 15106 41103 15162 41112
rect 15120 33998 15148 41103
rect 15292 37868 15344 37874
rect 15292 37810 15344 37816
rect 15200 35828 15252 35834
rect 15200 35770 15252 35776
rect 15212 35086 15240 35770
rect 15304 35154 15332 37810
rect 15292 35148 15344 35154
rect 15292 35090 15344 35096
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 15304 34898 15332 35090
rect 15212 34870 15332 34898
rect 15212 34066 15240 34870
rect 15396 34746 15424 41958
rect 15476 41540 15528 41546
rect 15476 41482 15528 41488
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15384 34740 15436 34746
rect 15384 34682 15436 34688
rect 15200 34060 15252 34066
rect 15200 34002 15252 34008
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15212 33454 15240 34002
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 14832 32982 14884 32988
rect 14936 32966 15056 32994
rect 14752 31878 14872 31906
rect 14648 31408 14700 31414
rect 14648 31350 14700 31356
rect 14648 31272 14700 31278
rect 14648 31214 14700 31220
rect 14660 30938 14688 31214
rect 14648 30932 14700 30938
rect 14648 30874 14700 30880
rect 14740 30048 14792 30054
rect 14740 29990 14792 29996
rect 14752 29578 14780 29990
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14752 29170 14780 29514
rect 14740 29164 14792 29170
rect 14740 29106 14792 29112
rect 14752 29050 14780 29106
rect 14660 29022 14780 29050
rect 14660 28014 14688 29022
rect 14738 28520 14794 28529
rect 14738 28455 14794 28464
rect 14752 28150 14780 28455
rect 14740 28144 14792 28150
rect 14740 28086 14792 28092
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14740 27872 14792 27878
rect 14740 27814 14792 27820
rect 14660 27470 14688 27814
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14752 27282 14780 27814
rect 14476 24138 14596 24154
rect 14464 24132 14596 24138
rect 14516 24126 14596 24132
rect 14660 27254 14780 27282
rect 14464 24074 14516 24080
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14476 23497 14504 23666
rect 14462 23488 14518 23497
rect 14462 23423 14518 23432
rect 14384 23174 14504 23202
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 14188 22500 14240 22506
rect 14188 22442 14240 22448
rect 14200 20777 14228 22442
rect 14186 20768 14242 20777
rect 14186 20703 14242 20712
rect 14292 20346 14320 22986
rect 14384 22506 14412 23054
rect 14476 22982 14504 23174
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 20466 14412 21286
rect 14476 20806 14504 22918
rect 14464 20800 14516 20806
rect 14464 20742 14516 20748
rect 14372 20460 14424 20466
rect 14424 20420 14504 20448
rect 14372 20402 14424 20408
rect 14108 20318 14320 20346
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14016 19446 14044 19994
rect 14004 19440 14056 19446
rect 14004 19382 14056 19388
rect 14016 18290 14044 19382
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13924 17224 14044 17252
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13636 14544 13688 14550
rect 13636 14486 13688 14492
rect 13740 14482 13768 14962
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13544 13898 13596 13904
rect 13544 13840 13596 13846
rect 13636 13864 13688 13870
rect 13556 13258 13584 13840
rect 13636 13806 13688 13812
rect 13648 13530 13676 13806
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 13464 12406 13584 12434
rect 13556 11762 13584 12406
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13188 8622 13308 8650
rect 13372 8634 13400 9046
rect 13176 8560 13228 8566
rect 13176 8502 13228 8508
rect 12676 8452 12756 8480
rect 12624 8434 12676 8440
rect 12360 8214 12572 8242
rect 12360 5370 12388 8214
rect 12636 8090 12664 8434
rect 12714 8392 12770 8401
rect 12714 8327 12770 8336
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12452 6458 12480 8026
rect 12440 6452 12492 6458
rect 12728 6440 12756 8327
rect 12818 7644 13126 7653
rect 12818 7642 12824 7644
rect 12880 7642 12904 7644
rect 12960 7642 12984 7644
rect 13040 7642 13064 7644
rect 13120 7642 13126 7644
rect 12880 7590 12882 7642
rect 13062 7590 13064 7642
rect 12818 7588 12824 7590
rect 12880 7588 12904 7590
rect 12960 7588 12984 7590
rect 13040 7588 13064 7590
rect 13120 7588 13126 7590
rect 12818 7579 13126 7588
rect 13188 7478 13216 8502
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 12806 6896 12862 6905
rect 12806 6831 12862 6840
rect 12820 6798 12848 6831
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 12440 6394 12492 6400
rect 12544 6412 12756 6440
rect 12544 6322 12572 6412
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12452 5846 12480 6054
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4826 12388 4966
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12268 4678 12388 4706
rect 12254 4040 12310 4049
rect 12254 3975 12310 3984
rect 12070 3632 12126 3641
rect 12070 3567 12126 3576
rect 12084 3194 12112 3567
rect 12268 3466 12296 3975
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12162 3224 12218 3233
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 12072 3188 12124 3194
rect 12162 3159 12218 3168
rect 12072 3130 12124 3136
rect 12176 3126 12204 3159
rect 11520 3120 11572 3126
rect 11520 3062 11572 3068
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 12164 2984 12216 2990
rect 12216 2932 12296 2938
rect 12164 2926 12296 2932
rect 12176 2910 12296 2926
rect 11888 2848 11940 2854
rect 11940 2796 12204 2802
rect 11888 2790 12204 2796
rect 11900 2774 12204 2790
rect 12176 2446 12204 2774
rect 12268 2650 12296 2910
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12360 2530 12388 4678
rect 12544 4604 12572 5646
rect 12636 5137 12664 6054
rect 12728 5914 12756 6258
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 13188 5250 13216 7414
rect 13280 6730 13308 8622
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13556 8498 13584 11698
rect 13648 11642 13676 13194
rect 13740 12918 13768 14418
rect 13832 13326 13860 16050
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13924 14074 13952 14894
rect 13912 14068 13964 14074
rect 13912 14010 13964 14016
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 12912 13780 12918
rect 13728 12854 13780 12860
rect 13818 12880 13874 12889
rect 13818 12815 13874 12824
rect 13832 12782 13860 12815
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 14016 12434 14044 17224
rect 14108 16454 14136 20318
rect 14188 20256 14240 20262
rect 14240 20216 14412 20244
rect 14188 20198 14240 20204
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14200 19514 14228 19858
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19514 14320 19654
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14280 19508 14332 19514
rect 14280 19450 14332 19456
rect 14200 18834 14228 19450
rect 14188 18828 14240 18834
rect 14188 18770 14240 18776
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 14292 18086 14320 18702
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14292 17882 14320 18022
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14096 16448 14148 16454
rect 14148 16408 14228 16436
rect 14096 16390 14148 16396
rect 14096 15428 14148 15434
rect 14096 15370 14148 15376
rect 14108 15026 14136 15370
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14016 12406 14136 12434
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13924 11898 13952 12242
rect 14004 12164 14056 12170
rect 14004 12106 14056 12112
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14016 11778 14044 12106
rect 13924 11750 14044 11778
rect 13648 11614 13768 11642
rect 13636 10736 13688 10742
rect 13636 10678 13688 10684
rect 13648 8566 13676 10678
rect 13740 9994 13768 11614
rect 13924 10674 13952 11750
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13636 8560 13688 8566
rect 13636 8502 13688 8508
rect 13544 8492 13596 8498
rect 13924 8480 13952 10610
rect 14016 10266 14044 10610
rect 14004 10260 14056 10266
rect 14004 10202 14056 10208
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9450 14044 9998
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 14016 9110 14044 9386
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 14004 8492 14056 8498
rect 13924 8452 14004 8480
rect 13544 8434 13596 8440
rect 14004 8434 14056 8440
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13372 7546 13400 7890
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13464 7002 13492 7278
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13280 6186 13308 6666
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13372 6089 13400 6258
rect 13358 6080 13414 6089
rect 13358 6015 13414 6024
rect 13096 5234 13216 5250
rect 13084 5228 13216 5234
rect 13136 5222 13216 5228
rect 13084 5170 13136 5176
rect 12622 5128 12678 5137
rect 12622 5063 12678 5072
rect 13360 5092 13412 5098
rect 13360 5034 13412 5040
rect 13372 4826 13400 5034
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13556 4622 13584 8434
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13832 8090 13860 8366
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13634 7576 13690 7585
rect 14016 7546 14044 8434
rect 13634 7511 13690 7520
rect 14004 7540 14056 7546
rect 12624 4616 12676 4622
rect 12544 4576 12624 4604
rect 12808 4616 12860 4622
rect 12624 4558 12676 4564
rect 12728 4576 12808 4604
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12544 3602 12572 3878
rect 12532 3596 12584 3602
rect 12532 3538 12584 3544
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12532 3460 12584 3466
rect 12636 3448 12664 4558
rect 12728 4146 12756 4576
rect 12808 4558 12860 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 13648 4264 13676 7511
rect 14004 7482 14056 7488
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13924 6458 13952 7346
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13924 5370 13952 5578
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13832 5166 13860 5306
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13464 4236 13676 4264
rect 13358 4176 13414 4185
rect 12716 4140 12768 4146
rect 13358 4111 13414 4120
rect 12716 4082 12768 4088
rect 13372 3738 13400 4111
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 12900 3460 12952 3466
rect 12636 3420 12900 3448
rect 12532 3402 12584 3408
rect 12900 3402 12952 3408
rect 12452 3194 12480 3402
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12544 2582 12572 3402
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 12268 2502 12388 2530
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12072 2440 12124 2446
rect 11794 2408 11850 2417
rect 12072 2382 12124 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 11794 2343 11850 2352
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11624 2106 11652 2246
rect 11612 2100 11664 2106
rect 11612 2042 11664 2048
rect 11716 2038 11744 2246
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11808 1970 11836 2343
rect 12084 2009 12112 2382
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 12070 2000 12126 2009
rect 11796 1964 11848 1970
rect 12070 1935 12126 1944
rect 11796 1906 11848 1912
rect 11796 1760 11848 1766
rect 12072 1760 12124 1766
rect 11796 1702 11848 1708
rect 11900 1720 12072 1748
rect 11428 1488 11480 1494
rect 11428 1430 11480 1436
rect 11808 1358 11836 1702
rect 11704 1352 11756 1358
rect 11348 1312 11704 1340
rect 11704 1294 11756 1300
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11256 678 11284 1158
rect 11900 898 11928 1720
rect 12072 1702 12124 1708
rect 12176 1358 12204 2246
rect 12164 1352 12216 1358
rect 12164 1294 12216 1300
rect 12268 950 12296 2502
rect 12636 2446 12664 3295
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 13464 2774 13492 4236
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13740 3534 13768 3975
rect 13924 3738 13952 5102
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 12728 2746 13492 2774
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 12452 2106 12480 2246
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 12440 1760 12492 1766
rect 12440 1702 12492 1708
rect 12452 1358 12480 1702
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 11808 870 11928 898
rect 12256 944 12308 950
rect 12256 886 12308 892
rect 11336 740 11388 746
rect 11388 700 11560 728
rect 11336 682 11388 688
rect 11244 672 11296 678
rect 11244 614 11296 620
rect 11532 160 11560 700
rect 11808 160 11836 870
rect 12072 672 12124 678
rect 12072 614 12124 620
rect 12084 160 12112 614
rect 12360 160 12388 1158
rect 12544 1018 12572 2246
rect 12622 2136 12678 2145
rect 12728 2122 12756 2746
rect 12898 2680 12954 2689
rect 12898 2615 12954 2624
rect 12912 2446 12940 2615
rect 12900 2440 12952 2446
rect 13268 2440 13320 2446
rect 12900 2382 12952 2388
rect 13266 2408 13268 2417
rect 13320 2408 13322 2417
rect 13266 2343 13322 2352
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 12678 2094 12756 2122
rect 13556 2106 13584 3334
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13544 2100 13596 2106
rect 12622 2071 12678 2080
rect 13544 2042 13596 2048
rect 13542 2000 13598 2009
rect 13542 1935 13544 1944
rect 13596 1935 13598 1944
rect 13544 1906 13596 1912
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 12532 1012 12584 1018
rect 12532 954 12584 960
rect 12636 160 12664 1702
rect 13648 1358 13676 1702
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 12716 1284 12768 1290
rect 12716 1226 12768 1232
rect 12728 626 12756 1226
rect 13084 1216 13136 1222
rect 13452 1216 13504 1222
rect 13136 1176 13216 1204
rect 13084 1158 13136 1164
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12728 598 12940 626
rect 12912 160 12940 598
rect 13188 160 13216 1176
rect 13452 1158 13504 1164
rect 13464 160 13492 1158
rect 13740 160 13768 1498
rect 13832 1358 13860 2790
rect 14108 2514 14136 12406
rect 14200 12102 14228 16408
rect 14278 14648 14334 14657
rect 14278 14583 14334 14592
rect 14292 14074 14320 14583
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 10742 14228 12038
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 8498 14320 10610
rect 14384 9722 14412 20216
rect 14476 19378 14504 20420
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14464 19168 14516 19174
rect 14464 19110 14516 19116
rect 14476 18902 14504 19110
rect 14464 18896 14516 18902
rect 14464 18838 14516 18844
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14476 17105 14504 18226
rect 14568 17270 14596 24006
rect 14660 20466 14688 27254
rect 14844 26330 14872 31878
rect 14936 31210 14964 32966
rect 15304 32910 15332 34682
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15396 33658 15424 33866
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15488 33289 15516 41482
rect 15580 41414 15608 43114
rect 15660 43104 15712 43110
rect 15660 43046 15712 43052
rect 15672 42945 15700 43046
rect 15785 43004 16093 43013
rect 15785 43002 15791 43004
rect 15847 43002 15871 43004
rect 15927 43002 15951 43004
rect 16007 43002 16031 43004
rect 16087 43002 16093 43004
rect 15847 42950 15849 43002
rect 16029 42950 16031 43002
rect 15785 42948 15791 42950
rect 15847 42948 15871 42950
rect 15927 42948 15951 42950
rect 16007 42948 16031 42950
rect 16087 42948 16093 42950
rect 15658 42936 15714 42945
rect 15785 42939 16093 42948
rect 15658 42871 15714 42880
rect 15844 42560 15896 42566
rect 15844 42502 15896 42508
rect 15856 42294 15884 42502
rect 15844 42288 15896 42294
rect 15844 42230 15896 42236
rect 16120 42084 16172 42090
rect 16120 42026 16172 42032
rect 15785 41916 16093 41925
rect 15785 41914 15791 41916
rect 15847 41914 15871 41916
rect 15927 41914 15951 41916
rect 16007 41914 16031 41916
rect 16087 41914 16093 41916
rect 15847 41862 15849 41914
rect 16029 41862 16031 41914
rect 15785 41860 15791 41862
rect 15847 41860 15871 41862
rect 15927 41860 15951 41862
rect 16007 41860 16031 41862
rect 16087 41860 16093 41862
rect 15785 41851 16093 41860
rect 15580 41386 15700 41414
rect 15566 36680 15622 36689
rect 15566 36615 15622 36624
rect 15474 33280 15530 33289
rect 15474 33215 15530 33224
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 15292 32904 15344 32910
rect 15292 32846 15344 32852
rect 15028 32609 15056 32846
rect 15200 32768 15252 32774
rect 15200 32710 15252 32716
rect 15384 32768 15436 32774
rect 15384 32710 15436 32716
rect 15014 32600 15070 32609
rect 15212 32570 15240 32710
rect 15396 32570 15424 32710
rect 15014 32535 15070 32544
rect 15200 32564 15252 32570
rect 15028 31906 15056 32535
rect 15200 32506 15252 32512
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15212 32366 15240 32506
rect 15580 32450 15608 36615
rect 15396 32422 15608 32450
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15200 32360 15252 32366
rect 15200 32302 15252 32308
rect 15120 32026 15148 32302
rect 15108 32020 15160 32026
rect 15108 31962 15160 31968
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 15198 31920 15254 31929
rect 15028 31878 15198 31906
rect 15198 31855 15254 31864
rect 15304 31822 15332 31962
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15108 31408 15160 31414
rect 15108 31350 15160 31356
rect 14924 31204 14976 31210
rect 14924 31146 14976 31152
rect 15120 31113 15148 31350
rect 15106 31104 15162 31113
rect 15106 31039 15162 31048
rect 15108 30796 15160 30802
rect 15028 30756 15108 30784
rect 14924 30048 14976 30054
rect 14924 29990 14976 29996
rect 14936 29102 14964 29990
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14924 28212 14976 28218
rect 14924 28154 14976 28160
rect 14936 27878 14964 28154
rect 15028 27985 15056 30756
rect 15108 30738 15160 30744
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15120 29170 15148 29446
rect 15212 29238 15240 29446
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15014 27976 15070 27985
rect 15014 27911 15070 27920
rect 14924 27872 14976 27878
rect 14924 27814 14976 27820
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 14936 26994 14964 27270
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14752 26302 14872 26330
rect 14752 25684 14780 26302
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14844 26042 14872 26182
rect 14832 26036 14884 26042
rect 14832 25978 14884 25984
rect 14832 25696 14884 25702
rect 14752 25656 14832 25684
rect 14832 25638 14884 25644
rect 14844 23118 14872 25638
rect 14936 24274 14964 26930
rect 15028 26042 15056 27270
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15120 24274 15148 29106
rect 15304 28558 15332 30670
rect 15396 29345 15424 32422
rect 15476 32360 15528 32366
rect 15476 32302 15528 32308
rect 15488 31890 15516 32302
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 32026 15608 32166
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15382 29336 15438 29345
rect 15382 29271 15438 29280
rect 15488 29186 15516 31826
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15580 30802 15608 31758
rect 15568 30796 15620 30802
rect 15568 30738 15620 30744
rect 15396 29158 15516 29186
rect 15568 29164 15620 29170
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15200 28008 15252 28014
rect 15200 27950 15252 27956
rect 15212 27334 15240 27950
rect 15304 27606 15332 28494
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15212 27062 15240 27270
rect 15200 27056 15252 27062
rect 15200 26998 15252 27004
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 14936 24070 14964 24210
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22098 14872 22374
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14832 22092 14884 22098
rect 14832 22034 14884 22040
rect 14752 21690 14780 22034
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14740 21684 14792 21690
rect 14740 21626 14792 21632
rect 14844 21146 14872 21830
rect 15120 21350 15148 21966
rect 15212 21706 15240 26318
rect 15304 24274 15332 27406
rect 15396 25430 15424 29158
rect 15568 29106 15620 29112
rect 15580 29073 15608 29106
rect 15566 29064 15622 29073
rect 15476 29028 15528 29034
rect 15566 28999 15622 29008
rect 15476 28970 15528 28976
rect 15384 25424 15436 25430
rect 15384 25366 15436 25372
rect 15488 24818 15516 28970
rect 15580 27470 15608 28999
rect 15568 27464 15620 27470
rect 15568 27406 15620 27412
rect 15672 26908 15700 41386
rect 15785 40828 16093 40837
rect 15785 40826 15791 40828
rect 15847 40826 15871 40828
rect 15927 40826 15951 40828
rect 16007 40826 16031 40828
rect 16087 40826 16093 40828
rect 15847 40774 15849 40826
rect 16029 40774 16031 40826
rect 15785 40772 15791 40774
rect 15847 40772 15871 40774
rect 15927 40772 15951 40774
rect 16007 40772 16031 40774
rect 16087 40772 16093 40774
rect 15785 40763 16093 40772
rect 15785 39740 16093 39749
rect 15785 39738 15791 39740
rect 15847 39738 15871 39740
rect 15927 39738 15951 39740
rect 16007 39738 16031 39740
rect 16087 39738 16093 39740
rect 15847 39686 15849 39738
rect 16029 39686 16031 39738
rect 15785 39684 15791 39686
rect 15847 39684 15871 39686
rect 15927 39684 15951 39686
rect 16007 39684 16031 39686
rect 16087 39684 16093 39686
rect 15785 39675 16093 39684
rect 15785 38652 16093 38661
rect 15785 38650 15791 38652
rect 15847 38650 15871 38652
rect 15927 38650 15951 38652
rect 16007 38650 16031 38652
rect 16087 38650 16093 38652
rect 15847 38598 15849 38650
rect 16029 38598 16031 38650
rect 15785 38596 15791 38598
rect 15847 38596 15871 38598
rect 15927 38596 15951 38598
rect 16007 38596 16031 38598
rect 16087 38596 16093 38598
rect 15785 38587 16093 38596
rect 15785 37564 16093 37573
rect 15785 37562 15791 37564
rect 15847 37562 15871 37564
rect 15927 37562 15951 37564
rect 16007 37562 16031 37564
rect 16087 37562 16093 37564
rect 15847 37510 15849 37562
rect 16029 37510 16031 37562
rect 15785 37508 15791 37510
rect 15847 37508 15871 37510
rect 15927 37508 15951 37510
rect 16007 37508 16031 37510
rect 16087 37508 16093 37510
rect 15785 37499 16093 37508
rect 15785 36476 16093 36485
rect 15785 36474 15791 36476
rect 15847 36474 15871 36476
rect 15927 36474 15951 36476
rect 16007 36474 16031 36476
rect 16087 36474 16093 36476
rect 15847 36422 15849 36474
rect 16029 36422 16031 36474
rect 15785 36420 15791 36422
rect 15847 36420 15871 36422
rect 15927 36420 15951 36422
rect 16007 36420 16031 36422
rect 16087 36420 16093 36422
rect 15785 36411 16093 36420
rect 15785 35388 16093 35397
rect 15785 35386 15791 35388
rect 15847 35386 15871 35388
rect 15927 35386 15951 35388
rect 16007 35386 16031 35388
rect 16087 35386 16093 35388
rect 15847 35334 15849 35386
rect 16029 35334 16031 35386
rect 15785 35332 15791 35334
rect 15847 35332 15871 35334
rect 15927 35332 15951 35334
rect 16007 35332 16031 35334
rect 16087 35332 16093 35334
rect 15785 35323 16093 35332
rect 15785 34300 16093 34309
rect 15785 34298 15791 34300
rect 15847 34298 15871 34300
rect 15927 34298 15951 34300
rect 16007 34298 16031 34300
rect 16087 34298 16093 34300
rect 15847 34246 15849 34298
rect 16029 34246 16031 34298
rect 15785 34244 15791 34246
rect 15847 34244 15871 34246
rect 15927 34244 15951 34246
rect 16007 34244 16031 34246
rect 16087 34244 16093 34246
rect 15785 34235 16093 34244
rect 15785 33212 16093 33221
rect 15785 33210 15791 33212
rect 15847 33210 15871 33212
rect 15927 33210 15951 33212
rect 16007 33210 16031 33212
rect 16087 33210 16093 33212
rect 15847 33158 15849 33210
rect 16029 33158 16031 33210
rect 15785 33156 15791 33158
rect 15847 33156 15871 33158
rect 15927 33156 15951 33158
rect 16007 33156 16031 33158
rect 16087 33156 16093 33158
rect 15785 33147 16093 33156
rect 16132 33114 16160 42026
rect 16316 41154 16344 43114
rect 16500 42786 16528 44463
rect 16776 43364 16804 44463
rect 17052 43450 17080 44463
rect 17328 44010 17356 44463
rect 17328 43982 17448 44010
rect 17040 43444 17092 43450
rect 17040 43386 17092 43392
rect 16856 43376 16908 43382
rect 16776 43336 16856 43364
rect 16856 43318 16908 43324
rect 17420 43246 17448 43982
rect 17500 43648 17552 43654
rect 17500 43590 17552 43596
rect 17408 43240 17460 43246
rect 17408 43182 17460 43188
rect 17512 43110 17540 43590
rect 17604 43330 17632 44463
rect 17880 43466 17908 44463
rect 18156 43602 18184 44463
rect 18432 43874 18460 44463
rect 18432 43858 18644 43874
rect 18432 43852 18656 43858
rect 18432 43846 18604 43852
rect 18604 43794 18656 43800
rect 18708 43738 18736 44463
rect 18432 43710 18736 43738
rect 18984 43738 19012 44463
rect 18984 43710 19196 43738
rect 18156 43574 18368 43602
rect 17880 43450 18184 43466
rect 17880 43444 18196 43450
rect 17880 43438 18144 43444
rect 18144 43386 18196 43392
rect 18236 43376 18288 43382
rect 17604 43324 18236 43330
rect 17604 43318 18288 43324
rect 17604 43302 18276 43318
rect 17776 43172 17828 43178
rect 17776 43114 17828 43120
rect 18236 43172 18288 43178
rect 18236 43114 18288 43120
rect 16856 43104 16908 43110
rect 16856 43046 16908 43052
rect 17500 43104 17552 43110
rect 17500 43046 17552 43052
rect 17592 43104 17644 43110
rect 17592 43046 17644 43052
rect 16868 42906 16896 43046
rect 16856 42900 16908 42906
rect 16856 42842 16908 42848
rect 17132 42832 17184 42838
rect 16500 42758 16620 42786
rect 17132 42774 17184 42780
rect 16592 42702 16620 42758
rect 16488 42696 16540 42702
rect 16488 42638 16540 42644
rect 16580 42696 16632 42702
rect 16580 42638 16632 42644
rect 16396 42084 16448 42090
rect 16396 42026 16448 42032
rect 16408 41721 16436 42026
rect 16500 42022 16528 42638
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 16948 42560 17000 42566
rect 16948 42502 17000 42508
rect 16488 42016 16540 42022
rect 16488 41958 16540 41964
rect 16394 41712 16450 41721
rect 16394 41647 16450 41656
rect 16316 41126 16436 41154
rect 16304 41064 16356 41070
rect 16304 41006 16356 41012
rect 16316 40730 16344 41006
rect 16408 40730 16436 41126
rect 16304 40724 16356 40730
rect 16304 40666 16356 40672
rect 16396 40724 16448 40730
rect 16396 40666 16448 40672
rect 16488 39432 16540 39438
rect 16488 39374 16540 39380
rect 16500 39030 16528 39374
rect 16488 39024 16540 39030
rect 16488 38966 16540 38972
rect 16396 37324 16448 37330
rect 16396 37266 16448 37272
rect 16304 35080 16356 35086
rect 16304 35022 16356 35028
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 16028 32904 16080 32910
rect 16026 32872 16028 32881
rect 16120 32904 16172 32910
rect 16080 32872 16082 32881
rect 16120 32846 16172 32852
rect 16026 32807 16082 32816
rect 15785 32124 16093 32133
rect 15785 32122 15791 32124
rect 15847 32122 15871 32124
rect 15927 32122 15951 32124
rect 16007 32122 16031 32124
rect 16087 32122 16093 32124
rect 15847 32070 15849 32122
rect 16029 32070 16031 32122
rect 15785 32068 15791 32070
rect 15847 32068 15871 32070
rect 15927 32068 15951 32070
rect 16007 32068 16031 32070
rect 16087 32068 16093 32070
rect 15785 32059 16093 32068
rect 16132 31686 16160 32846
rect 16224 31958 16252 33254
rect 16316 32230 16344 35022
rect 16304 32224 16356 32230
rect 16304 32166 16356 32172
rect 16212 31952 16264 31958
rect 16212 31894 16264 31900
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 16120 31136 16172 31142
rect 16120 31078 16172 31084
rect 15785 31036 16093 31045
rect 15785 31034 15791 31036
rect 15847 31034 15871 31036
rect 15927 31034 15951 31036
rect 16007 31034 16031 31036
rect 16087 31034 16093 31036
rect 15847 30982 15849 31034
rect 16029 30982 16031 31034
rect 15785 30980 15791 30982
rect 15847 30980 15871 30982
rect 15927 30980 15951 30982
rect 16007 30980 16031 30982
rect 16087 30980 16093 30982
rect 15785 30971 16093 30980
rect 16132 30938 16160 31078
rect 16120 30932 16172 30938
rect 16120 30874 16172 30880
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 15785 29948 16093 29957
rect 15785 29946 15791 29948
rect 15847 29946 15871 29948
rect 15927 29946 15951 29948
rect 16007 29946 16031 29948
rect 16087 29946 16093 29948
rect 15847 29894 15849 29946
rect 16029 29894 16031 29946
rect 15785 29892 15791 29894
rect 15847 29892 15871 29894
rect 15927 29892 15951 29894
rect 16007 29892 16031 29894
rect 16087 29892 16093 29894
rect 15785 29883 16093 29892
rect 15752 29708 15804 29714
rect 15752 29650 15804 29656
rect 15764 29073 15792 29650
rect 15750 29064 15806 29073
rect 15750 28999 15806 29008
rect 15785 28860 16093 28869
rect 15785 28858 15791 28860
rect 15847 28858 15871 28860
rect 15927 28858 15951 28860
rect 16007 28858 16031 28860
rect 16087 28858 16093 28860
rect 15847 28806 15849 28858
rect 16029 28806 16031 28858
rect 15785 28804 15791 28806
rect 15847 28804 15871 28806
rect 15927 28804 15951 28806
rect 16007 28804 16031 28806
rect 16087 28804 16093 28806
rect 15785 28795 16093 28804
rect 16132 28558 16160 30670
rect 16224 29782 16252 31894
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16316 30598 16344 31282
rect 16304 30592 16356 30598
rect 16304 30534 16356 30540
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16210 29336 16266 29345
rect 16210 29271 16266 29280
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 15785 27772 16093 27781
rect 15785 27770 15791 27772
rect 15847 27770 15871 27772
rect 15927 27770 15951 27772
rect 16007 27770 16031 27772
rect 16087 27770 16093 27772
rect 15847 27718 15849 27770
rect 16029 27718 16031 27770
rect 15785 27716 15791 27718
rect 15847 27716 15871 27718
rect 15927 27716 15951 27718
rect 16007 27716 16031 27718
rect 16087 27716 16093 27718
rect 15785 27707 16093 27716
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15856 27062 15884 27474
rect 15844 27056 15896 27062
rect 15844 26998 15896 27004
rect 15580 26880 15700 26908
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15384 24608 15436 24614
rect 15384 24550 15436 24556
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15304 22098 15332 22918
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15212 21678 15332 21706
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15028 21146 15056 21286
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 15120 21026 15148 21286
rect 15028 20998 15148 21026
rect 14738 20768 14794 20777
rect 14738 20703 14794 20712
rect 14752 20534 14780 20703
rect 14740 20528 14792 20534
rect 14740 20470 14792 20476
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 19854 14688 20402
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14752 19334 14780 20470
rect 14660 19306 14780 19334
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14660 17116 14688 19306
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 14462 17096 14518 17105
rect 14462 17031 14518 17040
rect 14568 17088 14688 17116
rect 14464 16992 14516 16998
rect 14464 16934 14516 16940
rect 14476 16590 14504 16934
rect 14464 16584 14516 16590
rect 14464 16526 14516 16532
rect 14568 16096 14596 17088
rect 14648 16516 14700 16522
rect 14648 16458 14700 16464
rect 14660 16250 14688 16458
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14648 16108 14700 16114
rect 14568 16068 14648 16096
rect 14648 16050 14700 16056
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14556 13864 14608 13870
rect 14660 13818 14688 15098
rect 14752 14550 14780 19110
rect 15028 18834 15056 20998
rect 15108 19780 15160 19786
rect 15108 19722 15160 19728
rect 15120 18834 15148 19722
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 14832 18624 14884 18630
rect 14832 18566 14884 18572
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 14608 13812 14688 13818
rect 14556 13806 14688 13812
rect 14568 13790 14688 13806
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14476 12102 14504 12174
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 10674 14504 12038
rect 14568 11830 14596 13670
rect 14660 12434 14688 13790
rect 14660 12406 14780 12434
rect 14752 12170 14780 12406
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14738 11792 14794 11801
rect 14738 11727 14794 11736
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14752 8922 14780 11727
rect 14660 8894 14780 8922
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14292 8378 14320 8434
rect 14200 8350 14320 8378
rect 14200 7410 14228 8350
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13924 1358 13952 2246
rect 14004 1828 14056 1834
rect 14004 1770 14056 1776
rect 14016 1358 14044 1770
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 14108 1494 14136 1702
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 14004 1352 14056 1358
rect 14004 1294 14056 1300
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14016 160 14044 1158
rect 14200 814 14228 7346
rect 14384 4758 14412 7346
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14568 4826 14596 4966
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14384 3194 14412 3470
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14660 2774 14688 8894
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 7886 14780 8774
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14752 4622 14780 6190
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 4146 14780 4558
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14660 2746 14780 2774
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 14188 808 14240 814
rect 14188 750 14240 756
rect 14292 160 14320 1702
rect 14476 1290 14504 2246
rect 14752 2106 14780 2746
rect 14844 2446 14872 18566
rect 15212 18034 15240 21558
rect 15304 20482 15332 21678
rect 15396 21185 15424 24550
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15382 21176 15438 21185
rect 15382 21111 15384 21120
rect 15436 21111 15438 21120
rect 15384 21082 15436 21088
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15396 20602 15424 20946
rect 15488 20602 15516 22510
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15304 20454 15516 20482
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15304 18426 15332 18702
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15028 18006 15240 18034
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14618 14964 14758
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14922 13968 14978 13977
rect 14922 13903 14924 13912
rect 14976 13903 14978 13912
rect 14924 13874 14976 13880
rect 15028 12918 15056 18006
rect 15396 17954 15424 20334
rect 15212 17926 15424 17954
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12238 14964 12582
rect 15120 12434 15148 15846
rect 15212 15609 15240 17926
rect 15488 17610 15516 20454
rect 15580 19174 15608 26880
rect 15785 26684 16093 26693
rect 15785 26682 15791 26684
rect 15847 26682 15871 26684
rect 15927 26682 15951 26684
rect 16007 26682 16031 26684
rect 16087 26682 16093 26684
rect 15847 26630 15849 26682
rect 16029 26630 16031 26682
rect 15785 26628 15791 26630
rect 15847 26628 15871 26630
rect 15927 26628 15951 26630
rect 16007 26628 16031 26630
rect 16087 26628 16093 26630
rect 15785 26619 16093 26628
rect 15936 26512 15988 26518
rect 15936 26454 15988 26460
rect 15660 26376 15712 26382
rect 15660 26318 15712 26324
rect 15672 26042 15700 26318
rect 15948 26042 15976 26454
rect 16132 26246 16160 28494
rect 16120 26240 16172 26246
rect 16120 26182 16172 26188
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16120 25832 16172 25838
rect 16120 25774 16172 25780
rect 15660 25764 15712 25770
rect 15660 25706 15712 25712
rect 15672 24392 15700 25706
rect 15785 25596 16093 25605
rect 15785 25594 15791 25596
rect 15847 25594 15871 25596
rect 15927 25594 15951 25596
rect 16007 25594 16031 25596
rect 16087 25594 16093 25596
rect 15847 25542 15849 25594
rect 16029 25542 16031 25594
rect 15785 25540 15791 25542
rect 15847 25540 15871 25542
rect 15927 25540 15951 25542
rect 16007 25540 16031 25542
rect 16087 25540 16093 25542
rect 15785 25531 16093 25540
rect 16132 24614 16160 25774
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 15785 24508 16093 24517
rect 15785 24506 15791 24508
rect 15847 24506 15871 24508
rect 15927 24506 15951 24508
rect 16007 24506 16031 24508
rect 16087 24506 16093 24508
rect 15847 24454 15849 24506
rect 16029 24454 16031 24506
rect 15785 24452 15791 24454
rect 15847 24452 15871 24454
rect 15927 24452 15951 24454
rect 16007 24452 16031 24454
rect 16087 24452 16093 24454
rect 15785 24443 16093 24452
rect 15672 24364 15792 24392
rect 15660 24268 15712 24274
rect 15660 24210 15712 24216
rect 15672 23866 15700 24210
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15764 23746 15792 24364
rect 15936 24200 15988 24206
rect 15936 24142 15988 24148
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15948 23866 15976 24142
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 15672 23718 15792 23746
rect 15672 22574 15700 23718
rect 16040 23594 16068 24142
rect 16224 23712 16252 29271
rect 16316 26586 16344 30534
rect 16304 26580 16356 26586
rect 16304 26522 16356 26528
rect 16302 25256 16358 25265
rect 16302 25191 16358 25200
rect 16132 23684 16252 23712
rect 16028 23588 16080 23594
rect 16028 23530 16080 23536
rect 15785 23420 16093 23429
rect 15785 23418 15791 23420
rect 15847 23418 15871 23420
rect 15927 23418 15951 23420
rect 16007 23418 16031 23420
rect 16087 23418 16093 23420
rect 15847 23366 15849 23418
rect 16029 23366 16031 23418
rect 15785 23364 15791 23366
rect 15847 23364 15871 23366
rect 15927 23364 15951 23366
rect 16007 23364 16031 23366
rect 16087 23364 16093 23366
rect 15785 23355 16093 23364
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15672 18714 15700 22510
rect 16040 22420 16068 22714
rect 16132 22545 16160 23684
rect 16212 23588 16264 23594
rect 16212 23530 16264 23536
rect 16118 22536 16174 22545
rect 16118 22471 16174 22480
rect 16040 22392 16160 22420
rect 15785 22332 16093 22341
rect 15785 22330 15791 22332
rect 15847 22330 15871 22332
rect 15927 22330 15951 22332
rect 16007 22330 16031 22332
rect 16087 22330 16093 22332
rect 15847 22278 15849 22330
rect 16029 22278 16031 22330
rect 15785 22276 15791 22278
rect 15847 22276 15871 22278
rect 15927 22276 15951 22278
rect 16007 22276 16031 22278
rect 16087 22276 16093 22278
rect 15785 22267 16093 22276
rect 16132 22030 16160 22392
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16132 21486 16160 21966
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 15785 21244 16093 21253
rect 15785 21242 15791 21244
rect 15847 21242 15871 21244
rect 15927 21242 15951 21244
rect 16007 21242 16031 21244
rect 16087 21242 16093 21244
rect 15847 21190 15849 21242
rect 16029 21190 16031 21242
rect 15785 21188 15791 21190
rect 15847 21188 15871 21190
rect 15927 21188 15951 21190
rect 16007 21188 16031 21190
rect 16087 21188 16093 21190
rect 15785 21179 16093 21188
rect 16132 21010 16160 21286
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 15752 20936 15804 20942
rect 16224 20890 16252 23530
rect 16316 21622 16344 25191
rect 16304 21616 16356 21622
rect 16304 21558 16356 21564
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 15752 20878 15804 20884
rect 15764 20806 15792 20878
rect 16132 20862 16252 20890
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15764 20398 15792 20742
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 16132 20262 16160 20862
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 15785 20156 16093 20165
rect 15785 20154 15791 20156
rect 15847 20154 15871 20156
rect 15927 20154 15951 20156
rect 16007 20154 16031 20156
rect 16087 20154 16093 20156
rect 15847 20102 15849 20154
rect 16029 20102 16031 20154
rect 15785 20100 15791 20102
rect 15847 20100 15871 20102
rect 15927 20100 15951 20102
rect 16007 20100 16031 20102
rect 16087 20100 16093 20102
rect 15785 20091 16093 20100
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 15785 19068 16093 19077
rect 15785 19066 15791 19068
rect 15847 19066 15871 19068
rect 15927 19066 15951 19068
rect 16007 19066 16031 19068
rect 16087 19066 16093 19068
rect 15847 19014 15849 19066
rect 16029 19014 16031 19066
rect 15785 19012 15791 19014
rect 15847 19012 15871 19014
rect 15927 19012 15951 19014
rect 16007 19012 16031 19014
rect 16087 19012 16093 19014
rect 15785 19003 16093 19012
rect 16132 18970 16160 19382
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15580 18686 15700 18714
rect 16224 18714 16252 20538
rect 16316 20466 16344 20946
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 16316 20058 16344 20402
rect 16304 20052 16356 20058
rect 16408 20040 16436 37266
rect 16500 35272 16528 38966
rect 16672 38820 16724 38826
rect 16672 38762 16724 38768
rect 16684 36786 16712 38762
rect 16776 37330 16804 42502
rect 16960 42294 16988 42502
rect 16948 42288 17000 42294
rect 16948 42230 17000 42236
rect 16856 42016 16908 42022
rect 16856 41958 16908 41964
rect 16868 39001 16896 41958
rect 16854 38992 16910 39001
rect 16854 38927 16910 38936
rect 17144 38758 17172 42774
rect 17604 42702 17632 43046
rect 17788 42702 17816 43114
rect 17868 43104 17920 43110
rect 17868 43046 17920 43052
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 17880 42906 17908 43046
rect 17868 42900 17920 42906
rect 17868 42842 17920 42848
rect 18064 42702 18092 43046
rect 18144 42900 18196 42906
rect 18144 42842 18196 42848
rect 17592 42696 17644 42702
rect 17592 42638 17644 42644
rect 17776 42696 17828 42702
rect 17776 42638 17828 42644
rect 18052 42696 18104 42702
rect 18052 42638 18104 42644
rect 17224 42560 17276 42566
rect 17224 42502 17276 42508
rect 17316 42560 17368 42566
rect 17316 42502 17368 42508
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 18052 42560 18104 42566
rect 18052 42502 18104 42508
rect 17236 42362 17264 42502
rect 17328 42362 17356 42502
rect 17788 42362 17816 42502
rect 18064 42362 18092 42502
rect 17224 42356 17276 42362
rect 17224 42298 17276 42304
rect 17316 42356 17368 42362
rect 17316 42298 17368 42304
rect 17776 42356 17828 42362
rect 17776 42298 17828 42304
rect 18052 42356 18104 42362
rect 18052 42298 18104 42304
rect 18156 42294 18184 42842
rect 18144 42288 18196 42294
rect 18144 42230 18196 42236
rect 17316 42084 17368 42090
rect 17316 42026 17368 42032
rect 17328 41857 17356 42026
rect 17592 42016 17644 42022
rect 17592 41958 17644 41964
rect 18144 42016 18196 42022
rect 18144 41958 18196 41964
rect 17314 41848 17370 41857
rect 17314 41783 17370 41792
rect 17604 41721 17632 41958
rect 17960 41812 18012 41818
rect 17960 41754 18012 41760
rect 18052 41812 18104 41818
rect 18052 41754 18104 41760
rect 17590 41712 17646 41721
rect 17590 41647 17646 41656
rect 17972 41614 18000 41754
rect 17960 41608 18012 41614
rect 17774 41576 17830 41585
rect 17960 41550 18012 41556
rect 17774 41511 17776 41520
rect 17828 41511 17830 41520
rect 17776 41482 17828 41488
rect 18064 41449 18092 41754
rect 18156 41614 18184 41958
rect 18248 41614 18276 43114
rect 18340 42838 18368 43574
rect 18328 42832 18380 42838
rect 18328 42774 18380 42780
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18340 42362 18368 42502
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 18432 42242 18460 43710
rect 18752 43548 19060 43557
rect 18752 43546 18758 43548
rect 18814 43546 18838 43548
rect 18894 43546 18918 43548
rect 18974 43546 18998 43548
rect 19054 43546 19060 43548
rect 18814 43494 18816 43546
rect 18996 43494 18998 43546
rect 18752 43492 18758 43494
rect 18814 43492 18838 43494
rect 18894 43492 18918 43494
rect 18974 43492 18998 43494
rect 19054 43492 19060 43494
rect 18752 43483 19060 43492
rect 19168 43178 19196 43710
rect 19156 43172 19208 43178
rect 19156 43114 19208 43120
rect 18604 43104 18656 43110
rect 18604 43046 18656 43052
rect 18616 42770 18644 43046
rect 19260 42922 19288 44463
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 19340 43308 19392 43314
rect 19340 43250 19392 43256
rect 19168 42894 19288 42922
rect 18708 42860 19104 42888
rect 18604 42764 18656 42770
rect 18604 42706 18656 42712
rect 18708 42650 18736 42860
rect 19076 42702 19104 42860
rect 18340 42214 18460 42242
rect 18524 42622 18736 42650
rect 18788 42696 18840 42702
rect 18788 42638 18840 42644
rect 19064 42696 19116 42702
rect 19064 42638 19116 42644
rect 18144 41608 18196 41614
rect 18144 41550 18196 41556
rect 18236 41608 18288 41614
rect 18236 41550 18288 41556
rect 18340 41562 18368 42214
rect 18420 42084 18472 42090
rect 18420 42026 18472 42032
rect 18432 41721 18460 42026
rect 18524 41818 18552 42622
rect 18604 42560 18656 42566
rect 18800 42548 18828 42638
rect 18972 42560 19024 42566
rect 18800 42520 18972 42548
rect 18604 42502 18656 42508
rect 18972 42502 19024 42508
rect 18616 42294 18644 42502
rect 18752 42460 19060 42469
rect 18752 42458 18758 42460
rect 18814 42458 18838 42460
rect 18894 42458 18918 42460
rect 18974 42458 18998 42460
rect 19054 42458 19060 42460
rect 18814 42406 18816 42458
rect 18996 42406 18998 42458
rect 18752 42404 18758 42406
rect 18814 42404 18838 42406
rect 18894 42404 18918 42406
rect 18974 42404 18998 42406
rect 19054 42404 19060 42406
rect 18752 42395 19060 42404
rect 19064 42356 19116 42362
rect 19064 42298 19116 42304
rect 18604 42288 18656 42294
rect 19076 42242 19104 42298
rect 18604 42230 18656 42236
rect 18880 42220 18932 42226
rect 18880 42162 18932 42168
rect 18984 42214 19104 42242
rect 18696 42016 18748 42022
rect 18696 41958 18748 41964
rect 18788 42016 18840 42022
rect 18788 41958 18840 41964
rect 18512 41812 18564 41818
rect 18512 41754 18564 41760
rect 18418 41712 18474 41721
rect 18708 41698 18736 41958
rect 18418 41647 18474 41656
rect 18524 41670 18736 41698
rect 18420 41608 18472 41614
rect 18340 41556 18420 41562
rect 18340 41550 18472 41556
rect 18340 41534 18460 41550
rect 18050 41440 18106 41449
rect 18050 41375 18106 41384
rect 17132 38752 17184 38758
rect 18524 38729 18552 41670
rect 18800 41562 18828 41958
rect 18892 41818 18920 42162
rect 18984 42090 19012 42214
rect 18972 42084 19024 42090
rect 18972 42026 19024 42032
rect 18880 41812 18932 41818
rect 18880 41754 18932 41760
rect 18616 41534 18828 41562
rect 17132 38694 17184 38700
rect 18510 38720 18566 38729
rect 18510 38655 18566 38664
rect 18616 37482 18644 41534
rect 18752 41372 19060 41381
rect 18752 41370 18758 41372
rect 18814 41370 18838 41372
rect 18894 41370 18918 41372
rect 18974 41370 18998 41372
rect 19054 41370 19060 41372
rect 18814 41318 18816 41370
rect 18996 41318 18998 41370
rect 18752 41316 18758 41318
rect 18814 41316 18838 41318
rect 18894 41316 18918 41318
rect 18974 41316 18998 41318
rect 19054 41316 19060 41318
rect 18752 41307 19060 41316
rect 19064 40928 19116 40934
rect 19064 40870 19116 40876
rect 19076 40594 19104 40870
rect 19064 40588 19116 40594
rect 19064 40530 19116 40536
rect 19168 40458 19196 42894
rect 19248 42628 19300 42634
rect 19248 42570 19300 42576
rect 19156 40452 19208 40458
rect 19156 40394 19208 40400
rect 18752 40284 19060 40293
rect 18752 40282 18758 40284
rect 18814 40282 18838 40284
rect 18894 40282 18918 40284
rect 18974 40282 18998 40284
rect 19054 40282 19060 40284
rect 18814 40230 18816 40282
rect 18996 40230 18998 40282
rect 18752 40228 18758 40230
rect 18814 40228 18838 40230
rect 18894 40228 18918 40230
rect 18974 40228 18998 40230
rect 19054 40228 19060 40230
rect 18752 40219 19060 40228
rect 18752 39196 19060 39205
rect 18752 39194 18758 39196
rect 18814 39194 18838 39196
rect 18894 39194 18918 39196
rect 18974 39194 18998 39196
rect 19054 39194 19060 39196
rect 18814 39142 18816 39194
rect 18996 39142 18998 39194
rect 18752 39140 18758 39142
rect 18814 39140 18838 39142
rect 18894 39140 18918 39142
rect 18974 39140 18998 39142
rect 19054 39140 19060 39142
rect 18752 39131 19060 39140
rect 19260 38962 19288 42570
rect 19352 42106 19380 43250
rect 19444 42362 19472 43726
rect 19536 43364 19564 44463
rect 19812 43790 19840 44463
rect 19800 43784 19852 43790
rect 19800 43726 19852 43732
rect 19984 43376 20036 43382
rect 19536 43336 19656 43364
rect 19524 43104 19576 43110
rect 19524 43046 19576 43052
rect 19432 42356 19484 42362
rect 19432 42298 19484 42304
rect 19536 42294 19564 43046
rect 19524 42288 19576 42294
rect 19524 42230 19576 42236
rect 19352 42078 19564 42106
rect 19432 42016 19484 42022
rect 19432 41958 19484 41964
rect 19444 41721 19472 41958
rect 19536 41818 19564 42078
rect 19524 41812 19576 41818
rect 19524 41754 19576 41760
rect 19430 41712 19486 41721
rect 19430 41647 19486 41656
rect 19340 41540 19392 41546
rect 19340 41482 19392 41488
rect 19352 41414 19380 41482
rect 19352 41386 19564 41414
rect 19536 40526 19564 41386
rect 19628 41120 19656 43336
rect 19984 43318 20036 43324
rect 19708 43308 19760 43314
rect 19892 43308 19944 43314
rect 19760 43268 19840 43296
rect 19708 43250 19760 43256
rect 19708 43172 19760 43178
rect 19708 43114 19760 43120
rect 19720 41614 19748 43114
rect 19708 41608 19760 41614
rect 19708 41550 19760 41556
rect 19708 41132 19760 41138
rect 19628 41092 19708 41120
rect 19708 41074 19760 41080
rect 19708 40996 19760 41002
rect 19708 40938 19760 40944
rect 19524 40520 19576 40526
rect 19524 40462 19576 40468
rect 19432 40384 19484 40390
rect 19352 40344 19432 40372
rect 19248 38956 19300 38962
rect 19248 38898 19300 38904
rect 18752 38108 19060 38117
rect 18752 38106 18758 38108
rect 18814 38106 18838 38108
rect 18894 38106 18918 38108
rect 18974 38106 18998 38108
rect 19054 38106 19060 38108
rect 18814 38054 18816 38106
rect 18996 38054 18998 38106
rect 18752 38052 18758 38054
rect 18814 38052 18838 38054
rect 18894 38052 18918 38054
rect 18974 38052 18998 38054
rect 19054 38052 19060 38054
rect 18752 38043 19060 38052
rect 18340 37454 18644 37482
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 17236 36922 17264 37198
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 16672 36780 16724 36786
rect 16672 36722 16724 36728
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 17316 36644 17368 36650
rect 17316 36586 17368 36592
rect 16764 35692 16816 35698
rect 16764 35634 16816 35640
rect 16500 35244 16620 35272
rect 16488 35148 16540 35154
rect 16488 35090 16540 35096
rect 16500 34678 16528 35090
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16592 34490 16620 35244
rect 16500 34462 16620 34490
rect 16500 27470 16528 34462
rect 16776 33998 16804 35634
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 16868 34678 16896 34886
rect 16856 34672 16908 34678
rect 16856 34614 16908 34620
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 16764 33992 16816 33998
rect 16764 33934 16816 33940
rect 16580 33516 16632 33522
rect 16580 33458 16632 33464
rect 16592 33114 16620 33458
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16776 32570 16804 33934
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16580 32496 16632 32502
rect 16580 32438 16632 32444
rect 16592 31890 16620 32438
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16592 31754 16620 31826
rect 16592 31726 16712 31754
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16592 29646 16620 31622
rect 16684 30818 16712 31726
rect 16776 30920 16804 31962
rect 16960 31890 16988 33798
rect 17052 33658 17080 34546
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17144 32026 17172 33458
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 16948 31884 17000 31890
rect 16948 31826 17000 31832
rect 16854 31376 16910 31385
rect 16854 31311 16856 31320
rect 16908 31311 16910 31320
rect 16856 31282 16908 31288
rect 16776 30892 16896 30920
rect 16684 30802 16804 30818
rect 16684 30796 16816 30802
rect 16684 30790 16764 30796
rect 16764 30738 16816 30744
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16592 29238 16620 29582
rect 16684 29510 16712 30670
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16580 29232 16632 29238
rect 16580 29174 16632 29180
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16684 28994 16712 29038
rect 16592 28966 16712 28994
rect 16488 27464 16540 27470
rect 16488 27406 16540 27412
rect 16500 25838 16528 27406
rect 16592 27334 16620 28966
rect 16672 28620 16724 28626
rect 16868 28608 16896 30892
rect 16960 29714 16988 31826
rect 17328 31414 17356 36586
rect 17420 36106 17448 36654
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 17408 36100 17460 36106
rect 17408 36042 17460 36048
rect 17592 35624 17644 35630
rect 17592 35566 17644 35572
rect 17408 34672 17460 34678
rect 17408 34614 17460 34620
rect 17420 33930 17448 34614
rect 17500 34604 17552 34610
rect 17500 34546 17552 34552
rect 17512 34202 17540 34546
rect 17604 34202 17632 35566
rect 17972 35086 18000 36518
rect 18052 35148 18104 35154
rect 18052 35090 18104 35096
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17960 34944 18012 34950
rect 17960 34886 18012 34892
rect 17500 34196 17552 34202
rect 17500 34138 17552 34144
rect 17592 34196 17644 34202
rect 17592 34138 17644 34144
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17408 33924 17460 33930
rect 17408 33866 17460 33872
rect 17420 32910 17448 33866
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 17316 31408 17368 31414
rect 17316 31350 17368 31356
rect 17328 29730 17356 31350
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17420 30938 17448 31078
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17512 29850 17540 33934
rect 17604 32978 17632 34138
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17684 33584 17736 33590
rect 17684 33526 17736 33532
rect 17592 32972 17644 32978
rect 17592 32914 17644 32920
rect 17604 30258 17632 32914
rect 17696 30802 17724 33526
rect 17788 33522 17816 33798
rect 17776 33516 17828 33522
rect 17776 33458 17828 33464
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 17592 30048 17644 30054
rect 17592 29990 17644 29996
rect 17604 29850 17632 29990
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17592 29844 17644 29850
rect 17592 29786 17644 29792
rect 16948 29708 17000 29714
rect 17328 29702 17540 29730
rect 16948 29650 17000 29656
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16946 29200 17002 29209
rect 16946 29135 16948 29144
rect 17000 29135 17002 29144
rect 16948 29106 17000 29112
rect 17052 28801 17080 29446
rect 17132 28960 17184 28966
rect 17132 28902 17184 28908
rect 17038 28792 17094 28801
rect 17038 28727 17094 28736
rect 17144 28744 17172 28902
rect 17144 28716 17262 28744
rect 17038 28656 17094 28665
rect 16948 28620 17000 28626
rect 16868 28580 16948 28608
rect 16672 28562 16724 28568
rect 17234 28626 17262 28716
rect 17038 28591 17094 28600
rect 17224 28620 17276 28626
rect 16948 28562 17000 28568
rect 16684 28218 16712 28562
rect 16958 28506 16986 28562
rect 17052 28558 17080 28591
rect 17224 28562 17276 28568
rect 17040 28552 17092 28558
rect 16958 28478 16988 28506
rect 17040 28494 17092 28500
rect 16672 28212 16724 28218
rect 16672 28154 16724 28160
rect 16960 27614 16988 28478
rect 17316 28144 17368 28150
rect 17316 28086 17368 28092
rect 17130 27840 17186 27849
rect 17130 27775 17186 27784
rect 16684 27586 16988 27614
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 16592 25498 16620 26862
rect 16684 25770 16712 27586
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16672 25764 16724 25770
rect 16672 25706 16724 25712
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16488 25424 16540 25430
rect 16488 25366 16540 25372
rect 16500 23474 16528 25366
rect 16776 25362 16804 26930
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16868 26042 16896 26250
rect 16856 26036 16908 26042
rect 16856 25978 16908 25984
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16762 24848 16818 24857
rect 16762 24783 16818 24792
rect 16672 24744 16724 24750
rect 16776 24732 16804 24783
rect 16724 24704 16804 24732
rect 16672 24686 16724 24692
rect 16580 24608 16632 24614
rect 16580 24550 16632 24556
rect 16592 24410 16620 24550
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16776 24274 16804 24704
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 16580 23792 16632 23798
rect 16578 23760 16580 23769
rect 16632 23760 16634 23769
rect 16578 23695 16634 23704
rect 16500 23446 16620 23474
rect 16592 22642 16620 23446
rect 16868 22778 16896 25434
rect 16960 24664 16988 26862
rect 17144 26858 17172 27775
rect 17224 27328 17276 27334
rect 17224 27270 17276 27276
rect 17236 26926 17264 27270
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17132 25968 17184 25974
rect 17132 25910 17184 25916
rect 17144 24886 17172 25910
rect 17328 25514 17356 28086
rect 17408 27328 17460 27334
rect 17408 27270 17460 27276
rect 17420 25702 17448 27270
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 17328 25486 17448 25514
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17328 24954 17356 25298
rect 17316 24948 17368 24954
rect 17316 24890 17368 24896
rect 17132 24880 17184 24886
rect 17132 24822 17184 24828
rect 17420 24818 17448 25486
rect 17512 24857 17540 29702
rect 17592 29232 17644 29238
rect 17592 29174 17644 29180
rect 17604 25294 17632 29174
rect 17696 28082 17724 30738
rect 17788 28150 17816 32846
rect 17972 31754 18000 34886
rect 18064 31890 18092 35090
rect 18156 34950 18184 37062
rect 18236 36644 18288 36650
rect 18236 36586 18288 36592
rect 18248 35834 18276 36586
rect 18236 35828 18288 35834
rect 18236 35770 18288 35776
rect 18144 34944 18196 34950
rect 18144 34886 18196 34892
rect 18248 34762 18276 35770
rect 18156 34734 18276 34762
rect 18156 33402 18184 34734
rect 18236 33856 18288 33862
rect 18236 33798 18288 33804
rect 18248 33522 18276 33798
rect 18236 33516 18288 33522
rect 18236 33458 18288 33464
rect 18156 33374 18276 33402
rect 18142 32328 18198 32337
rect 18142 32263 18198 32272
rect 18052 31884 18104 31890
rect 18052 31826 18104 31832
rect 17972 31726 18092 31754
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17972 30938 18000 31282
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 29510 17908 30194
rect 17868 29504 17920 29510
rect 17868 29446 17920 29452
rect 17880 29170 17908 29446
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17868 28960 17920 28966
rect 17868 28902 17920 28908
rect 17880 28393 17908 28902
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17866 28384 17922 28393
rect 17866 28319 17922 28328
rect 17776 28144 17828 28150
rect 17776 28086 17828 28092
rect 17972 28082 18000 28494
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17696 26450 17724 28018
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 26994 17908 27270
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17776 26920 17828 26926
rect 17776 26862 17828 26868
rect 17684 26444 17736 26450
rect 17684 26386 17736 26392
rect 17592 25288 17644 25294
rect 17592 25230 17644 25236
rect 17498 24848 17554 24857
rect 17408 24812 17460 24818
rect 17236 24772 17408 24800
rect 16960 24636 17080 24664
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16592 21593 16620 21966
rect 16578 21584 16634 21593
rect 16578 21519 16634 21528
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16500 21010 16528 21422
rect 16488 21004 16540 21010
rect 16488 20946 16540 20952
rect 16684 20874 16712 22374
rect 16868 22094 16896 22578
rect 16868 22066 16988 22094
rect 16960 21729 16988 22066
rect 16762 21720 16818 21729
rect 16762 21655 16818 21664
rect 16946 21720 17002 21729
rect 16946 21655 17002 21664
rect 16776 21622 16804 21655
rect 16764 21616 16816 21622
rect 16764 21558 16816 21564
rect 17052 21486 17080 24636
rect 17236 22438 17264 24772
rect 17498 24783 17500 24792
rect 17408 24754 17460 24760
rect 17552 24783 17554 24792
rect 17500 24754 17552 24760
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17408 24064 17460 24070
rect 17408 24006 17460 24012
rect 17316 22500 17368 22506
rect 17316 22442 17368 22448
rect 17224 22432 17276 22438
rect 17224 22374 17276 22380
rect 17328 22166 17356 22442
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 17224 21956 17276 21962
rect 17224 21898 17276 21904
rect 17236 21593 17264 21898
rect 17222 21584 17278 21593
rect 17222 21519 17278 21528
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 17040 21480 17092 21486
rect 17328 21434 17356 22102
rect 17040 21422 17092 21428
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16580 20800 16632 20806
rect 16580 20742 16632 20748
rect 16592 20058 16620 20742
rect 16672 20256 16724 20262
rect 16672 20198 16724 20204
rect 16580 20052 16632 20058
rect 16408 20012 16528 20040
rect 16304 19994 16356 20000
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16316 18970 16344 19858
rect 16408 19378 16436 19858
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16224 18698 16344 18714
rect 16224 18692 16356 18698
rect 16224 18686 16304 18692
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15488 16561 15516 17546
rect 15580 16658 15608 18686
rect 16304 18634 16356 18640
rect 15936 18624 15988 18630
rect 15672 18584 15936 18612
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15474 16552 15530 16561
rect 15474 16487 15530 16496
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15198 15600 15254 15609
rect 15198 15535 15254 15544
rect 15212 14006 15240 15535
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 15304 14074 15332 15302
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15028 12406 15148 12434
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14922 11112 14978 11121
rect 14922 11047 14924 11056
rect 14976 11047 14978 11056
rect 14924 11018 14976 11024
rect 14924 10668 14976 10674
rect 14924 10610 14976 10616
rect 14936 8566 14964 10610
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14936 7478 14964 8502
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14924 5636 14976 5642
rect 14924 5578 14976 5584
rect 14936 5166 14964 5578
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14936 2106 14964 2246
rect 14740 2100 14792 2106
rect 14740 2042 14792 2048
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 15028 1902 15056 12406
rect 15212 11762 15240 13262
rect 15396 12102 15424 16390
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15200 11756 15252 11762
rect 15252 11716 15332 11744
rect 15200 11698 15252 11704
rect 15108 11280 15160 11286
rect 15108 11222 15160 11228
rect 15120 10985 15148 11222
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15106 10976 15162 10985
rect 15106 10911 15162 10920
rect 15212 10606 15240 11086
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 8566 15148 8774
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15212 2774 15240 9658
rect 15304 6322 15332 11716
rect 15396 10674 15424 12038
rect 15474 10840 15530 10849
rect 15474 10775 15530 10784
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15488 9674 15516 10775
rect 15396 9646 15516 9674
rect 15396 8022 15424 9646
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 9042 15516 9318
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15396 6866 15424 7822
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15396 5710 15424 6802
rect 15488 5846 15516 8774
rect 15580 8430 15608 16594
rect 15568 8424 15620 8430
rect 15568 8366 15620 8372
rect 15580 7954 15608 8366
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15580 5846 15608 6394
rect 15672 5896 15700 18584
rect 15936 18566 15988 18572
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 15785 17980 16093 17989
rect 15785 17978 15791 17980
rect 15847 17978 15871 17980
rect 15927 17978 15951 17980
rect 16007 17978 16031 17980
rect 16087 17978 16093 17980
rect 15847 17926 15849 17978
rect 16029 17926 16031 17978
rect 15785 17924 15791 17926
rect 15847 17924 15871 17926
rect 15927 17924 15951 17926
rect 16007 17924 16031 17926
rect 16087 17924 16093 17926
rect 15785 17915 16093 17924
rect 15785 16892 16093 16901
rect 15785 16890 15791 16892
rect 15847 16890 15871 16892
rect 15927 16890 15951 16892
rect 16007 16890 16031 16892
rect 16087 16890 16093 16892
rect 15847 16838 15849 16890
rect 16029 16838 16031 16890
rect 15785 16836 15791 16838
rect 15847 16836 15871 16838
rect 15927 16836 15951 16838
rect 16007 16836 16031 16838
rect 16087 16836 16093 16838
rect 15785 16827 16093 16836
rect 16132 16794 16160 18022
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16316 16674 16344 18634
rect 16500 17320 16528 20012
rect 16580 19994 16632 20000
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16592 19446 16620 19654
rect 16580 19440 16632 19446
rect 16580 19382 16632 19388
rect 15936 16652 15988 16658
rect 15856 16612 15936 16640
rect 15856 16017 15884 16612
rect 15936 16594 15988 16600
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 16224 16646 16344 16674
rect 16408 17292 16528 17320
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15948 16250 15976 16458
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16040 16182 16068 16594
rect 16028 16176 16080 16182
rect 16028 16118 16080 16124
rect 15842 16008 15898 16017
rect 15842 15943 15898 15952
rect 15785 15804 16093 15813
rect 15785 15802 15791 15804
rect 15847 15802 15871 15804
rect 15927 15802 15951 15804
rect 16007 15802 16031 15804
rect 16087 15802 16093 15804
rect 15847 15750 15849 15802
rect 16029 15750 16031 15802
rect 15785 15748 15791 15750
rect 15847 15748 15871 15750
rect 15927 15748 15951 15750
rect 16007 15748 16031 15750
rect 16087 15748 16093 15750
rect 15785 15739 16093 15748
rect 16224 15201 16252 16646
rect 16304 16176 16356 16182
rect 16304 16118 16356 16124
rect 16210 15192 16266 15201
rect 16210 15127 16266 15136
rect 15785 14716 16093 14725
rect 15785 14714 15791 14716
rect 15847 14714 15871 14716
rect 15927 14714 15951 14716
rect 16007 14714 16031 14716
rect 16087 14714 16093 14716
rect 15847 14662 15849 14714
rect 16029 14662 16031 14714
rect 15785 14660 15791 14662
rect 15847 14660 15871 14662
rect 15927 14660 15951 14662
rect 16007 14660 16031 14662
rect 16087 14660 16093 14662
rect 15785 14651 16093 14660
rect 16120 14476 16172 14482
rect 16172 14436 16252 14464
rect 16120 14418 16172 14424
rect 16118 14376 16174 14385
rect 16118 14311 16120 14320
rect 16172 14311 16174 14320
rect 16120 14282 16172 14288
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15785 13628 16093 13637
rect 15785 13626 15791 13628
rect 15847 13626 15871 13628
rect 15927 13626 15951 13628
rect 16007 13626 16031 13628
rect 16087 13626 16093 13628
rect 15847 13574 15849 13626
rect 16029 13574 16031 13626
rect 15785 13572 15791 13574
rect 15847 13572 15871 13574
rect 15927 13572 15951 13574
rect 16007 13572 16031 13574
rect 16087 13572 16093 13574
rect 15785 13563 16093 13572
rect 15785 12540 16093 12549
rect 15785 12538 15791 12540
rect 15847 12538 15871 12540
rect 15927 12538 15951 12540
rect 16007 12538 16031 12540
rect 16087 12538 16093 12540
rect 15847 12486 15849 12538
rect 16029 12486 16031 12538
rect 15785 12484 15791 12486
rect 15847 12484 15871 12486
rect 15927 12484 15951 12486
rect 16007 12484 16031 12486
rect 16087 12484 16093 12486
rect 15785 12475 16093 12484
rect 15785 11452 16093 11461
rect 15785 11450 15791 11452
rect 15847 11450 15871 11452
rect 15927 11450 15951 11452
rect 16007 11450 16031 11452
rect 16087 11450 16093 11452
rect 15847 11398 15849 11450
rect 16029 11398 16031 11450
rect 15785 11396 15791 11398
rect 15847 11396 15871 11398
rect 15927 11396 15951 11398
rect 16007 11396 16031 11398
rect 16087 11396 16093 11398
rect 15785 11387 16093 11396
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15764 10742 15792 11222
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15856 10674 15884 11222
rect 16132 11218 16160 13874
rect 16224 11218 16252 14436
rect 16316 14414 16344 16118
rect 16408 15162 16436 17292
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16316 12374 16344 14350
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16408 12220 16436 14350
rect 16500 13938 16528 17070
rect 16592 16436 16620 17138
rect 16684 16590 16712 20198
rect 16776 16658 16804 21422
rect 17236 21418 17356 21434
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17224 21412 17356 21418
rect 17276 21406 17356 21412
rect 17224 21354 17276 21360
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16868 19514 16896 19790
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16854 17912 16910 17921
rect 16854 17847 16910 17856
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16592 16408 16712 16436
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 13932 16540 13938
rect 16488 13874 16540 13880
rect 16500 13394 16528 13874
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16592 13274 16620 14554
rect 16684 13410 16712 16408
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16776 14074 16804 15642
rect 16868 15502 16896 17847
rect 16856 15496 16908 15502
rect 16856 15438 16908 15444
rect 16960 14618 16988 20266
rect 17040 19916 17092 19922
rect 17040 19858 17092 19864
rect 17052 18873 17080 19858
rect 17144 19334 17172 21354
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17328 19446 17356 19654
rect 17316 19440 17368 19446
rect 17316 19382 17368 19388
rect 17144 19306 17356 19334
rect 17130 19000 17186 19009
rect 17186 18958 17264 18986
rect 17130 18935 17186 18944
rect 17038 18864 17094 18873
rect 17038 18799 17094 18808
rect 17052 17320 17080 18799
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17144 17678 17172 18702
rect 17236 18290 17264 18958
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17052 17292 17172 17320
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16868 13530 16896 14418
rect 16946 13832 17002 13841
rect 16946 13767 17002 13776
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16960 13462 16988 13767
rect 16948 13456 17000 13462
rect 16684 13382 16896 13410
rect 16948 13398 17000 13404
rect 16592 13246 16712 13274
rect 16488 12232 16540 12238
rect 16408 12192 16488 12220
rect 16488 12174 16540 12180
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15785 10364 16093 10373
rect 15785 10362 15791 10364
rect 15847 10362 15871 10364
rect 15927 10362 15951 10364
rect 16007 10362 16031 10364
rect 16087 10362 16093 10364
rect 15847 10310 15849 10362
rect 16029 10310 16031 10362
rect 15785 10308 15791 10310
rect 15847 10308 15871 10310
rect 15927 10308 15951 10310
rect 16007 10308 16031 10310
rect 16087 10308 16093 10310
rect 15785 10299 16093 10308
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15764 9722 15792 9930
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 16132 9636 16160 11154
rect 16224 10810 16252 11154
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16316 10674 16344 11494
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16408 10606 16436 12038
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16500 10713 16528 11698
rect 16592 11665 16620 12038
rect 16578 11656 16634 11665
rect 16578 11591 16634 11600
rect 16486 10704 16542 10713
rect 16486 10639 16542 10648
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16210 9752 16266 9761
rect 16266 9710 16344 9738
rect 16210 9687 16266 9696
rect 16132 9608 16252 9636
rect 15785 9276 16093 9285
rect 15785 9274 15791 9276
rect 15847 9274 15871 9276
rect 15927 9274 15951 9276
rect 16007 9274 16031 9276
rect 16087 9274 16093 9276
rect 15847 9222 15849 9274
rect 16029 9222 16031 9274
rect 15785 9220 15791 9222
rect 15847 9220 15871 9222
rect 15927 9220 15951 9222
rect 16007 9220 16031 9222
rect 16087 9220 16093 9222
rect 15785 9211 16093 9220
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 15785 8188 16093 8197
rect 15785 8186 15791 8188
rect 15847 8186 15871 8188
rect 15927 8186 15951 8188
rect 16007 8186 16031 8188
rect 16087 8186 16093 8188
rect 15847 8134 15849 8186
rect 16029 8134 16031 8186
rect 15785 8132 15791 8134
rect 15847 8132 15871 8134
rect 15927 8132 15951 8134
rect 16007 8132 16031 8134
rect 16087 8132 16093 8134
rect 15785 8123 16093 8132
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15856 7478 15884 7958
rect 15844 7472 15896 7478
rect 15844 7414 15896 7420
rect 15785 7100 16093 7109
rect 15785 7098 15791 7100
rect 15847 7098 15871 7100
rect 15927 7098 15951 7100
rect 16007 7098 16031 7100
rect 16087 7098 16093 7100
rect 15847 7046 15849 7098
rect 16029 7046 16031 7098
rect 15785 7044 15791 7046
rect 15847 7044 15871 7046
rect 15927 7044 15951 7046
rect 16007 7044 16031 7046
rect 16087 7044 16093 7046
rect 15785 7035 16093 7044
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 15672 5868 15792 5896
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 5166 15424 5646
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15304 4282 15332 5034
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15488 4214 15516 5782
rect 15764 5522 15792 5868
rect 15672 5494 15792 5522
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15580 5001 15608 5102
rect 15566 4992 15622 5001
rect 15566 4927 15622 4936
rect 15568 4616 15620 4622
rect 15566 4584 15568 4593
rect 15620 4584 15622 4593
rect 15566 4519 15622 4528
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15212 2746 15424 2774
rect 15396 1970 15424 2746
rect 15566 2544 15622 2553
rect 15566 2479 15622 2488
rect 15580 2446 15608 2479
rect 15672 2446 15700 5494
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15764 5030 15792 5102
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 16132 4622 16160 8774
rect 16224 7993 16252 9608
rect 16316 9042 16344 9710
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16210 7984 16266 7993
rect 16210 7919 16266 7928
rect 16224 7886 16252 7919
rect 16212 7880 16264 7886
rect 16264 7840 16344 7868
rect 16212 7822 16264 7828
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5914 16252 6054
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16316 5778 16344 7840
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16224 5137 16252 5646
rect 16210 5128 16266 5137
rect 16316 5098 16344 5714
rect 16408 5681 16436 10542
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8090 16528 8774
rect 16684 8634 16712 13246
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16776 10996 16804 12174
rect 16868 11762 16896 13382
rect 17052 12918 17080 17138
rect 17144 14414 17172 17292
rect 17236 16250 17264 18226
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17224 16040 17276 16046
rect 17224 15982 17276 15988
rect 17236 15094 17264 15982
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17328 14600 17356 19306
rect 17236 14572 17356 14600
rect 17236 14482 17264 14572
rect 17420 14498 17448 24006
rect 17512 21962 17540 24074
rect 17500 21956 17552 21962
rect 17500 21898 17552 21904
rect 17498 21720 17554 21729
rect 17604 21706 17632 25230
rect 17696 23730 17724 26386
rect 17788 24614 17816 26862
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17868 25288 17920 25294
rect 17868 25230 17920 25236
rect 17880 24682 17908 25230
rect 17972 24886 18000 25842
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17868 24676 17920 24682
rect 17868 24618 17920 24624
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17788 22642 17816 24550
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17776 21888 17828 21894
rect 17776 21830 17828 21836
rect 17604 21678 17724 21706
rect 17498 21655 17554 21664
rect 17512 18290 17540 21655
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17604 21350 17632 21490
rect 17696 21486 17724 21678
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17696 20330 17724 21422
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17788 19990 17816 21830
rect 17880 21554 17908 22510
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17880 21146 17908 21490
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17866 20496 17922 20505
rect 17972 20482 18000 24822
rect 18064 23050 18092 31726
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 20602 18092 21422
rect 18052 20596 18104 20602
rect 18052 20538 18104 20544
rect 17922 20466 18000 20482
rect 17922 20460 18012 20466
rect 17922 20454 17960 20460
rect 17866 20431 17922 20440
rect 17960 20402 18012 20408
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17500 18284 17552 18290
rect 17500 18226 17552 18232
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17882 17908 18090
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17512 15065 17540 17614
rect 17866 17096 17922 17105
rect 17866 17031 17922 17040
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17696 16794 17724 16934
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17880 16590 17908 17031
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17972 16182 18000 19654
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17814 18092 18158
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 18156 17252 18184 32263
rect 18248 30326 18276 33374
rect 18236 30320 18288 30326
rect 18236 30262 18288 30268
rect 18234 30152 18290 30161
rect 18234 30087 18290 30096
rect 18248 25809 18276 30087
rect 18234 25800 18290 25809
rect 18234 25735 18290 25744
rect 18340 22094 18368 37454
rect 18512 37324 18564 37330
rect 18512 37266 18564 37272
rect 18420 35760 18472 35766
rect 18420 35702 18472 35708
rect 18432 32026 18460 35702
rect 18420 32020 18472 32026
rect 18420 31962 18472 31968
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18432 30433 18460 31826
rect 18418 30424 18474 30433
rect 18418 30359 18474 30368
rect 18420 30320 18472 30326
rect 18420 30262 18472 30268
rect 18432 23848 18460 30262
rect 18524 24154 18552 37266
rect 18752 37020 19060 37029
rect 18752 37018 18758 37020
rect 18814 37018 18838 37020
rect 18894 37018 18918 37020
rect 18974 37018 18998 37020
rect 19054 37018 19060 37020
rect 18814 36966 18816 37018
rect 18996 36966 18998 37018
rect 18752 36964 18758 36966
rect 18814 36964 18838 36966
rect 18894 36964 18918 36966
rect 18974 36964 18998 36966
rect 19054 36964 19060 36966
rect 18752 36955 19060 36964
rect 19260 36174 19288 38898
rect 19352 37330 19380 40344
rect 19432 40326 19484 40332
rect 19616 40384 19668 40390
rect 19616 40326 19668 40332
rect 19628 40186 19656 40326
rect 19720 40225 19748 40938
rect 19812 40730 19840 43268
rect 19892 43250 19944 43256
rect 19904 42090 19932 43250
rect 19892 42084 19944 42090
rect 19892 42026 19944 42032
rect 19892 41132 19944 41138
rect 19892 41074 19944 41080
rect 19800 40724 19852 40730
rect 19800 40666 19852 40672
rect 19800 40384 19852 40390
rect 19800 40326 19852 40332
rect 19706 40216 19762 40225
rect 19616 40180 19668 40186
rect 19812 40186 19840 40326
rect 19706 40151 19762 40160
rect 19800 40180 19852 40186
rect 19616 40122 19668 40128
rect 19800 40122 19852 40128
rect 19432 39908 19484 39914
rect 19432 39850 19484 39856
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19352 36650 19380 36790
rect 19340 36644 19392 36650
rect 19340 36586 19392 36592
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 18752 35932 19060 35941
rect 18752 35930 18758 35932
rect 18814 35930 18838 35932
rect 18894 35930 18918 35932
rect 18974 35930 18998 35932
rect 19054 35930 19060 35932
rect 18814 35878 18816 35930
rect 18996 35878 18998 35930
rect 18752 35876 18758 35878
rect 18814 35876 18838 35878
rect 18894 35876 18918 35878
rect 18974 35876 18998 35878
rect 19054 35876 19060 35878
rect 18752 35867 19060 35876
rect 19064 35624 19116 35630
rect 18878 35592 18934 35601
rect 19064 35566 19116 35572
rect 18878 35527 18880 35536
rect 18932 35527 18934 35536
rect 18880 35498 18932 35504
rect 19076 35290 19104 35566
rect 19064 35284 19116 35290
rect 19064 35226 19116 35232
rect 19156 35012 19208 35018
rect 19156 34954 19208 34960
rect 18752 34844 19060 34853
rect 18752 34842 18758 34844
rect 18814 34842 18838 34844
rect 18894 34842 18918 34844
rect 18974 34842 18998 34844
rect 19054 34842 19060 34844
rect 18814 34790 18816 34842
rect 18996 34790 18998 34842
rect 18752 34788 18758 34790
rect 18814 34788 18838 34790
rect 18894 34788 18918 34790
rect 18974 34788 18998 34790
rect 19054 34788 19060 34790
rect 18752 34779 19060 34788
rect 19168 34746 19196 34954
rect 19156 34740 19208 34746
rect 19156 34682 19208 34688
rect 19260 34626 19288 36110
rect 19340 36032 19392 36038
rect 19340 35974 19392 35980
rect 19352 35834 19380 35974
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19168 34610 19288 34626
rect 19352 34610 19380 35022
rect 19156 34604 19288 34610
rect 19208 34598 19288 34604
rect 19340 34604 19392 34610
rect 19156 34546 19208 34552
rect 19340 34546 19392 34552
rect 18752 33756 19060 33765
rect 18752 33754 18758 33756
rect 18814 33754 18838 33756
rect 18894 33754 18918 33756
rect 18974 33754 18998 33756
rect 19054 33754 19060 33756
rect 18814 33702 18816 33754
rect 18996 33702 18998 33754
rect 18752 33700 18758 33702
rect 18814 33700 18838 33702
rect 18894 33700 18918 33702
rect 18974 33700 18998 33702
rect 19054 33700 19060 33702
rect 18752 33691 19060 33700
rect 18880 33652 18932 33658
rect 19064 33652 19116 33658
rect 18932 33612 19064 33640
rect 18880 33594 18932 33600
rect 19064 33594 19116 33600
rect 19168 33590 19196 34546
rect 19156 33584 19208 33590
rect 18878 33552 18934 33561
rect 18604 33516 18656 33522
rect 19156 33526 19208 33532
rect 18878 33487 18934 33496
rect 18604 33458 18656 33464
rect 18616 33114 18644 33458
rect 18892 33318 18920 33487
rect 19168 33402 19196 33526
rect 19168 33374 19288 33402
rect 18880 33312 18932 33318
rect 18880 33254 18932 33260
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 18752 32668 19060 32677
rect 18752 32666 18758 32668
rect 18814 32666 18838 32668
rect 18894 32666 18918 32668
rect 18974 32666 18998 32668
rect 19054 32666 19060 32668
rect 18814 32614 18816 32666
rect 18996 32614 18998 32666
rect 18752 32612 18758 32614
rect 18814 32612 18838 32614
rect 18894 32612 18918 32614
rect 18974 32612 18998 32614
rect 19054 32612 19060 32614
rect 18752 32603 19060 32612
rect 19260 32434 19288 33374
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19156 32224 19208 32230
rect 19156 32166 19208 32172
rect 18752 31580 19060 31589
rect 18752 31578 18758 31580
rect 18814 31578 18838 31580
rect 18894 31578 18918 31580
rect 18974 31578 18998 31580
rect 19054 31578 19060 31580
rect 18814 31526 18816 31578
rect 18996 31526 18998 31578
rect 18752 31524 18758 31526
rect 18814 31524 18838 31526
rect 18894 31524 18918 31526
rect 18974 31524 18998 31526
rect 19054 31524 19060 31526
rect 18752 31515 19060 31524
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18616 30938 18644 31078
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18616 30258 18644 30534
rect 18752 30492 19060 30501
rect 18752 30490 18758 30492
rect 18814 30490 18838 30492
rect 18894 30490 18918 30492
rect 18974 30490 18998 30492
rect 19054 30490 19060 30492
rect 18814 30438 18816 30490
rect 18996 30438 18998 30490
rect 18752 30436 18758 30438
rect 18814 30436 18838 30438
rect 18894 30436 18918 30438
rect 18974 30436 18998 30438
rect 19054 30436 19060 30438
rect 18752 30427 19060 30436
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18752 29404 19060 29413
rect 18752 29402 18758 29404
rect 18814 29402 18838 29404
rect 18894 29402 18918 29404
rect 18974 29402 18998 29404
rect 19054 29402 19060 29404
rect 18814 29350 18816 29402
rect 18996 29350 18998 29402
rect 18752 29348 18758 29350
rect 18814 29348 18838 29350
rect 18894 29348 18918 29350
rect 18974 29348 18998 29350
rect 19054 29348 19060 29350
rect 18752 29339 19060 29348
rect 19168 29238 19196 32166
rect 19444 31754 19472 39850
rect 19708 36644 19760 36650
rect 19708 36586 19760 36592
rect 19524 34944 19576 34950
rect 19524 34886 19576 34892
rect 19536 34678 19564 34886
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19524 32496 19576 32502
rect 19522 32464 19524 32473
rect 19576 32464 19578 32473
rect 19522 32399 19578 32408
rect 19536 31754 19564 32399
rect 19352 31726 19472 31754
rect 19524 31748 19576 31754
rect 19248 30592 19300 30598
rect 19248 30534 19300 30540
rect 19260 30122 19288 30534
rect 19352 30326 19380 31726
rect 19524 31690 19576 31696
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19432 30184 19484 30190
rect 19432 30126 19484 30132
rect 19248 30116 19300 30122
rect 19248 30058 19300 30064
rect 19248 29572 19300 29578
rect 19248 29514 19300 29520
rect 19156 29232 19208 29238
rect 19156 29174 19208 29180
rect 18696 28552 18748 28558
rect 18616 28500 18696 28506
rect 18616 28494 18748 28500
rect 18616 28478 18736 28494
rect 18616 28082 18644 28478
rect 18752 28316 19060 28325
rect 18752 28314 18758 28316
rect 18814 28314 18838 28316
rect 18894 28314 18918 28316
rect 18974 28314 18998 28316
rect 19054 28314 19060 28316
rect 18814 28262 18816 28314
rect 18996 28262 18998 28314
rect 18752 28260 18758 28262
rect 18814 28260 18838 28262
rect 18894 28260 18918 28262
rect 18974 28260 18998 28262
rect 19054 28260 19060 28262
rect 18752 28251 19060 28260
rect 19260 28098 19288 29514
rect 19444 28948 19472 30126
rect 19524 29232 19576 29238
rect 19524 29174 19576 29180
rect 19352 28920 19472 28948
rect 19352 28150 19380 28920
rect 19430 28792 19486 28801
rect 19536 28762 19564 29174
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19430 28727 19486 28736
rect 19524 28756 19576 28762
rect 19444 28694 19472 28727
rect 19524 28698 19576 28704
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19628 28558 19656 28902
rect 19616 28552 19668 28558
rect 19616 28494 19668 28500
rect 19616 28212 19668 28218
rect 19616 28154 19668 28160
rect 18604 28076 18656 28082
rect 18604 28018 18656 28024
rect 19168 28070 19288 28098
rect 19340 28144 19392 28150
rect 19432 28144 19484 28150
rect 19340 28086 19392 28092
rect 19430 28112 19432 28121
rect 19484 28112 19486 28121
rect 18752 27228 19060 27237
rect 18752 27226 18758 27228
rect 18814 27226 18838 27228
rect 18894 27226 18918 27228
rect 18974 27226 18998 27228
rect 19054 27226 19060 27228
rect 18814 27174 18816 27226
rect 18996 27174 18998 27226
rect 18752 27172 18758 27174
rect 18814 27172 18838 27174
rect 18894 27172 18918 27174
rect 18974 27172 18998 27174
rect 19054 27172 19060 27174
rect 18752 27163 19060 27172
rect 18752 26140 19060 26149
rect 18752 26138 18758 26140
rect 18814 26138 18838 26140
rect 18894 26138 18918 26140
rect 18974 26138 18998 26140
rect 19054 26138 19060 26140
rect 18814 26086 18816 26138
rect 18996 26086 18998 26138
rect 18752 26084 18758 26086
rect 18814 26084 18838 26086
rect 18894 26084 18918 26086
rect 18974 26084 18998 26086
rect 19054 26084 19060 26086
rect 18752 26075 19060 26084
rect 19168 25226 19196 28070
rect 19352 27996 19380 28086
rect 19430 28047 19486 28056
rect 19432 28008 19484 28014
rect 19352 27968 19432 27996
rect 19352 27334 19380 27968
rect 19432 27950 19484 27956
rect 19628 27878 19656 28154
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19628 27470 19656 27814
rect 19616 27464 19668 27470
rect 19616 27406 19668 27412
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 25294 19288 26182
rect 19248 25288 19300 25294
rect 19248 25230 19300 25236
rect 19156 25220 19208 25226
rect 19156 25162 19208 25168
rect 18752 25052 19060 25061
rect 18752 25050 18758 25052
rect 18814 25050 18838 25052
rect 18894 25050 18918 25052
rect 18974 25050 18998 25052
rect 19054 25050 19060 25052
rect 18814 24998 18816 25050
rect 18996 24998 18998 25050
rect 18752 24996 18758 24998
rect 18814 24996 18838 24998
rect 18894 24996 18918 24998
rect 18974 24996 18998 24998
rect 19054 24996 19060 24998
rect 18752 24987 19060 24996
rect 19248 24200 19300 24206
rect 18524 24126 18644 24154
rect 19248 24142 19300 24148
rect 18432 23820 18552 23848
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18432 23118 18460 23666
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18524 22964 18552 23820
rect 18064 17224 18184 17252
rect 18248 22066 18368 22094
rect 18432 22936 18552 22964
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17498 15056 17554 15065
rect 17498 14991 17554 15000
rect 17224 14476 17276 14482
rect 17224 14418 17276 14424
rect 17328 14470 17448 14498
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17328 14278 17356 14470
rect 17408 14408 17460 14414
rect 17408 14350 17460 14356
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17420 14074 17448 14350
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17040 12912 17092 12918
rect 16960 12872 17040 12900
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16856 11008 16908 11014
rect 16776 10968 16856 10996
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16684 7546 16712 8570
rect 16776 8072 16804 10968
rect 16856 10950 16908 10956
rect 16960 9586 16988 12872
rect 17040 12854 17092 12860
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11762 17080 12242
rect 17144 11830 17172 12582
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17144 11150 17172 11766
rect 17222 11384 17278 11393
rect 17222 11319 17278 11328
rect 17132 11144 17184 11150
rect 17038 11112 17094 11121
rect 17132 11086 17184 11092
rect 17038 11047 17040 11056
rect 17092 11047 17094 11056
rect 17040 11018 17092 11024
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17144 9382 17172 11086
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 16856 9036 16908 9042
rect 16908 8996 17080 9024
rect 16856 8978 16908 8984
rect 17052 8922 17080 8996
rect 17144 8922 17172 9318
rect 17052 8894 17172 8922
rect 16856 8084 16908 8090
rect 16776 8044 16856 8072
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16776 6458 16804 8044
rect 16856 8026 16908 8032
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16394 5672 16450 5681
rect 16394 5607 16450 5616
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 16210 5063 16266 5072
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 16408 4826 16436 5102
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16592 4729 16620 5510
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 16578 4720 16634 4729
rect 16578 4655 16634 4664
rect 16684 4622 16712 5170
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15660 2440 15712 2446
rect 16396 2440 16448 2446
rect 15660 2382 15712 2388
rect 16394 2408 16396 2417
rect 16448 2408 16450 2417
rect 16394 2343 16450 2352
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 15488 2106 15516 2246
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15016 1896 15068 1902
rect 15016 1838 15068 1844
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 14740 1760 14792 1766
rect 14568 1720 14740 1748
rect 14464 1284 14516 1290
rect 14464 1226 14516 1232
rect 14568 160 14596 1720
rect 14740 1702 14792 1708
rect 15108 1556 15160 1562
rect 14844 1516 15108 1544
rect 14844 160 14872 1516
rect 15108 1498 15160 1504
rect 15200 1488 15252 1494
rect 15120 1436 15200 1442
rect 15120 1430 15252 1436
rect 15120 1414 15240 1430
rect 15120 160 15148 1414
rect 15396 160 15424 1770
rect 15752 1760 15804 1766
rect 15672 1720 15752 1748
rect 15672 160 15700 1720
rect 15752 1702 15804 1708
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16120 1488 16172 1494
rect 15948 1448 16120 1476
rect 15948 160 15976 1448
rect 16120 1430 16172 1436
rect 16224 1290 16252 2246
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16316 1562 16344 1838
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16500 1442 16528 2246
rect 16776 2038 16804 3062
rect 16960 2446 16988 7414
rect 17052 2825 17080 8894
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17144 7954 17172 8774
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17132 5772 17184 5778
rect 17132 5714 17184 5720
rect 17144 5370 17172 5714
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17236 4162 17264 11319
rect 17328 9654 17356 12174
rect 17420 11150 17448 13874
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17604 9674 17632 15098
rect 17880 15094 17908 15982
rect 17972 15502 18000 16118
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 17776 15088 17828 15094
rect 17776 15030 17828 15036
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17788 14906 17816 15030
rect 17788 14878 17908 14906
rect 17774 14512 17830 14521
rect 17774 14447 17776 14456
rect 17828 14447 17830 14456
rect 17776 14418 17828 14424
rect 17880 14278 17908 14878
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17788 13326 17816 14010
rect 17972 13870 18000 15302
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17972 12850 18000 13806
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17788 12306 17816 12582
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17972 11914 18000 12786
rect 17880 11886 18000 11914
rect 17880 11762 17908 11886
rect 17868 11756 17920 11762
rect 17868 11698 17920 11704
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17776 11144 17828 11150
rect 17880 11132 17908 11698
rect 17972 11257 18000 11698
rect 17958 11248 18014 11257
rect 17958 11183 18014 11192
rect 17880 11104 18000 11132
rect 17776 11086 17828 11092
rect 17316 9648 17368 9654
rect 17316 9590 17368 9596
rect 17420 9646 17632 9674
rect 17328 8566 17356 9590
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17420 7886 17448 9646
rect 17788 9489 17816 11086
rect 17774 9480 17830 9489
rect 17774 9415 17830 9424
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17328 7478 17356 7754
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17512 5817 17540 9318
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 7750 17632 8910
rect 17684 8424 17736 8430
rect 17684 8366 17736 8372
rect 17696 7750 17724 8366
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17498 5808 17554 5817
rect 17498 5743 17554 5752
rect 17512 5710 17540 5743
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17604 5234 17632 7686
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17696 5642 17724 6598
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17604 4729 17632 5170
rect 17590 4720 17646 4729
rect 17590 4655 17646 4664
rect 17696 4282 17724 5170
rect 17788 5166 17816 9415
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 6866 17908 8434
rect 17972 8106 18000 11104
rect 18064 8242 18092 17224
rect 18144 14000 18196 14006
rect 18144 13942 18196 13948
rect 18156 9654 18184 13942
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18156 8838 18184 9386
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18156 8401 18184 8502
rect 18142 8392 18198 8401
rect 18142 8327 18198 8336
rect 18064 8214 18184 8242
rect 17972 8078 18092 8106
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17972 7002 18000 7958
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6458 17908 6802
rect 17958 6760 18014 6769
rect 17958 6695 18014 6704
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17972 6225 18000 6695
rect 18064 6662 18092 8078
rect 18156 6769 18184 8214
rect 18142 6760 18198 6769
rect 18142 6695 18198 6704
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18248 6440 18276 22066
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 18290 18368 18566
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18340 11354 18368 11494
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 9586 18368 10202
rect 18328 9580 18380 9586
rect 18328 9522 18380 9528
rect 18432 8276 18460 22936
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18524 22166 18552 22374
rect 18512 22160 18564 22166
rect 18512 22102 18564 22108
rect 18616 21978 18644 24126
rect 18752 23964 19060 23973
rect 18752 23962 18758 23964
rect 18814 23962 18838 23964
rect 18894 23962 18918 23964
rect 18974 23962 18998 23964
rect 19054 23962 19060 23964
rect 18814 23910 18816 23962
rect 18996 23910 18998 23962
rect 18752 23908 18758 23910
rect 18814 23908 18838 23910
rect 18894 23908 18918 23910
rect 18974 23908 18998 23910
rect 19054 23908 19060 23910
rect 18752 23899 19060 23908
rect 19260 23866 19288 24142
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19352 23050 19380 27066
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 19720 26738 19748 36586
rect 19904 34354 19932 41074
rect 19996 41002 20024 43318
rect 20088 42129 20116 44463
rect 20364 43450 20392 44463
rect 20640 43450 20668 44463
rect 20720 43852 20772 43858
rect 20720 43794 20772 43800
rect 20352 43444 20404 43450
rect 20352 43386 20404 43392
rect 20628 43444 20680 43450
rect 20628 43386 20680 43392
rect 20444 43308 20496 43314
rect 20444 43250 20496 43256
rect 20260 42152 20312 42158
rect 20074 42120 20130 42129
rect 20260 42094 20312 42100
rect 20074 42055 20130 42064
rect 20272 41818 20300 42094
rect 20456 42090 20484 43250
rect 20536 42560 20588 42566
rect 20536 42502 20588 42508
rect 20444 42084 20496 42090
rect 20444 42026 20496 42032
rect 20548 41818 20576 42502
rect 20732 42242 20760 43794
rect 20916 43178 20944 44463
rect 21192 43450 21220 44463
rect 21272 43648 21324 43654
rect 21272 43590 21324 43596
rect 21180 43444 21232 43450
rect 21180 43386 21232 43392
rect 20904 43172 20956 43178
rect 20904 43114 20956 43120
rect 21284 42838 21312 43590
rect 21468 43364 21496 44463
rect 21548 43376 21600 43382
rect 21468 43336 21548 43364
rect 21548 43318 21600 43324
rect 21640 43308 21692 43314
rect 21640 43250 21692 43256
rect 21364 43104 21416 43110
rect 21364 43046 21416 43052
rect 21272 42832 21324 42838
rect 21272 42774 21324 42780
rect 20812 42628 20864 42634
rect 20812 42570 20864 42576
rect 21088 42628 21140 42634
rect 21088 42570 21140 42576
rect 20824 42362 20852 42570
rect 20996 42560 21048 42566
rect 20996 42502 21048 42508
rect 20812 42356 20864 42362
rect 20812 42298 20864 42304
rect 20732 42226 20852 42242
rect 20732 42220 20864 42226
rect 20732 42214 20812 42220
rect 20812 42162 20864 42168
rect 20904 42152 20956 42158
rect 20718 42120 20774 42129
rect 20904 42094 20956 42100
rect 20718 42055 20774 42064
rect 20732 41818 20760 42055
rect 20260 41812 20312 41818
rect 20260 41754 20312 41760
rect 20536 41812 20588 41818
rect 20536 41754 20588 41760
rect 20720 41812 20772 41818
rect 20720 41754 20772 41760
rect 20352 41744 20404 41750
rect 20350 41712 20352 41721
rect 20404 41712 20406 41721
rect 20350 41647 20406 41656
rect 20260 41608 20312 41614
rect 20260 41550 20312 41556
rect 20272 41274 20300 41550
rect 20260 41268 20312 41274
rect 20260 41210 20312 41216
rect 20536 41132 20588 41138
rect 20536 41074 20588 41080
rect 20444 41064 20496 41070
rect 20444 41006 20496 41012
rect 19984 40996 20036 41002
rect 19984 40938 20036 40944
rect 20260 40656 20312 40662
rect 20260 40598 20312 40604
rect 20168 40520 20220 40526
rect 20168 40462 20220 40468
rect 20076 40180 20128 40186
rect 20076 40122 20128 40128
rect 20088 40089 20116 40122
rect 20074 40080 20130 40089
rect 19984 40044 20036 40050
rect 20074 40015 20130 40024
rect 19984 39986 20036 39992
rect 19996 39409 20024 39986
rect 19982 39400 20038 39409
rect 19982 39335 20038 39344
rect 20076 39364 20128 39370
rect 20076 39306 20128 39312
rect 20088 38826 20116 39306
rect 20076 38820 20128 38826
rect 20076 38762 20128 38768
rect 20180 38010 20208 40462
rect 20272 40361 20300 40598
rect 20258 40352 20314 40361
rect 20258 40287 20314 40296
rect 20456 39506 20484 41006
rect 20444 39500 20496 39506
rect 20444 39442 20496 39448
rect 20444 39296 20496 39302
rect 20444 39238 20496 39244
rect 20456 39098 20484 39238
rect 20444 39092 20496 39098
rect 20444 39034 20496 39040
rect 20444 38888 20496 38894
rect 20442 38856 20444 38865
rect 20496 38856 20498 38865
rect 20442 38791 20498 38800
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 20260 37800 20312 37806
rect 20180 37760 20260 37788
rect 19984 34400 20036 34406
rect 19904 34348 19984 34354
rect 19904 34342 20036 34348
rect 19904 34326 20024 34342
rect 19904 34202 19932 34326
rect 19892 34196 19944 34202
rect 19892 34138 19944 34144
rect 20180 31346 20208 37760
rect 20260 37742 20312 37748
rect 20548 37126 20576 41074
rect 20812 40996 20864 41002
rect 20812 40938 20864 40944
rect 20628 40928 20680 40934
rect 20628 40870 20680 40876
rect 20720 40928 20772 40934
rect 20720 40870 20772 40876
rect 20640 40497 20668 40870
rect 20626 40488 20682 40497
rect 20626 40423 20682 40432
rect 20732 40118 20760 40870
rect 20824 40730 20852 40938
rect 20812 40724 20864 40730
rect 20812 40666 20864 40672
rect 20810 40216 20866 40225
rect 20810 40151 20866 40160
rect 20720 40112 20772 40118
rect 20720 40054 20772 40060
rect 20824 40050 20852 40151
rect 20812 40044 20864 40050
rect 20812 39986 20864 39992
rect 20812 39908 20864 39914
rect 20812 39850 20864 39856
rect 20824 39545 20852 39850
rect 20916 39642 20944 42094
rect 21008 40730 21036 42502
rect 21100 41274 21128 42570
rect 21272 42220 21324 42226
rect 21272 42162 21324 42168
rect 21180 42016 21232 42022
rect 21180 41958 21232 41964
rect 21192 41818 21220 41958
rect 21180 41812 21232 41818
rect 21180 41754 21232 41760
rect 21180 41608 21232 41614
rect 21180 41550 21232 41556
rect 21192 41274 21220 41550
rect 21284 41274 21312 42162
rect 21376 41818 21404 43046
rect 21548 42628 21600 42634
rect 21548 42570 21600 42576
rect 21364 41812 21416 41818
rect 21364 41754 21416 41760
rect 21362 41712 21418 41721
rect 21362 41647 21418 41656
rect 21376 41614 21404 41647
rect 21364 41608 21416 41614
rect 21364 41550 21416 41556
rect 21456 41472 21508 41478
rect 21456 41414 21508 41420
rect 21088 41268 21140 41274
rect 21088 41210 21140 41216
rect 21180 41268 21232 41274
rect 21180 41210 21232 41216
rect 21272 41268 21324 41274
rect 21272 41210 21324 41216
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 21180 41132 21232 41138
rect 21180 41074 21232 41080
rect 21364 41132 21416 41138
rect 21364 41074 21416 41080
rect 20996 40724 21048 40730
rect 20996 40666 21048 40672
rect 20996 40520 21048 40526
rect 20996 40462 21048 40468
rect 21008 39642 21036 40462
rect 21100 40202 21128 41074
rect 21192 40594 21220 41074
rect 21376 40594 21404 41074
rect 21180 40588 21232 40594
rect 21180 40530 21232 40536
rect 21364 40588 21416 40594
rect 21364 40530 21416 40536
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21100 40174 21220 40202
rect 21088 40044 21140 40050
rect 21088 39986 21140 39992
rect 21100 39846 21128 39986
rect 21088 39840 21140 39846
rect 21088 39782 21140 39788
rect 21192 39658 21220 40174
rect 20904 39636 20956 39642
rect 20904 39578 20956 39584
rect 20996 39636 21048 39642
rect 20996 39578 21048 39584
rect 21100 39630 21220 39658
rect 20810 39536 20866 39545
rect 20720 39500 20772 39506
rect 20810 39471 20866 39480
rect 20720 39442 20772 39448
rect 20628 38940 20680 38946
rect 20628 38882 20680 38888
rect 20640 38554 20668 38882
rect 20628 38548 20680 38554
rect 20628 38490 20680 38496
rect 20732 38486 20760 39442
rect 20904 39432 20956 39438
rect 20904 39374 20956 39380
rect 20812 39364 20864 39370
rect 20812 39306 20864 39312
rect 20824 38978 20852 39306
rect 20916 39098 20944 39374
rect 20904 39092 20956 39098
rect 20904 39034 20956 39040
rect 20824 38962 20944 38978
rect 20824 38956 20956 38962
rect 20824 38950 20904 38956
rect 20904 38898 20956 38904
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20720 38480 20772 38486
rect 20720 38422 20772 38428
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 20732 36922 20760 37198
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20536 36780 20588 36786
rect 20536 36722 20588 36728
rect 20548 36582 20576 36722
rect 20536 36576 20588 36582
rect 20536 36518 20588 36524
rect 20260 36168 20312 36174
rect 20260 36110 20312 36116
rect 20272 33998 20300 36110
rect 20444 34672 20496 34678
rect 20444 34614 20496 34620
rect 20456 34406 20484 34614
rect 20444 34400 20496 34406
rect 20444 34342 20496 34348
rect 20260 33992 20312 33998
rect 20260 33934 20312 33940
rect 20628 33108 20680 33114
rect 20628 33050 20680 33056
rect 20536 32224 20588 32230
rect 20536 32166 20588 32172
rect 20548 31958 20576 32166
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20640 31754 20668 33050
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20456 31726 20668 31754
rect 20732 31754 20760 31894
rect 20732 31726 20852 31754
rect 19800 31340 19852 31346
rect 19800 31282 19852 31288
rect 20168 31340 20220 31346
rect 20168 31282 20220 31288
rect 19812 29034 19840 31282
rect 19984 30048 20036 30054
rect 19984 29990 20036 29996
rect 19996 29510 20024 29990
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19800 29028 19852 29034
rect 19800 28970 19852 28976
rect 19812 27062 19840 28970
rect 19996 28558 20024 29446
rect 19984 28552 20036 28558
rect 20036 28512 20116 28540
rect 19984 28494 20036 28500
rect 19800 27056 19852 27062
rect 19800 26998 19852 27004
rect 20088 26994 20116 28512
rect 20076 26988 20128 26994
rect 19996 26948 20076 26976
rect 19444 26382 19472 26726
rect 19720 26710 19932 26738
rect 19708 26580 19760 26586
rect 19708 26522 19760 26528
rect 19524 26512 19576 26518
rect 19524 26454 19576 26460
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19444 25242 19472 25638
rect 19536 25430 19564 26454
rect 19616 26308 19668 26314
rect 19616 26250 19668 26256
rect 19524 25424 19576 25430
rect 19524 25366 19576 25372
rect 19444 25214 19564 25242
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 24886 19472 25094
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 19536 24256 19564 25214
rect 19444 24228 19564 24256
rect 19444 23526 19472 24228
rect 19628 24154 19656 26250
rect 19720 25242 19748 26522
rect 19720 25214 19840 25242
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19720 24954 19748 25094
rect 19708 24948 19760 24954
rect 19708 24890 19760 24896
rect 19706 24848 19762 24857
rect 19706 24783 19762 24792
rect 19536 24126 19656 24154
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19340 23044 19392 23050
rect 19340 22986 19392 22992
rect 18752 22876 19060 22885
rect 18752 22874 18758 22876
rect 18814 22874 18838 22876
rect 18894 22874 18918 22876
rect 18974 22874 18998 22876
rect 19054 22874 19060 22876
rect 18814 22822 18816 22874
rect 18996 22822 18998 22874
rect 18752 22820 18758 22822
rect 18814 22820 18838 22822
rect 18894 22820 18918 22822
rect 18974 22820 18998 22822
rect 19054 22820 19060 22822
rect 18752 22811 19060 22820
rect 19156 22228 19208 22234
rect 19444 22216 19472 23462
rect 19536 22778 19564 24126
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19628 23526 19656 24006
rect 19720 23866 19748 24783
rect 19708 23860 19760 23866
rect 19708 23802 19760 23808
rect 19616 23520 19668 23526
rect 19616 23462 19668 23468
rect 19628 23118 19656 23462
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19208 22188 19288 22216
rect 19444 22188 19564 22216
rect 19156 22170 19208 22176
rect 19260 22114 19288 22188
rect 19260 22086 19380 22114
rect 18524 21950 18644 21978
rect 19248 22024 19300 22030
rect 19352 22012 19380 22086
rect 19352 21984 19472 22012
rect 19248 21966 19300 21972
rect 18524 20466 18552 21950
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18616 21622 18644 21830
rect 18752 21788 19060 21797
rect 18752 21786 18758 21788
rect 18814 21786 18838 21788
rect 18894 21786 18918 21788
rect 18974 21786 18998 21788
rect 19054 21786 19060 21788
rect 18814 21734 18816 21786
rect 18996 21734 18998 21786
rect 18752 21732 18758 21734
rect 18814 21732 18838 21734
rect 18894 21732 18918 21734
rect 18974 21732 18998 21734
rect 19054 21732 19060 21734
rect 18752 21723 19060 21732
rect 18604 21616 18656 21622
rect 18604 21558 18656 21564
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18800 21010 18828 21286
rect 18788 21004 18840 21010
rect 18788 20946 18840 20952
rect 19156 20936 19208 20942
rect 19156 20878 19208 20884
rect 18752 20700 19060 20709
rect 18752 20698 18758 20700
rect 18814 20698 18838 20700
rect 18894 20698 18918 20700
rect 18974 20698 18998 20700
rect 19054 20698 19060 20700
rect 18814 20646 18816 20698
rect 18996 20646 18998 20698
rect 18752 20644 18758 20646
rect 18814 20644 18838 20646
rect 18894 20644 18918 20646
rect 18974 20644 18998 20646
rect 19054 20644 19060 20646
rect 18752 20635 19060 20644
rect 19168 20602 19196 20878
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 18970 18644 19654
rect 18752 19612 19060 19621
rect 18752 19610 18758 19612
rect 18814 19610 18838 19612
rect 18894 19610 18918 19612
rect 18974 19610 18998 19612
rect 19054 19610 19060 19612
rect 18814 19558 18816 19610
rect 18996 19558 18998 19610
rect 18752 19556 18758 19558
rect 18814 19556 18838 19558
rect 18894 19556 18918 19558
rect 18974 19556 18998 19558
rect 19054 19556 19060 19558
rect 18752 19547 19060 19556
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18752 18524 19060 18533
rect 18752 18522 18758 18524
rect 18814 18522 18838 18524
rect 18894 18522 18918 18524
rect 18974 18522 18998 18524
rect 19054 18522 19060 18524
rect 18814 18470 18816 18522
rect 18996 18470 18998 18522
rect 18752 18468 18758 18470
rect 18814 18468 18838 18470
rect 18894 18468 18918 18470
rect 18974 18468 18998 18470
rect 19054 18468 19060 18470
rect 18752 18459 19060 18468
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18524 15026 18552 17478
rect 18752 17436 19060 17445
rect 18752 17434 18758 17436
rect 18814 17434 18838 17436
rect 18894 17434 18918 17436
rect 18974 17434 18998 17436
rect 19054 17434 19060 17436
rect 18814 17382 18816 17434
rect 18996 17382 18998 17434
rect 18752 17380 18758 17382
rect 18814 17380 18838 17382
rect 18894 17380 18918 17382
rect 18974 17380 18998 17382
rect 19054 17380 19060 17382
rect 18752 17371 19060 17380
rect 19168 17252 19196 20402
rect 19260 19854 19288 21966
rect 19340 21412 19392 21418
rect 19340 21354 19392 21360
rect 19352 21010 19380 21354
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19444 18170 19472 21984
rect 19536 21554 19564 22188
rect 19812 22094 19840 25214
rect 19904 24834 19932 26710
rect 19996 25702 20024 26948
rect 20076 26930 20128 26936
rect 19984 25696 20036 25702
rect 19984 25638 20036 25644
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 19996 25362 20024 25638
rect 20088 25498 20116 25638
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20180 25378 20208 31282
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 20352 28960 20404 28966
rect 20352 28902 20404 28908
rect 20272 28801 20300 28902
rect 20258 28792 20314 28801
rect 20364 28762 20392 28902
rect 20258 28727 20314 28736
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20456 28642 20484 31726
rect 20640 31686 20668 31726
rect 20536 31680 20588 31686
rect 20536 31622 20588 31628
rect 20628 31680 20680 31686
rect 20628 31622 20680 31628
rect 20548 31498 20576 31622
rect 20548 31470 20760 31498
rect 20732 31346 20760 31470
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20628 31204 20680 31210
rect 20628 31146 20680 31152
rect 20640 30938 20668 31146
rect 20628 30932 20680 30938
rect 20628 30874 20680 30880
rect 20824 30734 20852 31726
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20536 30252 20588 30258
rect 20536 30194 20588 30200
rect 20548 29578 20576 30194
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20364 28614 20484 28642
rect 20364 28558 20392 28614
rect 20352 28552 20404 28558
rect 20352 28494 20404 28500
rect 20536 28416 20588 28422
rect 20536 28358 20588 28364
rect 20444 26512 20496 26518
rect 20444 26454 20496 26460
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20364 25498 20392 25706
rect 20352 25492 20404 25498
rect 20352 25434 20404 25440
rect 19984 25356 20036 25362
rect 20180 25350 20392 25378
rect 19984 25298 20036 25304
rect 19996 24954 20024 25298
rect 20076 25288 20128 25294
rect 20074 25256 20076 25265
rect 20128 25256 20130 25265
rect 20074 25191 20130 25200
rect 19984 24948 20036 24954
rect 19984 24890 20036 24896
rect 19904 24806 20024 24834
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23322 19932 24006
rect 19996 23798 20024 24806
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24206 20208 24754
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19984 23792 20036 23798
rect 19984 23734 20036 23740
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19812 22066 20024 22094
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19812 21554 19840 21966
rect 19892 21956 19944 21962
rect 19892 21898 19944 21904
rect 19524 21548 19576 21554
rect 19524 21490 19576 21496
rect 19800 21548 19852 21554
rect 19800 21490 19852 21496
rect 19536 19446 19564 21490
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19628 21146 19656 21286
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19616 20528 19668 20534
rect 19616 20470 19668 20476
rect 19628 19446 19656 20470
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 19444 18142 19564 18170
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19444 17610 19472 18022
rect 19432 17604 19484 17610
rect 19432 17546 19484 17552
rect 19444 17338 19472 17546
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19168 17224 19288 17252
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14618 18552 14758
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18524 13530 18552 14214
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18616 12850 18644 16526
rect 18752 16348 19060 16357
rect 18752 16346 18758 16348
rect 18814 16346 18838 16348
rect 18894 16346 18918 16348
rect 18974 16346 18998 16348
rect 19054 16346 19060 16348
rect 18814 16294 18816 16346
rect 18996 16294 18998 16346
rect 18752 16292 18758 16294
rect 18814 16292 18838 16294
rect 18894 16292 18918 16294
rect 18974 16292 18998 16294
rect 19054 16292 19060 16294
rect 18752 16283 19060 16292
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18892 15706 18920 16050
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18752 15260 19060 15269
rect 18752 15258 18758 15260
rect 18814 15258 18838 15260
rect 18894 15258 18918 15260
rect 18974 15258 18998 15260
rect 19054 15258 19060 15260
rect 18814 15206 18816 15258
rect 18996 15206 18998 15258
rect 18752 15204 18758 15206
rect 18814 15204 18838 15206
rect 18894 15204 18918 15206
rect 18974 15204 18998 15206
rect 19054 15204 19060 15206
rect 18752 15195 19060 15204
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 18752 14172 19060 14181
rect 18752 14170 18758 14172
rect 18814 14170 18838 14172
rect 18894 14170 18918 14172
rect 18974 14170 18998 14172
rect 19054 14170 19060 14172
rect 18814 14118 18816 14170
rect 18996 14118 18998 14170
rect 18752 14116 18758 14118
rect 18814 14116 18838 14118
rect 18894 14116 18918 14118
rect 18974 14116 18998 14118
rect 19054 14116 19060 14118
rect 18752 14107 19060 14116
rect 19168 14006 19196 14214
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19156 13864 19208 13870
rect 18984 13812 19156 13818
rect 18984 13806 19208 13812
rect 18880 13796 18932 13802
rect 18880 13738 18932 13744
rect 18984 13790 19196 13806
rect 18892 13326 18920 13738
rect 18984 13394 19012 13790
rect 19260 13682 19288 17224
rect 19536 15994 19564 18142
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19444 15966 19564 15994
rect 19340 15428 19392 15434
rect 19340 15370 19392 15376
rect 19352 15162 19380 15370
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19168 13654 19288 13682
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18752 13084 19060 13093
rect 18752 13082 18758 13084
rect 18814 13082 18838 13084
rect 18894 13082 18918 13084
rect 18974 13082 18998 13084
rect 19054 13082 19060 13084
rect 18814 13030 18816 13082
rect 18996 13030 18998 13082
rect 18752 13028 18758 13030
rect 18814 13028 18838 13030
rect 18894 13028 18918 13030
rect 18974 13028 18998 13030
rect 19054 13028 19060 13030
rect 18752 13019 19060 13028
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 19168 12434 19196 13654
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19260 12714 19288 13126
rect 19352 12918 19380 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19248 12708 19300 12714
rect 19248 12650 19300 12656
rect 18064 6412 18276 6440
rect 18340 8248 18460 8276
rect 18524 12406 19196 12434
rect 17958 6216 18014 6225
rect 17958 6151 18014 6160
rect 17868 6112 17920 6118
rect 17868 6054 17920 6060
rect 17880 5642 17908 6054
rect 17958 5672 18014 5681
rect 17868 5636 17920 5642
rect 17958 5607 18014 5616
rect 17868 5578 17920 5584
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 17972 5098 18000 5607
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17144 4134 17264 4162
rect 17880 4146 17908 4490
rect 17958 4176 18014 4185
rect 17868 4140 17920 4146
rect 17038 2816 17094 2825
rect 17038 2751 17094 2760
rect 17144 2774 17172 4134
rect 17958 4111 18014 4120
rect 17868 4082 17920 4088
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17236 2938 17264 2994
rect 17604 2990 17632 3674
rect 17972 3618 18000 4111
rect 17788 3590 18000 3618
rect 17788 3482 17816 3590
rect 18064 3516 18092 6412
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5370 18184 6122
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18248 5370 18276 5850
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18340 4146 18368 8248
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18432 7546 18460 8026
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18432 5370 18460 6190
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 18524 5250 18552 12406
rect 18752 11996 19060 12005
rect 18752 11994 18758 11996
rect 18814 11994 18838 11996
rect 18894 11994 18918 11996
rect 18974 11994 18998 11996
rect 19054 11994 19060 11996
rect 18814 11942 18816 11994
rect 18996 11942 18998 11994
rect 18752 11940 18758 11942
rect 18814 11940 18838 11942
rect 18894 11940 18918 11942
rect 18974 11940 18998 11942
rect 19054 11940 19060 11942
rect 18752 11931 19060 11940
rect 19444 11801 19472 15966
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19536 15026 19564 15846
rect 19628 15094 19656 17478
rect 19616 15088 19668 15094
rect 19616 15030 19668 15036
rect 19524 15020 19576 15026
rect 19524 14962 19576 14968
rect 19524 13456 19576 13462
rect 19522 13424 19524 13433
rect 19576 13424 19578 13433
rect 19522 13359 19578 13368
rect 19720 12434 19748 20742
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 15978 19840 19314
rect 19904 17134 19932 21898
rect 19892 17128 19944 17134
rect 19892 17070 19944 17076
rect 19904 16794 19932 17070
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19996 16425 20024 22066
rect 20088 22030 20116 22714
rect 20260 22092 20312 22098
rect 20260 22034 20312 22040
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20272 21690 20300 22034
rect 20364 21962 20392 25350
rect 20352 21956 20404 21962
rect 20352 21898 20404 21904
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20456 21162 20484 26454
rect 20548 26382 20576 28358
rect 20732 28098 20760 29786
rect 20640 28070 20760 28098
rect 20640 27452 20668 28070
rect 20720 28008 20772 28014
rect 20720 27950 20772 27956
rect 20732 27606 20760 27950
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 27606 20852 27814
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20640 27424 20760 27452
rect 20732 27010 20760 27424
rect 20916 27146 20944 38694
rect 21100 38554 21128 39630
rect 21180 39568 21232 39574
rect 21180 39510 21232 39516
rect 21192 39030 21220 39510
rect 21180 39024 21232 39030
rect 21180 38966 21232 38972
rect 21284 38654 21312 40462
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21376 39574 21404 39986
rect 21364 39568 21416 39574
rect 21364 39510 21416 39516
rect 21468 39438 21496 41414
rect 21560 41138 21588 42570
rect 21652 42362 21680 43250
rect 21744 43092 21772 44463
rect 22020 43160 22048 44463
rect 22192 43172 22244 43178
rect 22020 43132 22140 43160
rect 21916 43104 21968 43110
rect 21744 43064 21916 43092
rect 21916 43046 21968 43052
rect 21719 43004 22027 43013
rect 21719 43002 21725 43004
rect 21781 43002 21805 43004
rect 21861 43002 21885 43004
rect 21941 43002 21965 43004
rect 22021 43002 22027 43004
rect 21781 42950 21783 43002
rect 21963 42950 21965 43002
rect 21719 42948 21725 42950
rect 21781 42948 21805 42950
rect 21861 42948 21885 42950
rect 21941 42948 21965 42950
rect 22021 42948 22027 42950
rect 21719 42939 22027 42948
rect 22112 42786 22140 43132
rect 22192 43114 22244 43120
rect 21928 42758 22140 42786
rect 21928 42702 21956 42758
rect 21916 42696 21968 42702
rect 22204 42650 22232 43114
rect 22296 42770 22324 44463
rect 22376 43308 22428 43314
rect 22376 43250 22428 43256
rect 22388 42838 22416 43250
rect 22572 43246 22600 44463
rect 22652 43308 22704 43314
rect 22652 43250 22704 43256
rect 22560 43240 22612 43246
rect 22560 43182 22612 43188
rect 22376 42832 22428 42838
rect 22376 42774 22428 42780
rect 22284 42764 22336 42770
rect 22284 42706 22336 42712
rect 21916 42638 21968 42644
rect 22112 42622 22232 42650
rect 21916 42560 21968 42566
rect 21968 42520 22048 42548
rect 21916 42502 21968 42508
rect 21640 42356 21692 42362
rect 21640 42298 21692 42304
rect 21914 42120 21970 42129
rect 22020 42090 22048 42520
rect 21914 42055 21916 42064
rect 21968 42055 21970 42064
rect 22008 42084 22060 42090
rect 21916 42026 21968 42032
rect 22008 42026 22060 42032
rect 21719 41916 22027 41925
rect 21719 41914 21725 41916
rect 21781 41914 21805 41916
rect 21861 41914 21885 41916
rect 21941 41914 21965 41916
rect 22021 41914 22027 41916
rect 21781 41862 21783 41914
rect 21963 41862 21965 41914
rect 21719 41860 21725 41862
rect 21781 41860 21805 41862
rect 21861 41860 21885 41862
rect 21941 41860 21965 41862
rect 22021 41860 22027 41862
rect 21719 41851 22027 41860
rect 21640 41608 21692 41614
rect 21638 41576 21640 41585
rect 21692 41576 21694 41585
rect 22112 41562 22140 42622
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22204 42226 22232 42502
rect 22192 42220 22244 42226
rect 22192 42162 22244 42168
rect 22284 41812 22336 41818
rect 22284 41754 22336 41760
rect 21638 41511 21694 41520
rect 21824 41540 21876 41546
rect 21824 41482 21876 41488
rect 22020 41534 22140 41562
rect 21836 41414 21864 41482
rect 21652 41386 21864 41414
rect 21548 41132 21600 41138
rect 21548 41074 21600 41080
rect 21546 41032 21602 41041
rect 21546 40967 21602 40976
rect 21560 40202 21588 40967
rect 21652 40390 21680 41386
rect 21732 41268 21784 41274
rect 21732 41210 21784 41216
rect 21744 41177 21772 41210
rect 21730 41168 21786 41177
rect 21730 41103 21786 41112
rect 21916 41132 21968 41138
rect 21916 41074 21968 41080
rect 21928 40934 21956 41074
rect 22020 41002 22048 41534
rect 22296 41274 22324 41754
rect 22376 41472 22428 41478
rect 22376 41414 22428 41420
rect 22284 41268 22336 41274
rect 22284 41210 22336 41216
rect 22100 41200 22152 41206
rect 22100 41142 22152 41148
rect 22008 40996 22060 41002
rect 22008 40938 22060 40944
rect 21916 40928 21968 40934
rect 21916 40870 21968 40876
rect 21719 40828 22027 40837
rect 21719 40826 21725 40828
rect 21781 40826 21805 40828
rect 21861 40826 21885 40828
rect 21941 40826 21965 40828
rect 22021 40826 22027 40828
rect 21781 40774 21783 40826
rect 21963 40774 21965 40826
rect 21719 40772 21725 40774
rect 21781 40772 21805 40774
rect 21861 40772 21885 40774
rect 21941 40772 21965 40774
rect 22021 40772 22027 40774
rect 21719 40763 22027 40772
rect 22112 40730 22140 41142
rect 22192 41132 22244 41138
rect 22192 41074 22244 41080
rect 22100 40724 22152 40730
rect 22100 40666 22152 40672
rect 21732 40452 21784 40458
rect 21732 40394 21784 40400
rect 21640 40384 21692 40390
rect 21640 40326 21692 40332
rect 21560 40174 21680 40202
rect 21548 40112 21600 40118
rect 21548 40054 21600 40060
rect 21456 39432 21508 39438
rect 21456 39374 21508 39380
rect 21456 39296 21508 39302
rect 21456 39238 21508 39244
rect 21468 39098 21496 39238
rect 21456 39092 21508 39098
rect 21456 39034 21508 39040
rect 21192 38626 21312 38654
rect 21088 38548 21140 38554
rect 21088 38490 21140 38496
rect 21088 34536 21140 34542
rect 21088 34478 21140 34484
rect 21100 34202 21128 34478
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 20996 33652 21048 33658
rect 20996 33594 21048 33600
rect 21008 33522 21036 33594
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21192 31686 21220 38626
rect 21560 37856 21588 40054
rect 21652 39846 21680 40174
rect 21744 40050 21772 40394
rect 21732 40044 21784 40050
rect 21732 39986 21784 39992
rect 21640 39840 21692 39846
rect 21640 39782 21692 39788
rect 21719 39740 22027 39749
rect 21719 39738 21725 39740
rect 21781 39738 21805 39740
rect 21861 39738 21885 39740
rect 21941 39738 21965 39740
rect 22021 39738 22027 39740
rect 21781 39686 21783 39738
rect 21963 39686 21965 39738
rect 21719 39684 21725 39686
rect 21781 39684 21805 39686
rect 21861 39684 21885 39686
rect 21941 39684 21965 39686
rect 22021 39684 22027 39686
rect 21719 39675 22027 39684
rect 22204 39642 22232 41074
rect 22388 40984 22416 41414
rect 22560 41132 22612 41138
rect 22560 41074 22612 41080
rect 22388 40956 22508 40984
rect 22284 40928 22336 40934
rect 22284 40870 22336 40876
rect 22296 40458 22324 40870
rect 22376 40520 22428 40526
rect 22376 40462 22428 40468
rect 22284 40452 22336 40458
rect 22284 40394 22336 40400
rect 22282 39944 22338 39953
rect 22282 39879 22338 39888
rect 22296 39846 22324 39879
rect 22284 39840 22336 39846
rect 22284 39782 22336 39788
rect 22388 39642 22416 40462
rect 22480 40372 22508 40956
rect 22572 40730 22600 41074
rect 22664 41002 22692 43250
rect 22848 42362 22876 44463
rect 23124 43450 23152 44463
rect 23112 43444 23164 43450
rect 23112 43386 23164 43392
rect 23202 43344 23258 43353
rect 23202 43279 23258 43288
rect 23020 42832 23072 42838
rect 23020 42774 23072 42780
rect 22836 42356 22888 42362
rect 22836 42298 22888 42304
rect 22836 42220 22888 42226
rect 22836 42162 22888 42168
rect 22744 41064 22796 41070
rect 22744 41006 22796 41012
rect 22652 40996 22704 41002
rect 22652 40938 22704 40944
rect 22756 40730 22784 41006
rect 22560 40724 22612 40730
rect 22560 40666 22612 40672
rect 22744 40724 22796 40730
rect 22744 40666 22796 40672
rect 22650 40624 22706 40633
rect 22650 40559 22706 40568
rect 22744 40588 22796 40594
rect 22664 40526 22692 40559
rect 22744 40530 22796 40536
rect 22652 40520 22704 40526
rect 22652 40462 22704 40468
rect 22756 40372 22784 40530
rect 22480 40344 22784 40372
rect 22468 40044 22520 40050
rect 22468 39986 22520 39992
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22376 39636 22428 39642
rect 22376 39578 22428 39584
rect 22008 39432 22060 39438
rect 21284 37828 21588 37856
rect 21652 39392 22008 39420
rect 21284 32978 21312 37828
rect 21652 37754 21680 39392
rect 22008 39374 22060 39380
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 21824 38888 21876 38894
rect 21822 38856 21824 38865
rect 21876 38856 21878 38865
rect 21822 38791 21878 38800
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 21719 38652 22027 38661
rect 21719 38650 21725 38652
rect 21781 38650 21805 38652
rect 21861 38650 21885 38652
rect 21941 38650 21965 38652
rect 22021 38650 22027 38652
rect 21781 38598 21783 38650
rect 21963 38598 21965 38650
rect 21719 38596 21725 38598
rect 21781 38596 21805 38598
rect 21861 38596 21885 38598
rect 21941 38596 21965 38598
rect 22021 38596 22027 38598
rect 21719 38587 22027 38596
rect 22112 38350 22140 38694
rect 22100 38344 22152 38350
rect 22100 38286 22152 38292
rect 22192 38208 22244 38214
rect 22192 38150 22244 38156
rect 22204 38010 22232 38150
rect 22192 38004 22244 38010
rect 22192 37946 22244 37952
rect 21376 37726 21680 37754
rect 21272 32972 21324 32978
rect 21272 32914 21324 32920
rect 21376 31754 21404 37726
rect 21640 37664 21692 37670
rect 21640 37606 21692 37612
rect 21652 37466 21680 37606
rect 21719 37564 22027 37573
rect 21719 37562 21725 37564
rect 21781 37562 21805 37564
rect 21861 37562 21885 37564
rect 21941 37562 21965 37564
rect 22021 37562 22027 37564
rect 21781 37510 21783 37562
rect 21963 37510 21965 37562
rect 21719 37508 21725 37510
rect 21781 37508 21805 37510
rect 21861 37508 21885 37510
rect 21941 37508 21965 37510
rect 22021 37508 22027 37510
rect 21719 37499 22027 37508
rect 21640 37460 21692 37466
rect 21640 37402 21692 37408
rect 22296 37330 22324 39374
rect 22284 37324 22336 37330
rect 22284 37266 22336 37272
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22192 37256 22244 37262
rect 22192 37198 22244 37204
rect 21836 36922 21864 37198
rect 21824 36916 21876 36922
rect 21824 36858 21876 36864
rect 21719 36476 22027 36485
rect 21719 36474 21725 36476
rect 21781 36474 21805 36476
rect 21861 36474 21885 36476
rect 21941 36474 21965 36476
rect 22021 36474 22027 36476
rect 21781 36422 21783 36474
rect 21963 36422 21965 36474
rect 21719 36420 21725 36422
rect 21781 36420 21805 36422
rect 21861 36420 21885 36422
rect 21941 36420 21965 36422
rect 22021 36420 22027 36422
rect 21719 36411 22027 36420
rect 22112 36378 22140 37198
rect 22204 37126 22232 37198
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 22100 36372 22152 36378
rect 22100 36314 22152 36320
rect 21719 35388 22027 35397
rect 21719 35386 21725 35388
rect 21781 35386 21805 35388
rect 21861 35386 21885 35388
rect 21941 35386 21965 35388
rect 22021 35386 22027 35388
rect 21781 35334 21783 35386
rect 21963 35334 21965 35386
rect 21719 35332 21725 35334
rect 21781 35332 21805 35334
rect 21861 35332 21885 35334
rect 21941 35332 21965 35334
rect 22021 35332 22027 35334
rect 21719 35323 22027 35332
rect 22204 34610 22232 37062
rect 22376 36712 22428 36718
rect 22376 36654 22428 36660
rect 22388 36378 22416 36654
rect 22376 36372 22428 36378
rect 22376 36314 22428 36320
rect 22480 35290 22508 39986
rect 22848 39914 22876 42162
rect 23032 40730 23060 42774
rect 23216 42362 23244 43279
rect 23204 42356 23256 42362
rect 23204 42298 23256 42304
rect 23400 41274 23428 44463
rect 23480 43308 23532 43314
rect 23480 43250 23532 43256
rect 23492 42022 23520 43250
rect 23570 42120 23626 42129
rect 23570 42055 23626 42064
rect 23480 42016 23532 42022
rect 23480 41958 23532 41964
rect 23584 41614 23612 42055
rect 23572 41608 23624 41614
rect 23572 41550 23624 41556
rect 23676 41478 23704 44463
rect 23756 42628 23808 42634
rect 23756 42570 23808 42576
rect 23664 41472 23716 41478
rect 23664 41414 23716 41420
rect 23388 41268 23440 41274
rect 23388 41210 23440 41216
rect 23112 41132 23164 41138
rect 23112 41074 23164 41080
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 22928 40520 22980 40526
rect 22926 40488 22928 40497
rect 22980 40488 22982 40497
rect 22926 40423 22982 40432
rect 22928 40384 22980 40390
rect 22928 40326 22980 40332
rect 22836 39908 22888 39914
rect 22836 39850 22888 39856
rect 22940 39846 22968 40326
rect 23018 40216 23074 40225
rect 23018 40151 23074 40160
rect 23032 40050 23060 40151
rect 23124 40089 23152 41074
rect 23204 41064 23256 41070
rect 23768 41041 23796 42570
rect 23952 41818 23980 44463
rect 24124 43104 24176 43110
rect 24124 43046 24176 43052
rect 24032 42220 24084 42226
rect 24032 42162 24084 42168
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 23848 41540 23900 41546
rect 23848 41482 23900 41488
rect 23204 41006 23256 41012
rect 23754 41032 23810 41041
rect 23110 40080 23166 40089
rect 23020 40044 23072 40050
rect 23110 40015 23166 40024
rect 23020 39986 23072 39992
rect 23216 39953 23244 41006
rect 23754 40967 23810 40976
rect 23664 40928 23716 40934
rect 23662 40896 23664 40905
rect 23716 40896 23718 40905
rect 23662 40831 23718 40840
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23676 40361 23704 40462
rect 23662 40352 23718 40361
rect 23662 40287 23718 40296
rect 23860 40186 23888 41482
rect 23940 41472 23992 41478
rect 23940 41414 23992 41420
rect 23952 40202 23980 41414
rect 24044 40730 24072 42162
rect 24136 41993 24164 43046
rect 24228 42702 24256 44463
rect 24400 43648 24452 43654
rect 24400 43590 24452 43596
rect 24216 42696 24268 42702
rect 24216 42638 24268 42644
rect 24412 42242 24440 43590
rect 24504 42362 24532 44463
rect 24780 43738 24808 44463
rect 24596 43710 24808 43738
rect 24596 42702 24624 43710
rect 24686 43548 24994 43557
rect 24686 43546 24692 43548
rect 24748 43546 24772 43548
rect 24828 43546 24852 43548
rect 24908 43546 24932 43548
rect 24988 43546 24994 43548
rect 24748 43494 24750 43546
rect 24930 43494 24932 43546
rect 24686 43492 24692 43494
rect 24748 43492 24772 43494
rect 24828 43492 24852 43494
rect 24908 43492 24932 43494
rect 24988 43492 24994 43494
rect 24686 43483 24994 43492
rect 24584 42696 24636 42702
rect 24584 42638 24636 42644
rect 24686 42460 24994 42469
rect 24686 42458 24692 42460
rect 24748 42458 24772 42460
rect 24828 42458 24852 42460
rect 24908 42458 24932 42460
rect 24988 42458 24994 42460
rect 24748 42406 24750 42458
rect 24930 42406 24932 42458
rect 24686 42404 24692 42406
rect 24748 42404 24772 42406
rect 24828 42404 24852 42406
rect 24908 42404 24932 42406
rect 24988 42404 24994 42406
rect 24686 42395 24994 42404
rect 24492 42356 24544 42362
rect 24492 42298 24544 42304
rect 24584 42288 24636 42294
rect 24412 42214 24532 42242
rect 24584 42230 24636 42236
rect 24216 42084 24268 42090
rect 24216 42026 24268 42032
rect 24122 41984 24178 41993
rect 24122 41919 24178 41928
rect 24032 40724 24084 40730
rect 24032 40666 24084 40672
rect 23848 40180 23900 40186
rect 23952 40174 24164 40202
rect 23848 40122 23900 40128
rect 23756 40044 23808 40050
rect 23756 39986 23808 39992
rect 24032 40044 24084 40050
rect 24032 39986 24084 39992
rect 23202 39944 23258 39953
rect 23020 39908 23072 39914
rect 23202 39879 23258 39888
rect 23020 39850 23072 39856
rect 22928 39840 22980 39846
rect 22928 39782 22980 39788
rect 22836 39636 22888 39642
rect 22836 39578 22888 39584
rect 22560 39432 22612 39438
rect 22848 39409 22876 39578
rect 23032 39545 23060 39850
rect 23018 39536 23074 39545
rect 23018 39471 23074 39480
rect 22560 39374 22612 39380
rect 22834 39400 22890 39409
rect 22572 37942 22600 39374
rect 22834 39335 22890 39344
rect 23572 38956 23624 38962
rect 23572 38898 23624 38904
rect 23664 38956 23716 38962
rect 23664 38898 23716 38904
rect 23480 38820 23532 38826
rect 23480 38762 23532 38768
rect 22928 38548 22980 38554
rect 22928 38490 22980 38496
rect 22744 38480 22796 38486
rect 22744 38422 22796 38428
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22560 37936 22612 37942
rect 22560 37878 22612 37884
rect 22664 37466 22692 38286
rect 22756 38010 22784 38422
rect 22940 38350 22968 38490
rect 23112 38412 23164 38418
rect 23112 38354 23164 38360
rect 22928 38344 22980 38350
rect 22928 38286 22980 38292
rect 23020 38276 23072 38282
rect 23020 38218 23072 38224
rect 22836 38208 22888 38214
rect 22836 38150 22888 38156
rect 22928 38208 22980 38214
rect 22928 38150 22980 38156
rect 22744 38004 22796 38010
rect 22744 37946 22796 37952
rect 22848 37738 22876 38150
rect 22940 38010 22968 38150
rect 22928 38004 22980 38010
rect 22928 37946 22980 37952
rect 22928 37800 22980 37806
rect 22928 37742 22980 37748
rect 22836 37732 22888 37738
rect 22836 37674 22888 37680
rect 22652 37460 22704 37466
rect 22652 37402 22704 37408
rect 22744 37256 22796 37262
rect 22744 37198 22796 37204
rect 22756 36009 22784 37198
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22848 36378 22876 36518
rect 22836 36372 22888 36378
rect 22836 36314 22888 36320
rect 22742 36000 22798 36009
rect 22742 35935 22798 35944
rect 22468 35284 22520 35290
rect 22468 35226 22520 35232
rect 22192 34604 22244 34610
rect 22192 34546 22244 34552
rect 21548 34400 21600 34406
rect 21548 34342 21600 34348
rect 21560 33998 21588 34342
rect 21719 34300 22027 34309
rect 21719 34298 21725 34300
rect 21781 34298 21805 34300
rect 21861 34298 21885 34300
rect 21941 34298 21965 34300
rect 22021 34298 22027 34300
rect 21781 34246 21783 34298
rect 21963 34246 21965 34298
rect 21719 34244 21725 34246
rect 21781 34244 21805 34246
rect 21861 34244 21885 34246
rect 21941 34244 21965 34246
rect 22021 34244 22027 34246
rect 21719 34235 22027 34244
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 22560 33992 22612 33998
rect 22560 33934 22612 33940
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 21640 33856 21692 33862
rect 21640 33798 21692 33804
rect 21546 31920 21602 31929
rect 21652 31906 21680 33798
rect 22374 33552 22430 33561
rect 22374 33487 22430 33496
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 21719 33212 22027 33221
rect 21719 33210 21725 33212
rect 21781 33210 21805 33212
rect 21861 33210 21885 33212
rect 21941 33210 21965 33212
rect 22021 33210 22027 33212
rect 21781 33158 21783 33210
rect 21963 33158 21965 33210
rect 21719 33156 21725 33158
rect 21781 33156 21805 33158
rect 21861 33156 21885 33158
rect 21941 33156 21965 33158
rect 22021 33156 22027 33158
rect 21719 33147 22027 33156
rect 22204 32910 22232 33254
rect 22100 32904 22152 32910
rect 22100 32846 22152 32852
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 21719 32124 22027 32133
rect 21719 32122 21725 32124
rect 21781 32122 21805 32124
rect 21861 32122 21885 32124
rect 21941 32122 21965 32124
rect 22021 32122 22027 32124
rect 21781 32070 21783 32122
rect 21963 32070 21965 32122
rect 21719 32068 21725 32070
rect 21781 32068 21805 32070
rect 21861 32068 21885 32070
rect 21941 32068 21965 32070
rect 22021 32068 22027 32070
rect 21719 32059 22027 32068
rect 21652 31890 21772 31906
rect 21652 31884 21784 31890
rect 21652 31878 21732 31884
rect 21546 31855 21602 31864
rect 21284 31726 21404 31754
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 21008 28218 21036 28358
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 21088 28212 21140 28218
rect 21088 28154 21140 28160
rect 21100 27606 21128 28154
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 21180 27464 21232 27470
rect 21180 27406 21232 27412
rect 21192 27334 21220 27406
rect 21180 27328 21232 27334
rect 21180 27270 21232 27276
rect 20916 27118 21128 27146
rect 21100 27062 21128 27118
rect 21088 27056 21140 27062
rect 20732 26982 20944 27010
rect 21088 26998 21140 27004
rect 20810 26888 20866 26897
rect 20810 26823 20866 26832
rect 20536 26376 20588 26382
rect 20720 26376 20772 26382
rect 20536 26318 20588 26324
rect 20718 26344 20720 26353
rect 20772 26344 20774 26353
rect 20718 26279 20774 26288
rect 20720 25968 20772 25974
rect 20720 25910 20772 25916
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 23118 20668 24550
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20548 22778 20576 22986
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20640 22234 20668 23054
rect 20732 22234 20760 25910
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20824 22094 20852 26823
rect 20916 24070 20944 26982
rect 21088 26920 21140 26926
rect 21008 26880 21088 26908
rect 21008 24154 21036 26880
rect 21088 26862 21140 26868
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21100 24274 21128 25638
rect 21192 25294 21220 27270
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 21192 24614 21220 25230
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21284 24290 21312 31726
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21376 30433 21404 31078
rect 21468 30938 21496 31282
rect 21456 30932 21508 30938
rect 21456 30874 21508 30880
rect 21362 30424 21418 30433
rect 21362 30359 21418 30368
rect 21560 26926 21588 31855
rect 21732 31826 21784 31832
rect 21719 31036 22027 31045
rect 21719 31034 21725 31036
rect 21781 31034 21805 31036
rect 21861 31034 21885 31036
rect 21941 31034 21965 31036
rect 22021 31034 22027 31036
rect 21781 30982 21783 31034
rect 21963 30982 21965 31034
rect 21719 30980 21725 30982
rect 21781 30980 21805 30982
rect 21861 30980 21885 30982
rect 21941 30980 21965 30982
rect 22021 30980 22027 30982
rect 21719 30971 22027 30980
rect 21719 29948 22027 29957
rect 21719 29946 21725 29948
rect 21781 29946 21805 29948
rect 21861 29946 21885 29948
rect 21941 29946 21965 29948
rect 22021 29946 22027 29948
rect 21781 29894 21783 29946
rect 21963 29894 21965 29946
rect 21719 29892 21725 29894
rect 21781 29892 21805 29894
rect 21861 29892 21885 29894
rect 21941 29892 21965 29894
rect 22021 29892 22027 29894
rect 21719 29883 22027 29892
rect 22112 28994 22140 32846
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22204 31346 22232 31418
rect 22192 31340 22244 31346
rect 22192 31282 22244 31288
rect 22204 30258 22232 31282
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22296 30054 22324 30670
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22112 28966 22324 28994
rect 21719 28860 22027 28869
rect 21719 28858 21725 28860
rect 21781 28858 21805 28860
rect 21861 28858 21885 28860
rect 21941 28858 21965 28860
rect 22021 28858 22027 28860
rect 21781 28806 21783 28858
rect 21963 28806 21965 28858
rect 21719 28804 21725 28806
rect 21781 28804 21805 28806
rect 21861 28804 21885 28806
rect 21941 28804 21965 28806
rect 22021 28804 22027 28806
rect 21719 28795 22027 28804
rect 22192 28144 22244 28150
rect 22190 28112 22192 28121
rect 22244 28112 22246 28121
rect 22100 28076 22152 28082
rect 22190 28047 22246 28056
rect 22100 28018 22152 28024
rect 21719 27772 22027 27781
rect 21719 27770 21725 27772
rect 21781 27770 21805 27772
rect 21861 27770 21885 27772
rect 21941 27770 21965 27772
rect 22021 27770 22027 27772
rect 21781 27718 21783 27770
rect 21963 27718 21965 27770
rect 21719 27716 21725 27718
rect 21781 27716 21805 27718
rect 21861 27716 21885 27718
rect 21941 27716 21965 27718
rect 22021 27716 22027 27718
rect 21719 27707 22027 27716
rect 22112 27554 22140 28018
rect 22020 27526 22140 27554
rect 22020 27402 22048 27526
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21376 25498 21404 25842
rect 21456 25696 21508 25702
rect 21456 25638 21508 25644
rect 21364 25492 21416 25498
rect 21364 25434 21416 25440
rect 21376 24818 21404 25434
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21468 24732 21496 25638
rect 21560 24954 21588 25842
rect 21548 24948 21600 24954
rect 21548 24890 21600 24896
rect 21548 24744 21600 24750
rect 21468 24704 21548 24732
rect 21548 24686 21600 24692
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21468 24410 21496 24550
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21088 24268 21140 24274
rect 21284 24262 21588 24290
rect 21088 24210 21140 24216
rect 21008 24126 21128 24154
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20732 22080 20852 22094
rect 20088 21134 20484 21162
rect 20640 22066 20852 22080
rect 20640 22052 20760 22066
rect 19982 16416 20038 16425
rect 19982 16351 20038 16360
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 15026 19840 15302
rect 19800 15020 19852 15026
rect 19800 14962 19852 14968
rect 19720 12406 19840 12434
rect 19430 11792 19486 11801
rect 19430 11727 19486 11736
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11354 19104 11494
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18616 10266 18644 11086
rect 18752 10908 19060 10917
rect 18752 10906 18758 10908
rect 18814 10906 18838 10908
rect 18894 10906 18918 10908
rect 18974 10906 18998 10908
rect 19054 10906 19060 10908
rect 18814 10854 18816 10906
rect 18996 10854 18998 10906
rect 18752 10852 18758 10854
rect 18814 10852 18838 10854
rect 18894 10852 18918 10854
rect 18974 10852 18998 10854
rect 19054 10852 19060 10854
rect 18752 10843 19060 10852
rect 19064 10804 19116 10810
rect 19168 10792 19196 11562
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19246 11112 19302 11121
rect 19246 11047 19302 11056
rect 19116 10764 19196 10792
rect 19064 10746 19116 10752
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 19076 10198 19104 10542
rect 19156 10464 19208 10470
rect 19156 10406 19208 10412
rect 19168 10266 19196 10406
rect 19156 10260 19208 10266
rect 19156 10202 19208 10208
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 18752 9820 19060 9829
rect 18752 9818 18758 9820
rect 18814 9818 18838 9820
rect 18894 9818 18918 9820
rect 18974 9818 18998 9820
rect 19054 9818 19060 9820
rect 18814 9766 18816 9818
rect 18996 9766 18998 9818
rect 18752 9764 18758 9766
rect 18814 9764 18838 9766
rect 18894 9764 18918 9766
rect 18974 9764 18998 9766
rect 19054 9764 19060 9766
rect 18752 9755 19060 9764
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18616 8498 18644 8842
rect 18752 8732 19060 8741
rect 18752 8730 18758 8732
rect 18814 8730 18838 8732
rect 18894 8730 18918 8732
rect 18974 8730 18998 8732
rect 19054 8730 19060 8732
rect 18814 8678 18816 8730
rect 18996 8678 18998 8730
rect 18752 8676 18758 8678
rect 18814 8676 18838 8678
rect 18894 8676 18918 8678
rect 18974 8676 18998 8678
rect 19054 8676 19060 8678
rect 18752 8667 19060 8676
rect 18694 8528 18750 8537
rect 18604 8492 18656 8498
rect 18788 8492 18840 8498
rect 18750 8472 18788 8480
rect 18694 8463 18788 8472
rect 18708 8452 18788 8463
rect 18604 8434 18656 8440
rect 18788 8434 18840 8440
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18616 8022 18644 8230
rect 18708 8090 18736 8230
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18604 8016 18656 8022
rect 18604 7958 18656 7964
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18616 7002 18644 7822
rect 18752 7644 19060 7653
rect 18752 7642 18758 7644
rect 18814 7642 18838 7644
rect 18894 7642 18918 7644
rect 18974 7642 18998 7644
rect 19054 7642 19060 7644
rect 18814 7590 18816 7642
rect 18996 7590 18998 7642
rect 18752 7588 18758 7590
rect 18814 7588 18838 7590
rect 18894 7588 18918 7590
rect 18974 7588 18998 7590
rect 19054 7588 19060 7590
rect 18752 7579 19060 7588
rect 18788 7404 18840 7410
rect 18788 7346 18840 7352
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18800 6798 18828 7346
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 19168 5370 19196 6598
rect 19156 5364 19208 5370
rect 19156 5306 19208 5312
rect 18432 5222 18552 5250
rect 18788 5228 18840 5234
rect 18432 4264 18460 5222
rect 18788 5170 18840 5176
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 18800 4826 18828 5170
rect 19062 5128 19118 5137
rect 19062 5063 19118 5072
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 19076 4622 19104 5063
rect 19168 4826 19196 5170
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19260 4706 19288 11047
rect 19430 10840 19486 10849
rect 19430 10775 19432 10784
rect 19484 10775 19486 10784
rect 19432 10746 19484 10752
rect 19338 10704 19394 10713
rect 19338 10646 19340 10648
rect 19392 10646 19394 10648
rect 19338 10639 19394 10646
rect 19515 10668 19567 10674
rect 19515 10610 19567 10616
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 19536 10418 19564 10610
rect 19628 10418 19656 11290
rect 19706 10840 19762 10849
rect 19706 10775 19762 10784
rect 19352 10266 19380 10406
rect 19536 10390 19656 10418
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19536 9674 19564 10390
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19352 9646 19564 9674
rect 19352 8498 19380 9646
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19536 8498 19564 9318
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19536 7886 19564 8434
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 19352 6882 19380 7754
rect 19352 6854 19564 6882
rect 19536 6798 19564 6854
rect 19340 6792 19392 6798
rect 19524 6792 19576 6798
rect 19430 6760 19486 6769
rect 19392 6740 19430 6746
rect 19340 6734 19430 6740
rect 19352 6718 19430 6734
rect 19524 6734 19576 6740
rect 19430 6695 19486 6704
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5234 19380 5510
rect 19340 5228 19392 5234
rect 19340 5170 19392 5176
rect 19168 4678 19288 4706
rect 19352 4690 19380 5170
rect 19340 4684 19392 4690
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18512 4276 18564 4282
rect 18432 4236 18512 4264
rect 18616 4264 18644 4558
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18880 4276 18932 4282
rect 18616 4236 18828 4264
rect 18512 4218 18564 4224
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18326 4040 18382 4049
rect 18326 3975 18382 3984
rect 18234 3904 18290 3913
rect 18234 3839 18290 3848
rect 18144 3596 18196 3602
rect 18248 3584 18276 3839
rect 18196 3556 18276 3584
rect 18144 3538 18196 3544
rect 17972 3510 18092 3516
rect 17696 3454 17816 3482
rect 17960 3504 18092 3510
rect 17696 3194 17724 3454
rect 18012 3488 18092 3504
rect 18234 3496 18290 3505
rect 17960 3446 18012 3452
rect 18234 3431 18290 3440
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18142 3360 18198 3369
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17592 2984 17644 2990
rect 17236 2910 17448 2938
rect 17592 2926 17644 2932
rect 17144 2746 17356 2774
rect 17222 2680 17278 2689
rect 17040 2644 17092 2650
rect 17222 2615 17278 2624
rect 17040 2586 17092 2592
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 16764 2032 16816 2038
rect 16764 1974 16816 1980
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16672 1556 16724 1562
rect 16672 1498 16724 1504
rect 16396 1420 16448 1426
rect 16500 1414 16620 1442
rect 16396 1362 16448 1368
rect 16212 1284 16264 1290
rect 16212 1226 16264 1232
rect 16408 762 16436 1362
rect 16592 1358 16620 1414
rect 16488 1352 16540 1358
rect 16486 1320 16488 1329
rect 16580 1352 16632 1358
rect 16540 1320 16542 1329
rect 16580 1294 16632 1300
rect 16486 1255 16542 1264
rect 16684 1170 16712 1498
rect 16224 734 16436 762
rect 16500 1142 16712 1170
rect 16224 160 16252 734
rect 16500 160 16528 1142
rect 11242 82 11298 160
rect 11164 54 11298 82
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 12070 0 12126 160
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 0 14610 160
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 82 16818 160
rect 16868 82 16896 1702
rect 17052 160 17080 2586
rect 17236 2446 17264 2615
rect 17328 2514 17356 2746
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17224 2440 17276 2446
rect 17420 2428 17448 2910
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17512 2689 17540 2790
rect 17498 2680 17554 2689
rect 17498 2615 17554 2624
rect 17420 2400 17724 2428
rect 17224 2382 17276 2388
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17408 1760 17460 1766
rect 17408 1702 17460 1708
rect 16762 54 16896 82
rect 16762 0 16818 54
rect 17038 0 17094 160
rect 17314 82 17370 160
rect 17420 82 17448 1702
rect 17512 1358 17540 2246
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17500 1352 17552 1358
rect 17500 1294 17552 1300
rect 17604 160 17632 1702
rect 17696 1426 17724 2400
rect 17788 2038 17816 3334
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17880 2650 17908 2994
rect 17972 2961 18000 2994
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 17958 2680 18014 2689
rect 17868 2644 17920 2650
rect 17958 2615 18014 2624
rect 17868 2586 17920 2592
rect 17972 2514 18000 2615
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 2106 18000 2314
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17868 1488 17920 1494
rect 17868 1430 17920 1436
rect 17684 1420 17736 1426
rect 17684 1362 17736 1368
rect 17880 160 17908 1430
rect 18064 542 18092 3334
rect 18142 3295 18198 3304
rect 18156 2417 18184 3295
rect 18248 3058 18276 3431
rect 18340 3194 18368 3975
rect 18708 3777 18736 4082
rect 18694 3768 18750 3777
rect 18800 3738 18828 4236
rect 19168 4264 19196 4678
rect 19340 4626 19392 4632
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19260 4282 19288 4558
rect 18880 4218 18932 4224
rect 19076 4236 19196 4264
rect 19248 4276 19300 4282
rect 18694 3703 18750 3712
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18788 3528 18840 3534
rect 18423 3488 18736 3516
rect 18423 3380 18451 3488
rect 18708 3398 18736 3488
rect 18892 3516 18920 4218
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 4010 19012 4082
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 19076 3534 19104 4236
rect 19444 4264 19472 6598
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19248 4218 19300 4224
rect 19352 4236 19472 4264
rect 19536 5148 19564 5850
rect 19628 5284 19656 10202
rect 19720 9518 19748 10775
rect 19708 9512 19760 9518
rect 19708 9454 19760 9460
rect 19720 7478 19748 9454
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 19708 5296 19760 5302
rect 19628 5256 19708 5284
rect 19708 5238 19760 5244
rect 19616 5160 19668 5166
rect 19536 5120 19616 5148
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19168 3777 19196 3878
rect 19154 3768 19210 3777
rect 19154 3703 19210 3712
rect 19156 3664 19208 3670
rect 19156 3606 19208 3612
rect 18840 3488 18920 3516
rect 19064 3528 19116 3534
rect 18788 3470 18840 3476
rect 19064 3470 19116 3476
rect 18604 3392 18656 3398
rect 18423 3352 18460 3380
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18142 2408 18198 2417
rect 18142 2343 18198 2352
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 18052 536 18104 542
rect 18052 478 18104 484
rect 17314 54 17448 82
rect 17314 0 17370 54
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 82 18198 160
rect 18248 82 18276 2246
rect 18340 1358 18368 2790
rect 18432 2446 18460 3352
rect 18602 3360 18604 3369
rect 18696 3392 18748 3398
rect 18656 3360 18658 3369
rect 18696 3334 18748 3340
rect 18602 3295 18658 3304
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 19168 3233 19196 3606
rect 19154 3224 19210 3233
rect 19064 3188 19116 3194
rect 19154 3159 19210 3168
rect 19064 3130 19116 3136
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18696 3052 18748 3058
rect 18880 3052 18932 3058
rect 18748 3012 18828 3040
rect 18696 2994 18748 3000
rect 18694 2952 18750 2961
rect 18694 2887 18696 2896
rect 18748 2887 18750 2896
rect 18696 2858 18748 2864
rect 18510 2680 18566 2689
rect 18510 2615 18566 2624
rect 18694 2680 18750 2689
rect 18800 2666 18828 3012
rect 18880 2994 18932 3000
rect 18750 2638 18828 2666
rect 18694 2615 18750 2624
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 18432 160 18460 2246
rect 18524 1970 18552 2615
rect 18892 2582 18920 2994
rect 18984 2854 19012 3062
rect 18972 2848 19024 2854
rect 18972 2790 19024 2796
rect 18880 2576 18932 2582
rect 18880 2518 18932 2524
rect 18604 2440 18656 2446
rect 18602 2408 18604 2417
rect 18656 2408 18658 2417
rect 18602 2343 18658 2352
rect 19076 2292 19104 3130
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 18616 2264 19104 2292
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18616 1000 18644 2264
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 18616 972 18736 1000
rect 18708 160 18736 972
rect 18142 54 18276 82
rect 18142 0 18198 54
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 82 19026 160
rect 19168 82 19196 2790
rect 19260 2394 19288 3878
rect 19352 3466 19380 4236
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19340 3460 19392 3466
rect 19444 3448 19472 4082
rect 19536 4049 19564 5120
rect 19616 5102 19668 5108
rect 19616 5024 19668 5030
rect 19616 4966 19668 4972
rect 19628 4826 19656 4966
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19812 4622 19840 12406
rect 19904 12322 19932 15438
rect 19996 15026 20024 15846
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 20088 12434 20116 21134
rect 20260 21004 20312 21010
rect 20312 20964 20392 20992
rect 20260 20946 20312 20952
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18970 20300 19110
rect 20260 18964 20312 18970
rect 20260 18906 20312 18912
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16794 20208 16934
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20168 15904 20220 15910
rect 20168 15846 20220 15852
rect 20180 15502 20208 15846
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20260 14884 20312 14890
rect 20260 14826 20312 14832
rect 20272 14618 20300 14826
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20364 13410 20392 20964
rect 20640 20924 20668 22052
rect 20812 22024 20864 22030
rect 20812 21966 20864 21972
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21078 20760 21898
rect 20824 21690 20852 21966
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20916 20942 20944 21830
rect 21008 21690 21036 21830
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 20904 20936 20956 20942
rect 20640 20896 20760 20924
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20536 19236 20588 19242
rect 20536 19178 20588 19184
rect 20548 17626 20576 19178
rect 20640 18766 20668 19654
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20732 18057 20760 20896
rect 20904 20878 20956 20884
rect 20812 19712 20864 19718
rect 20812 19654 20864 19660
rect 20824 19514 20852 19654
rect 21100 19530 21128 24126
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 21008 19502 21128 19530
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20718 18048 20774 18057
rect 20718 17983 20774 17992
rect 20548 17598 20760 17626
rect 20548 17134 20576 17598
rect 20732 17542 20760 17598
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20640 17338 20668 17478
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20536 17128 20588 17134
rect 20536 17070 20588 17076
rect 20456 16674 20484 17070
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20456 16658 20576 16674
rect 20456 16652 20588 16658
rect 20456 16646 20536 16652
rect 20536 16594 20588 16600
rect 20732 16250 20760 16934
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20626 15056 20682 15065
rect 20626 14991 20682 15000
rect 20812 15020 20864 15026
rect 20444 13796 20496 13802
rect 20444 13738 20496 13744
rect 20456 13530 20484 13738
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20364 13382 20484 13410
rect 20352 13320 20404 13326
rect 20352 13262 20404 13268
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20180 12986 20208 13194
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20364 12646 20392 13262
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20456 12434 20484 13382
rect 20088 12406 20392 12434
rect 20456 12406 20576 12434
rect 20364 12322 20392 12406
rect 19904 12294 20208 12322
rect 20364 12294 20484 12322
rect 20180 12238 20208 12294
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 19904 9926 19932 11086
rect 20088 10810 20116 11086
rect 20076 10804 20128 10810
rect 20076 10746 20128 10752
rect 20272 10266 20300 11086
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20168 8492 20220 8498
rect 20168 8434 20220 8440
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19904 7546 19932 7822
rect 19996 7818 20024 8230
rect 20180 8090 20208 8434
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20076 8016 20128 8022
rect 20076 7958 20128 7964
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 20088 6780 20116 7958
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 19904 6752 20116 6780
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19522 4040 19578 4049
rect 19522 3975 19578 3984
rect 19524 3460 19576 3466
rect 19444 3420 19524 3448
rect 19340 3402 19392 3408
rect 19524 3402 19576 3408
rect 19536 3194 19564 3402
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19430 2680 19486 2689
rect 19430 2615 19486 2624
rect 19444 2446 19472 2615
rect 19628 2582 19656 2926
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 19432 2440 19484 2446
rect 19260 2366 19380 2394
rect 19432 2382 19484 2388
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19260 2106 19288 2246
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19352 1986 19380 2366
rect 19536 2106 19564 2382
rect 19524 2100 19576 2106
rect 19524 2042 19576 2048
rect 19260 1958 19380 1986
rect 19260 160 19288 1958
rect 19432 1896 19484 1902
rect 19432 1838 19484 1844
rect 19444 1562 19472 1838
rect 19720 1714 19748 3334
rect 19812 3058 19840 4422
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19904 2990 19932 6752
rect 20180 5778 20208 7278
rect 20168 5772 20220 5778
rect 20168 5714 20220 5720
rect 20272 5409 20300 8774
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 20364 7002 20392 7822
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20258 5400 20314 5409
rect 20258 5335 20314 5344
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20088 4622 20116 4966
rect 20364 4826 20392 5646
rect 20352 4820 20404 4826
rect 20352 4762 20404 4768
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 4282 20300 4422
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20364 4146 20392 4762
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20076 4072 20128 4078
rect 20456 4026 20484 12294
rect 20548 6798 20576 12406
rect 20640 10690 20668 14991
rect 20812 14962 20864 14968
rect 20824 14074 20852 14962
rect 20916 14929 20944 18566
rect 21008 18290 21036 19502
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21100 18970 21128 19314
rect 21192 19242 21220 24006
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21284 21026 21312 22918
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21468 22166 21496 22578
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 21560 21690 21588 24262
rect 21652 22094 21680 26998
rect 21719 26684 22027 26693
rect 21719 26682 21725 26684
rect 21781 26682 21805 26684
rect 21861 26682 21885 26684
rect 21941 26682 21965 26684
rect 22021 26682 22027 26684
rect 21781 26630 21783 26682
rect 21963 26630 21965 26682
rect 21719 26628 21725 26630
rect 21781 26628 21805 26630
rect 21861 26628 21885 26630
rect 21941 26628 21965 26630
rect 22021 26628 22027 26630
rect 21719 26619 22027 26628
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21719 25596 22027 25605
rect 21719 25594 21725 25596
rect 21781 25594 21805 25596
rect 21861 25594 21885 25596
rect 21941 25594 21965 25596
rect 22021 25594 22027 25596
rect 21781 25542 21783 25594
rect 21963 25542 21965 25594
rect 21719 25540 21725 25542
rect 21781 25540 21805 25542
rect 21861 25540 21885 25542
rect 21941 25540 21965 25542
rect 22021 25540 22027 25542
rect 21719 25531 22027 25540
rect 22112 25226 22140 25842
rect 21732 25220 21784 25226
rect 21732 25162 21784 25168
rect 22100 25220 22152 25226
rect 22100 25162 22152 25168
rect 21744 24857 21772 25162
rect 21730 24848 21786 24857
rect 21730 24783 21786 24792
rect 22192 24744 22244 24750
rect 22192 24686 22244 24692
rect 21719 24508 22027 24517
rect 21719 24506 21725 24508
rect 21781 24506 21805 24508
rect 21861 24506 21885 24508
rect 21941 24506 21965 24508
rect 22021 24506 22027 24508
rect 21781 24454 21783 24506
rect 21963 24454 21965 24506
rect 21719 24452 21725 24454
rect 21781 24452 21805 24454
rect 21861 24452 21885 24454
rect 21941 24452 21965 24454
rect 22021 24452 22027 24454
rect 21719 24443 22027 24452
rect 21719 23420 22027 23429
rect 21719 23418 21725 23420
rect 21781 23418 21805 23420
rect 21861 23418 21885 23420
rect 21941 23418 21965 23420
rect 22021 23418 22027 23420
rect 21781 23366 21783 23418
rect 21963 23366 21965 23418
rect 21719 23364 21725 23366
rect 21781 23364 21805 23366
rect 21861 23364 21885 23366
rect 21941 23364 21965 23366
rect 22021 23364 22027 23366
rect 21719 23355 22027 23364
rect 21732 23112 21784 23118
rect 22204 23066 22232 24686
rect 21732 23054 21784 23060
rect 21744 22778 21772 23054
rect 22020 23038 22232 23066
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 22020 22642 22048 23038
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 21744 22545 21772 22578
rect 21730 22536 21786 22545
rect 21730 22471 21786 22480
rect 21719 22332 22027 22341
rect 21719 22330 21725 22332
rect 21781 22330 21805 22332
rect 21861 22330 21885 22332
rect 21941 22330 21965 22332
rect 22021 22330 22027 22332
rect 21781 22278 21783 22330
rect 21963 22278 21965 22330
rect 21719 22276 21725 22278
rect 21781 22276 21805 22278
rect 21861 22276 21885 22278
rect 21941 22276 21965 22278
rect 22021 22276 22027 22278
rect 21719 22267 22027 22276
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 21652 22066 21772 22094
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21364 21344 21416 21350
rect 21364 21286 21416 21292
rect 21376 21146 21404 21286
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21284 20998 21404 21026
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21284 19378 21312 19790
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 21180 19236 21232 19242
rect 21180 19178 21232 19184
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 21376 18426 21404 20998
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21284 17678 21312 18158
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21088 17264 21140 17270
rect 21468 17218 21496 21490
rect 21744 21434 21772 22066
rect 21652 21406 21772 21434
rect 21546 19952 21602 19961
rect 21546 19887 21602 19896
rect 21560 19854 21588 19887
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21560 17513 21588 19790
rect 21652 18329 21680 21406
rect 22020 21332 22048 22170
rect 22112 22030 22140 22918
rect 22204 22234 22232 22918
rect 22296 22710 22324 28966
rect 22388 24970 22416 33487
rect 22572 33425 22600 33934
rect 22652 33856 22704 33862
rect 22652 33798 22704 33804
rect 22664 33658 22692 33798
rect 22848 33658 22876 33934
rect 22652 33652 22704 33658
rect 22652 33594 22704 33600
rect 22836 33652 22888 33658
rect 22836 33594 22888 33600
rect 22558 33416 22614 33425
rect 22558 33351 22614 33360
rect 22652 32972 22704 32978
rect 22652 32914 22704 32920
rect 22560 30592 22612 30598
rect 22560 30534 22612 30540
rect 22572 29646 22600 30534
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22560 27940 22612 27946
rect 22560 27882 22612 27888
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22480 27674 22508 27814
rect 22468 27668 22520 27674
rect 22468 27610 22520 27616
rect 22572 25294 22600 27882
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22560 25152 22612 25158
rect 22560 25094 22612 25100
rect 22388 24942 22508 24970
rect 22376 24812 22428 24818
rect 22376 24754 22428 24760
rect 22388 24410 22416 24754
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22480 24206 22508 24942
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22572 23866 22600 25094
rect 22664 24410 22692 32914
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 22756 28966 22784 30194
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22848 29850 22876 29990
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22744 28960 22796 28966
rect 22744 28902 22796 28908
rect 22756 25752 22784 28902
rect 22940 28150 22968 37742
rect 23032 37398 23060 38218
rect 23124 37466 23152 38354
rect 23492 38350 23520 38762
rect 23584 38554 23612 38898
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 23480 38344 23532 38350
rect 23480 38286 23532 38292
rect 23112 37460 23164 37466
rect 23112 37402 23164 37408
rect 23020 37392 23072 37398
rect 23020 37334 23072 37340
rect 23676 37262 23704 38898
rect 23768 38554 23796 39986
rect 23940 39840 23992 39846
rect 23940 39782 23992 39788
rect 23952 39438 23980 39782
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23940 39432 23992 39438
rect 23940 39374 23992 39380
rect 23860 39098 23888 39374
rect 23940 39296 23992 39302
rect 23940 39238 23992 39244
rect 23848 39092 23900 39098
rect 23848 39034 23900 39040
rect 23756 38548 23808 38554
rect 23756 38490 23808 38496
rect 23952 38350 23980 39238
rect 24044 38962 24072 39986
rect 24032 38956 24084 38962
rect 24032 38898 24084 38904
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 24136 38026 24164 40174
rect 23952 37998 24164 38026
rect 23952 37262 23980 37998
rect 24032 37868 24084 37874
rect 24032 37810 24084 37816
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23664 37256 23716 37262
rect 23664 37198 23716 37204
rect 23940 37256 23992 37262
rect 23940 37198 23992 37204
rect 23020 36780 23072 36786
rect 23020 36722 23072 36728
rect 23032 35834 23060 36722
rect 23584 36378 23612 37198
rect 23848 37188 23900 37194
rect 23848 37130 23900 37136
rect 23860 36922 23888 37130
rect 24044 36922 24072 37810
rect 24124 37324 24176 37330
rect 24124 37266 24176 37272
rect 24136 37233 24164 37266
rect 24122 37224 24178 37233
rect 24122 37159 24178 37168
rect 23848 36916 23900 36922
rect 23848 36858 23900 36864
rect 24032 36916 24084 36922
rect 24032 36858 24084 36864
rect 24032 36780 24084 36786
rect 24032 36722 24084 36728
rect 23572 36372 23624 36378
rect 23572 36314 23624 36320
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23584 35834 23612 36110
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23572 35828 23624 35834
rect 23572 35770 23624 35776
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 23112 34400 23164 34406
rect 23112 34342 23164 34348
rect 23124 33522 23152 34342
rect 23112 33516 23164 33522
rect 23112 33458 23164 33464
rect 23216 31754 23244 35634
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23388 35080 23440 35086
rect 23388 35022 23440 35028
rect 23400 34202 23428 35022
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23388 34196 23440 34202
rect 23388 34138 23440 34144
rect 23492 33998 23520 34886
rect 23676 34746 23704 35226
rect 23768 34746 23796 35430
rect 23664 34740 23716 34746
rect 23664 34682 23716 34688
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 23952 34678 23980 35634
rect 23940 34672 23992 34678
rect 23940 34614 23992 34620
rect 23756 34604 23808 34610
rect 23756 34546 23808 34552
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23480 33856 23532 33862
rect 23308 33816 23480 33844
rect 23308 32842 23336 33816
rect 23480 33798 23532 33804
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33658 23704 33798
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23388 33312 23440 33318
rect 23388 33254 23440 33260
rect 23480 33312 23532 33318
rect 23480 33254 23532 33260
rect 23400 33114 23428 33254
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23296 32836 23348 32842
rect 23296 32778 23348 32784
rect 23492 32586 23520 33254
rect 23768 32910 23796 34546
rect 23756 32904 23808 32910
rect 23756 32846 23808 32852
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 23492 32558 23704 32586
rect 23952 32570 23980 32846
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23124 31726 23244 31754
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 22836 28076 22888 28082
rect 22836 28018 22888 28024
rect 22848 27674 22876 28018
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23032 27674 23060 27814
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 23020 27668 23072 27674
rect 23020 27610 23072 27616
rect 22836 27396 22888 27402
rect 22836 27338 22888 27344
rect 22848 27130 22876 27338
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 22836 27124 22888 27130
rect 22836 27066 22888 27072
rect 22940 26790 22968 27270
rect 23032 27130 23060 27270
rect 23020 27124 23072 27130
rect 23020 27066 23072 27072
rect 23124 27010 23152 31726
rect 23296 31408 23348 31414
rect 23296 31350 23348 31356
rect 23308 30734 23336 31350
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 23204 30048 23256 30054
rect 23204 29990 23256 29996
rect 23216 29850 23244 29990
rect 23204 29844 23256 29850
rect 23204 29786 23256 29792
rect 23032 26994 23152 27010
rect 23020 26988 23152 26994
rect 23072 26982 23152 26988
rect 23020 26930 23072 26936
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 22756 25724 23060 25752
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22664 23118 22692 23666
rect 22376 23112 22428 23118
rect 22376 23054 22428 23060
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22284 22704 22336 22710
rect 22284 22646 22336 22652
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22192 22228 22244 22234
rect 22192 22170 22244 22176
rect 22296 22098 22324 22374
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21690 22324 21830
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22190 21448 22246 21457
rect 22190 21383 22246 21392
rect 22020 21304 22140 21332
rect 21719 21244 22027 21253
rect 21719 21242 21725 21244
rect 21781 21242 21805 21244
rect 21861 21242 21885 21244
rect 21941 21242 21965 21244
rect 22021 21242 22027 21244
rect 21781 21190 21783 21242
rect 21963 21190 21965 21242
rect 21719 21188 21725 21190
rect 21781 21188 21805 21190
rect 21861 21188 21885 21190
rect 21941 21188 21965 21190
rect 22021 21188 22027 21190
rect 21719 21179 22027 21188
rect 22112 20942 22140 21304
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22112 20602 22140 20878
rect 22100 20596 22152 20602
rect 22100 20538 22152 20544
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21719 20156 22027 20165
rect 21719 20154 21725 20156
rect 21781 20154 21805 20156
rect 21861 20154 21885 20156
rect 21941 20154 21965 20156
rect 22021 20154 22027 20156
rect 21781 20102 21783 20154
rect 21963 20102 21965 20154
rect 21719 20100 21725 20102
rect 21781 20100 21805 20102
rect 21861 20100 21885 20102
rect 21941 20100 21965 20102
rect 22021 20100 22027 20102
rect 21719 20091 22027 20100
rect 22112 20058 22140 20402
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21719 19068 22027 19077
rect 21719 19066 21725 19068
rect 21781 19066 21805 19068
rect 21861 19066 21885 19068
rect 21941 19066 21965 19068
rect 22021 19066 22027 19068
rect 21781 19014 21783 19066
rect 21963 19014 21965 19066
rect 21719 19012 21725 19014
rect 21781 19012 21805 19014
rect 21861 19012 21885 19014
rect 21941 19012 21965 19014
rect 22021 19012 22027 19014
rect 21719 19003 22027 19012
rect 21638 18320 21694 18329
rect 21638 18255 21694 18264
rect 21719 17980 22027 17989
rect 21719 17978 21725 17980
rect 21781 17978 21805 17980
rect 21861 17978 21885 17980
rect 21941 17978 21965 17980
rect 22021 17978 22027 17980
rect 21781 17926 21783 17978
rect 21963 17926 21965 17978
rect 21719 17924 21725 17926
rect 21781 17924 21805 17926
rect 21861 17924 21885 17926
rect 21941 17924 21965 17926
rect 22021 17924 22027 17926
rect 21719 17915 22027 17924
rect 22204 17762 22232 21383
rect 22388 21010 22416 23054
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22466 22536 22522 22545
rect 22466 22471 22522 22480
rect 22480 22166 22508 22471
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22282 19952 22338 19961
rect 22282 19887 22338 19896
rect 22296 17785 22324 19887
rect 22388 18222 22416 20946
rect 22572 20466 22600 22578
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22848 22234 22876 22374
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22652 20868 22704 20874
rect 22652 20810 22704 20816
rect 22664 20482 22692 20810
rect 22836 20528 22888 20534
rect 22664 20476 22836 20482
rect 22664 20470 22888 20476
rect 22560 20460 22612 20466
rect 22664 20454 22876 20470
rect 22560 20402 22612 20408
rect 22572 20058 22600 20402
rect 22652 20324 22704 20330
rect 22652 20266 22704 20272
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22376 18216 22428 18222
rect 22376 18158 22428 18164
rect 22572 17882 22600 19994
rect 22664 19378 22692 20266
rect 22756 19825 22784 20454
rect 22742 19816 22798 19825
rect 22742 19751 22798 19760
rect 23032 19700 23060 25724
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23124 25498 23152 25638
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 23308 24290 23336 30534
rect 23492 26874 23520 31758
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30394 23612 30534
rect 23572 30388 23624 30394
rect 23572 30330 23624 30336
rect 23572 27532 23624 27538
rect 23572 27474 23624 27480
rect 23584 27130 23612 27474
rect 23572 27124 23624 27130
rect 23572 27066 23624 27072
rect 23492 26846 23612 26874
rect 23584 26518 23612 26846
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23676 26466 23704 32558
rect 23940 32564 23992 32570
rect 23940 32506 23992 32512
rect 24044 32230 24072 36722
rect 24228 36650 24256 42026
rect 24400 39840 24452 39846
rect 24398 39808 24400 39817
rect 24452 39808 24454 39817
rect 24398 39743 24454 39752
rect 24400 38752 24452 38758
rect 24398 38720 24400 38729
rect 24452 38720 24454 38729
rect 24398 38655 24454 38664
rect 24400 37664 24452 37670
rect 24398 37632 24400 37641
rect 24452 37632 24454 37641
rect 24398 37567 24454 37576
rect 24216 36644 24268 36650
rect 24216 36586 24268 36592
rect 24400 36576 24452 36582
rect 24398 36544 24400 36553
rect 24452 36544 24454 36553
rect 24398 36479 24454 36488
rect 24400 35488 24452 35494
rect 24398 35456 24400 35465
rect 24452 35456 24454 35465
rect 24398 35391 24454 35400
rect 24400 34536 24452 34542
rect 24398 34504 24400 34513
rect 24452 34504 24454 34513
rect 24398 34439 24454 34448
rect 24400 33312 24452 33318
rect 24398 33280 24400 33289
rect 24452 33280 24454 33289
rect 24398 33215 24454 33224
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 24136 32026 24164 32370
rect 24400 32224 24452 32230
rect 24398 32192 24400 32201
rect 24452 32192 24454 32201
rect 24398 32127 24454 32136
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 23756 31952 23808 31958
rect 23756 31894 23808 31900
rect 23768 27962 23796 31894
rect 24308 31680 24360 31686
rect 24308 31622 24360 31628
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23860 30394 23888 31282
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 30394 23980 31078
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 24216 29572 24268 29578
rect 24216 29514 24268 29520
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23768 27934 23888 27962
rect 23756 27872 23808 27878
rect 23756 27814 23808 27820
rect 23768 27130 23796 27814
rect 23756 27124 23808 27130
rect 23756 27066 23808 27072
rect 23756 26988 23808 26994
rect 23756 26930 23808 26936
rect 23768 26586 23796 26930
rect 23756 26580 23808 26586
rect 23756 26522 23808 26528
rect 23676 26438 23796 26466
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23400 24410 23428 25774
rect 23492 25362 23520 26318
rect 23584 26042 23612 26318
rect 23664 26240 23716 26246
rect 23664 26182 23716 26188
rect 23572 26036 23624 26042
rect 23572 25978 23624 25984
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23584 25498 23612 25842
rect 23676 25498 23704 26182
rect 23768 25786 23796 26438
rect 23860 25974 23888 27934
rect 23952 27674 23980 28018
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 24124 26784 24176 26790
rect 24124 26726 24176 26732
rect 23848 25968 23900 25974
rect 23848 25910 23900 25916
rect 23768 25758 23888 25786
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23664 25492 23716 25498
rect 23664 25434 23716 25440
rect 23480 25356 23532 25362
rect 23480 25298 23532 25304
rect 23492 24954 23520 25298
rect 23756 25152 23808 25158
rect 23756 25094 23808 25100
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23388 24404 23440 24410
rect 23388 24346 23440 24352
rect 23308 24262 23520 24290
rect 23296 24200 23348 24206
rect 23296 24142 23348 24148
rect 23308 23866 23336 24142
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 23216 22778 23244 23666
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23216 22094 23244 22714
rect 23124 22066 23244 22094
rect 23308 22094 23336 23462
rect 23492 22982 23520 24262
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23584 23633 23612 24142
rect 23570 23624 23626 23633
rect 23570 23559 23626 23568
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23388 22094 23440 22098
rect 23308 22092 23440 22094
rect 23308 22066 23388 22092
rect 23124 22030 23152 22066
rect 23388 22034 23440 22040
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23492 21962 23520 22578
rect 23584 22234 23612 23462
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 23676 22094 23704 24142
rect 23768 23118 23796 25094
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23860 22930 23888 25758
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23952 23322 23980 23666
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 24032 22976 24084 22982
rect 23860 22902 23980 22930
rect 24032 22918 24084 22924
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23676 22066 23796 22094
rect 23768 22030 23796 22066
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23480 21956 23532 21962
rect 23480 21898 23532 21904
rect 23388 21888 23440 21894
rect 23860 21842 23888 22646
rect 23388 21830 23440 21836
rect 23112 21480 23164 21486
rect 23112 21422 23164 21428
rect 22756 19672 23060 19700
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22112 17734 22232 17762
rect 22282 17776 22338 17785
rect 21640 17536 21692 17542
rect 21546 17504 21602 17513
rect 21640 17478 21692 17484
rect 21546 17439 21602 17448
rect 21088 17206 21140 17212
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16114 21036 16390
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20902 14920 20958 14929
rect 20902 14855 20958 14864
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20916 13938 20944 14855
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 21008 13818 21036 15914
rect 20916 13790 21036 13818
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20824 12986 20852 13262
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20812 12164 20864 12170
rect 20812 12106 20864 12112
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10810 20760 11086
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20824 10713 20852 12106
rect 20810 10704 20866 10713
rect 20640 10674 20760 10690
rect 20640 10668 20772 10674
rect 20640 10662 20720 10668
rect 20810 10639 20866 10648
rect 20720 10610 20772 10616
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20640 9654 20668 9862
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20640 8430 20668 9590
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20640 7546 20668 7822
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20628 6928 20680 6934
rect 20732 6905 20760 10610
rect 20824 10130 20852 10639
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20810 9888 20866 9897
rect 20810 9823 20866 9832
rect 20824 7750 20852 9823
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20916 7562 20944 13790
rect 21100 11354 21128 17206
rect 21376 17190 21496 17218
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21192 15094 21220 15438
rect 21180 15088 21232 15094
rect 21180 15030 21232 15036
rect 21192 13326 21220 15030
rect 21284 14958 21312 16594
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21192 12918 21220 13262
rect 21180 12912 21232 12918
rect 21180 12854 21232 12860
rect 21192 12628 21220 12854
rect 21284 12753 21312 13670
rect 21270 12744 21326 12753
rect 21270 12679 21326 12688
rect 21192 12600 21312 12628
rect 21178 12336 21234 12345
rect 21178 12271 21234 12280
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21100 9722 21128 10610
rect 21192 10062 21220 12271
rect 21284 12238 21312 12600
rect 21376 12434 21404 17190
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21468 16794 21496 17002
rect 21548 16992 21600 16998
rect 21548 16934 21600 16940
rect 21560 16794 21588 16934
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21652 16726 21680 17478
rect 22112 17218 22140 17734
rect 22282 17711 22338 17720
rect 22192 17672 22244 17678
rect 22192 17614 22244 17620
rect 22204 17338 22232 17614
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17338 22508 17478
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22112 17190 22232 17218
rect 21824 17128 21876 17134
rect 21876 17076 22140 17082
rect 21824 17070 22140 17076
rect 21836 17054 22140 17070
rect 21719 16892 22027 16901
rect 21719 16890 21725 16892
rect 21781 16890 21805 16892
rect 21861 16890 21885 16892
rect 21941 16890 21965 16892
rect 22021 16890 22027 16892
rect 21781 16838 21783 16890
rect 21963 16838 21965 16890
rect 21719 16836 21725 16838
rect 21781 16836 21805 16838
rect 21861 16836 21885 16838
rect 21941 16836 21965 16838
rect 22021 16836 22027 16838
rect 21719 16827 22027 16836
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21468 16250 21496 16594
rect 22112 16454 22140 17054
rect 21640 16448 21692 16454
rect 21640 16390 21692 16396
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21456 16244 21508 16250
rect 21456 16186 21508 16192
rect 21652 15638 21680 16390
rect 21719 15804 22027 15813
rect 21719 15802 21725 15804
rect 21781 15802 21805 15804
rect 21861 15802 21885 15804
rect 21941 15802 21965 15804
rect 22021 15802 22027 15804
rect 21781 15750 21783 15802
rect 21963 15750 21965 15802
rect 21719 15748 21725 15750
rect 21781 15748 21805 15750
rect 21861 15748 21885 15750
rect 21941 15748 21965 15750
rect 22021 15748 22027 15750
rect 21719 15739 22027 15748
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21468 12646 21496 13126
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21560 12442 21588 14894
rect 21719 14716 22027 14725
rect 21719 14714 21725 14716
rect 21781 14714 21805 14716
rect 21861 14714 21885 14716
rect 21941 14714 21965 14716
rect 22021 14714 22027 14716
rect 21781 14662 21783 14714
rect 21963 14662 21965 14714
rect 21719 14660 21725 14662
rect 21781 14660 21805 14662
rect 21861 14660 21885 14662
rect 21941 14660 21965 14662
rect 22021 14660 22027 14662
rect 21719 14651 22027 14660
rect 21640 14272 21692 14278
rect 21640 14214 21692 14220
rect 21548 12436 21600 12442
rect 21376 12406 21496 12434
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21008 8090 21036 9658
rect 21192 8906 21220 9862
rect 21284 8974 21312 12174
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21376 8276 21404 11018
rect 21468 10146 21496 12406
rect 21652 12434 21680 14214
rect 21719 13628 22027 13637
rect 21719 13626 21725 13628
rect 21781 13626 21805 13628
rect 21861 13626 21885 13628
rect 21941 13626 21965 13628
rect 22021 13626 22027 13628
rect 21781 13574 21783 13626
rect 21963 13574 21965 13626
rect 21719 13572 21725 13574
rect 21781 13572 21805 13574
rect 21861 13572 21885 13574
rect 21941 13572 21965 13574
rect 22021 13572 22027 13574
rect 21719 13563 22027 13572
rect 22112 12866 22140 16390
rect 22204 15502 22232 17190
rect 22572 16454 22600 17818
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22572 16046 22600 16390
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22756 15722 22784 19672
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22848 17202 22876 19450
rect 23124 19378 23152 21422
rect 23296 20800 23348 20806
rect 23296 20742 23348 20748
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23216 19514 23244 19654
rect 23308 19514 23336 20742
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23112 19236 23164 19242
rect 23112 19178 23164 19184
rect 23124 19122 23152 19178
rect 23124 19094 23244 19122
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22836 17196 22888 17202
rect 22836 17138 22888 17144
rect 22940 16590 22968 18702
rect 23020 18624 23072 18630
rect 23020 18566 23072 18572
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 23032 17338 23060 18566
rect 23124 18358 23152 18566
rect 23112 18352 23164 18358
rect 23112 18294 23164 18300
rect 23216 17542 23244 19094
rect 23400 18766 23428 21830
rect 23676 21814 23888 21842
rect 23676 21554 23704 21814
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23492 21434 23520 21490
rect 23492 21406 23612 21434
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 20398 23520 21286
rect 23584 20602 23612 21406
rect 23664 21412 23716 21418
rect 23664 21354 23716 21360
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23480 20392 23532 20398
rect 23480 20334 23532 20340
rect 23676 19854 23704 21354
rect 23848 21344 23900 21350
rect 23846 21312 23848 21321
rect 23900 21312 23902 21321
rect 23846 21247 23902 21256
rect 23664 19848 23716 19854
rect 23664 19790 23716 19796
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23860 19258 23888 19722
rect 23952 19446 23980 22902
rect 24044 22098 24072 22918
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24032 20936 24084 20942
rect 24032 20878 24084 20884
rect 24044 20330 24072 20878
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 24030 20224 24086 20233
rect 24030 20159 24086 20168
rect 24044 20058 24072 20159
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24136 19446 24164 26726
rect 24228 24818 24256 29514
rect 24320 26042 24348 31622
rect 24400 31136 24452 31142
rect 24398 31104 24400 31113
rect 24452 31104 24454 31113
rect 24398 31039 24454 31048
rect 24504 30818 24532 42214
rect 24596 35290 24624 42230
rect 24686 41372 24994 41381
rect 24686 41370 24692 41372
rect 24748 41370 24772 41372
rect 24828 41370 24852 41372
rect 24908 41370 24932 41372
rect 24988 41370 24994 41372
rect 24748 41318 24750 41370
rect 24930 41318 24932 41370
rect 24686 41316 24692 41318
rect 24748 41316 24772 41318
rect 24828 41316 24852 41318
rect 24908 41316 24932 41318
rect 24988 41316 24994 41318
rect 24686 41307 24994 41316
rect 25056 41274 25084 44463
rect 25332 43160 25360 44463
rect 25332 43132 25452 43160
rect 25318 43072 25374 43081
rect 25318 43007 25374 43016
rect 25136 42764 25188 42770
rect 25136 42706 25188 42712
rect 25148 42537 25176 42706
rect 25134 42528 25190 42537
rect 25134 42463 25190 42472
rect 25228 42016 25280 42022
rect 25228 41958 25280 41964
rect 25240 41449 25268 41958
rect 25332 41818 25360 43007
rect 25424 41818 25452 43132
rect 25608 42158 25636 44463
rect 25596 42152 25648 42158
rect 25596 42094 25648 42100
rect 25320 41812 25372 41818
rect 25320 41754 25372 41760
rect 25412 41812 25464 41818
rect 25412 41754 25464 41760
rect 25780 41608 25832 41614
rect 25780 41550 25832 41556
rect 25226 41440 25282 41449
rect 25226 41375 25282 41384
rect 25044 41268 25096 41274
rect 25044 41210 25096 41216
rect 25320 40656 25372 40662
rect 25320 40598 25372 40604
rect 25136 40452 25188 40458
rect 25136 40394 25188 40400
rect 25148 40361 25176 40394
rect 25134 40352 25190 40361
rect 24686 40284 24994 40293
rect 25134 40287 25190 40296
rect 24686 40282 24692 40284
rect 24748 40282 24772 40284
rect 24828 40282 24852 40284
rect 24908 40282 24932 40284
rect 24988 40282 24994 40284
rect 24748 40230 24750 40282
rect 24930 40230 24932 40282
rect 24686 40228 24692 40230
rect 24748 40228 24772 40230
rect 24828 40228 24852 40230
rect 24908 40228 24932 40230
rect 24988 40228 24994 40230
rect 24686 40219 24994 40228
rect 25228 39296 25280 39302
rect 25226 39264 25228 39273
rect 25280 39264 25282 39273
rect 24686 39196 24994 39205
rect 25226 39199 25282 39208
rect 24686 39194 24692 39196
rect 24748 39194 24772 39196
rect 24828 39194 24852 39196
rect 24908 39194 24932 39196
rect 24988 39194 24994 39196
rect 24748 39142 24750 39194
rect 24930 39142 24932 39194
rect 24686 39140 24692 39142
rect 24748 39140 24772 39142
rect 24828 39140 24852 39142
rect 24908 39140 24932 39142
rect 24988 39140 24994 39142
rect 24686 39131 24994 39140
rect 25228 38208 25280 38214
rect 25226 38176 25228 38185
rect 25280 38176 25282 38185
rect 24686 38108 24994 38117
rect 25226 38111 25282 38120
rect 24686 38106 24692 38108
rect 24748 38106 24772 38108
rect 24828 38106 24852 38108
rect 24908 38106 24932 38108
rect 24988 38106 24994 38108
rect 24748 38054 24750 38106
rect 24930 38054 24932 38106
rect 24686 38052 24692 38054
rect 24748 38052 24772 38054
rect 24828 38052 24852 38054
rect 24908 38052 24932 38054
rect 24988 38052 24994 38054
rect 24686 38043 24994 38052
rect 24686 37020 24994 37029
rect 24686 37018 24692 37020
rect 24748 37018 24772 37020
rect 24828 37018 24852 37020
rect 24908 37018 24932 37020
rect 24988 37018 24994 37020
rect 24748 36966 24750 37018
rect 24930 36966 24932 37018
rect 24686 36964 24692 36966
rect 24748 36964 24772 36966
rect 24828 36964 24852 36966
rect 24908 36964 24932 36966
rect 24988 36964 24994 36966
rect 24686 36955 24994 36964
rect 25136 36100 25188 36106
rect 25136 36042 25188 36048
rect 25148 36009 25176 36042
rect 25134 36000 25190 36009
rect 24686 35932 24994 35941
rect 25134 35935 25190 35944
rect 24686 35930 24692 35932
rect 24748 35930 24772 35932
rect 24828 35930 24852 35932
rect 24908 35930 24932 35932
rect 24988 35930 24994 35932
rect 24748 35878 24750 35930
rect 24930 35878 24932 35930
rect 24686 35876 24692 35878
rect 24748 35876 24772 35878
rect 24828 35876 24852 35878
rect 24908 35876 24932 35878
rect 24988 35876 24994 35878
rect 24686 35867 24994 35876
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 24686 34844 24994 34853
rect 24686 34842 24692 34844
rect 24748 34842 24772 34844
rect 24828 34842 24852 34844
rect 24908 34842 24932 34844
rect 24988 34842 24994 34844
rect 24748 34790 24750 34842
rect 24930 34790 24932 34842
rect 24686 34788 24692 34790
rect 24748 34788 24772 34790
rect 24828 34788 24852 34790
rect 24908 34788 24932 34790
rect 24988 34788 24994 34790
rect 24686 34779 24994 34788
rect 24686 33756 24994 33765
rect 24686 33754 24692 33756
rect 24748 33754 24772 33756
rect 24828 33754 24852 33756
rect 24908 33754 24932 33756
rect 24988 33754 24994 33756
rect 24748 33702 24750 33754
rect 24930 33702 24932 33754
rect 24686 33700 24692 33702
rect 24748 33700 24772 33702
rect 24828 33700 24852 33702
rect 24908 33700 24932 33702
rect 24988 33700 24994 33702
rect 24686 33691 24994 33700
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 24686 32668 24994 32677
rect 24686 32666 24692 32668
rect 24748 32666 24772 32668
rect 24828 32666 24852 32668
rect 24908 32666 24932 32668
rect 24988 32666 24994 32668
rect 24748 32614 24750 32666
rect 24930 32614 24932 32666
rect 24686 32612 24692 32614
rect 24748 32612 24772 32614
rect 24828 32612 24852 32614
rect 24908 32612 24932 32614
rect 24988 32612 24994 32614
rect 24686 32603 24994 32612
rect 24686 31580 24994 31589
rect 24686 31578 24692 31580
rect 24748 31578 24772 31580
rect 24828 31578 24852 31580
rect 24908 31578 24932 31580
rect 24988 31578 24994 31580
rect 24748 31526 24750 31578
rect 24930 31526 24932 31578
rect 24686 31524 24692 31526
rect 24748 31524 24772 31526
rect 24828 31524 24852 31526
rect 24908 31524 24932 31526
rect 24988 31524 24994 31526
rect 24686 31515 24994 31524
rect 24504 30790 24624 30818
rect 24596 30734 24624 30790
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24400 30048 24452 30054
rect 24398 30016 24400 30025
rect 24452 30016 24454 30025
rect 24398 29951 24454 29960
rect 24400 28960 24452 28966
rect 24398 28928 24400 28937
rect 24452 28928 24454 28937
rect 24398 28863 24454 28872
rect 24400 27872 24452 27878
rect 24398 27840 24400 27849
rect 24452 27840 24454 27849
rect 24398 27775 24454 27784
rect 24400 26784 24452 26790
rect 24398 26752 24400 26761
rect 24452 26752 24454 26761
rect 24398 26687 24454 26696
rect 24492 26512 24544 26518
rect 24492 26454 24544 26460
rect 24308 26036 24360 26042
rect 24308 25978 24360 25984
rect 24400 25696 24452 25702
rect 24398 25664 24400 25673
rect 24452 25664 24454 25673
rect 24398 25599 24454 25608
rect 24216 24812 24268 24818
rect 24216 24754 24268 24760
rect 24308 24676 24360 24682
rect 24308 24618 24360 24624
rect 24216 22024 24268 22030
rect 24216 21966 24268 21972
rect 24228 21146 24256 21966
rect 24216 21140 24268 21146
rect 24216 21082 24268 21088
rect 24216 20800 24268 20806
rect 24216 20742 24268 20748
rect 24228 20466 24256 20742
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24216 20256 24268 20262
rect 24216 20198 24268 20204
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 23860 19230 23980 19258
rect 23848 19168 23900 19174
rect 23846 19136 23848 19145
rect 23900 19136 23902 19145
rect 23846 19071 23902 19080
rect 23480 18896 23532 18902
rect 23480 18838 23532 18844
rect 23388 18760 23440 18766
rect 23388 18702 23440 18708
rect 23492 17882 23520 18838
rect 23664 18828 23716 18834
rect 23664 18770 23716 18776
rect 23572 18080 23624 18086
rect 23572 18022 23624 18028
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 23018 17232 23074 17241
rect 23018 17167 23074 17176
rect 22928 16584 22980 16590
rect 22928 16526 22980 16532
rect 23032 16402 23060 17167
rect 22664 15694 22784 15722
rect 22940 16374 23060 16402
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22480 15162 22508 15438
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22204 14414 22232 14758
rect 22468 14544 22520 14550
rect 22572 14498 22600 14758
rect 22520 14492 22600 14498
rect 22468 14486 22600 14492
rect 22480 14470 22600 14486
rect 22480 14414 22508 14470
rect 22192 14408 22244 14414
rect 22192 14350 22244 14356
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22190 13696 22246 13705
rect 22190 13631 22246 13640
rect 22204 12986 22232 13631
rect 22296 13462 22324 14010
rect 22468 13932 22520 13938
rect 22468 13874 22520 13880
rect 22284 13456 22336 13462
rect 22284 13398 22336 13404
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22376 12912 22428 12918
rect 22112 12850 22232 12866
rect 22376 12854 22428 12860
rect 22112 12844 22244 12850
rect 22112 12838 22192 12844
rect 22192 12786 22244 12792
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 21719 12540 22027 12549
rect 21719 12538 21725 12540
rect 21781 12538 21805 12540
rect 21861 12538 21885 12540
rect 21941 12538 21965 12540
rect 22021 12538 22027 12540
rect 21781 12486 21783 12538
rect 21963 12486 21965 12538
rect 21719 12484 21725 12486
rect 21781 12484 21805 12486
rect 21861 12484 21885 12486
rect 21941 12484 21965 12486
rect 22021 12484 22027 12486
rect 21719 12475 22027 12484
rect 21652 12406 21772 12434
rect 21548 12378 21600 12384
rect 21640 12164 21692 12170
rect 21640 12106 21692 12112
rect 21652 11762 21680 12106
rect 21744 11762 21772 12406
rect 22112 12238 22140 12650
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21468 10118 21588 10146
rect 21456 9988 21508 9994
rect 21456 9930 21508 9936
rect 21468 8378 21496 9930
rect 21560 9926 21588 10118
rect 21548 9920 21600 9926
rect 21548 9862 21600 9868
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21560 8498 21588 9658
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21468 8350 21588 8378
rect 21192 8248 21404 8276
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21088 7880 21140 7886
rect 21088 7822 21140 7828
rect 20916 7534 21036 7562
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 7002 20852 7142
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20628 6870 20680 6876
rect 20718 6896 20774 6905
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 6322 20576 6598
rect 20640 6322 20668 6870
rect 20774 6854 20852 6882
rect 20718 6831 20774 6840
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20718 5264 20774 5273
rect 20718 5199 20774 5208
rect 20732 5098 20760 5199
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20536 4616 20588 4622
rect 20536 4558 20588 4564
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20548 4282 20576 4558
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20076 4014 20128 4020
rect 19984 3732 20036 3738
rect 20088 3720 20116 4014
rect 20036 3692 20116 3720
rect 19984 3674 20036 3680
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 19798 2680 19854 2689
rect 19798 2615 19854 2624
rect 19812 2514 19840 2615
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19892 2372 19944 2378
rect 19892 2314 19944 2320
rect 19904 1970 19932 2314
rect 19892 1964 19944 1970
rect 19892 1906 19944 1912
rect 19536 1686 19748 1714
rect 19432 1556 19484 1562
rect 19432 1498 19484 1504
rect 19536 160 19564 1686
rect 18970 54 19196 82
rect 18970 0 19026 54
rect 19246 0 19302 160
rect 19522 0 19578 160
rect 19798 82 19854 160
rect 19996 82 20024 2790
rect 20088 1902 20116 3692
rect 20272 3998 20484 4026
rect 20272 2774 20300 3998
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 20534 3904 20590 3913
rect 20180 2746 20300 2774
rect 20076 1896 20128 1902
rect 20076 1838 20128 1844
rect 20088 160 20116 1838
rect 20180 1562 20208 2746
rect 20352 1760 20404 1766
rect 20352 1702 20404 1708
rect 20168 1556 20220 1562
rect 20168 1498 20220 1504
rect 20364 160 20392 1702
rect 20456 649 20484 3878
rect 20534 3839 20590 3848
rect 20548 1562 20576 3839
rect 20640 3738 20668 4558
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20732 3534 20760 4762
rect 20824 3942 20852 6854
rect 20916 6798 20944 7346
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 20902 6488 20958 6497
rect 20902 6423 20958 6432
rect 20916 6322 20944 6423
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20904 6112 20956 6118
rect 20902 6080 20904 6089
rect 20956 6080 20958 6089
rect 20902 6015 20958 6024
rect 21008 5794 21036 7534
rect 21100 7002 21128 7822
rect 21088 6996 21140 7002
rect 21088 6938 21140 6944
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 21100 6497 21128 6666
rect 21086 6488 21142 6497
rect 21086 6423 21142 6432
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 5914 21128 6258
rect 21192 5914 21220 8248
rect 21560 7342 21588 8350
rect 21548 7336 21600 7342
rect 21548 7278 21600 7284
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21284 6662 21312 6938
rect 21376 6798 21404 7142
rect 21454 6896 21510 6905
rect 21454 6831 21510 6840
rect 21468 6798 21496 6831
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21456 6792 21508 6798
rect 21456 6734 21508 6740
rect 21652 6662 21680 11698
rect 21836 11694 21864 12038
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21719 11452 22027 11461
rect 21719 11450 21725 11452
rect 21781 11450 21805 11452
rect 21861 11450 21885 11452
rect 21941 11450 21965 11452
rect 22021 11450 22027 11452
rect 21781 11398 21783 11450
rect 21963 11398 21965 11450
rect 21719 11396 21725 11398
rect 21781 11396 21805 11398
rect 21861 11396 21885 11398
rect 21941 11396 21965 11398
rect 22021 11396 22027 11398
rect 21719 11387 22027 11396
rect 22296 11014 22324 12378
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22388 10810 22416 12854
rect 22480 11150 22508 13874
rect 22664 12986 22692 15694
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 15162 22784 15302
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 22836 14952 22888 14958
rect 22836 14894 22888 14900
rect 22744 14272 22796 14278
rect 22744 14214 22796 14220
rect 22756 13938 22784 14214
rect 22848 14006 22876 14894
rect 22836 14000 22888 14006
rect 22836 13942 22888 13948
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22652 12640 22704 12646
rect 22558 12608 22614 12617
rect 22652 12582 22704 12588
rect 22558 12543 22614 12552
rect 22468 11144 22520 11150
rect 22468 11086 22520 11092
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 21719 10364 22027 10373
rect 21719 10362 21725 10364
rect 21781 10362 21805 10364
rect 21861 10362 21885 10364
rect 21941 10362 21965 10364
rect 22021 10362 22027 10364
rect 21781 10310 21783 10362
rect 21963 10310 21965 10362
rect 21719 10308 21725 10310
rect 21781 10308 21805 10310
rect 21861 10308 21885 10310
rect 21941 10308 21965 10310
rect 22021 10308 22027 10310
rect 21719 10299 22027 10308
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 21836 9722 21864 9862
rect 22296 9722 22324 9862
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22100 9376 22152 9382
rect 22100 9318 22152 9324
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 21719 9276 22027 9285
rect 21719 9274 21725 9276
rect 21781 9274 21805 9276
rect 21861 9274 21885 9276
rect 21941 9274 21965 9276
rect 22021 9274 22027 9276
rect 21781 9222 21783 9274
rect 21963 9222 21965 9274
rect 21719 9220 21725 9222
rect 21781 9220 21805 9222
rect 21861 9220 21885 9222
rect 21941 9220 21965 9222
rect 22021 9220 22027 9222
rect 21719 9211 22027 9220
rect 22112 8498 22140 9318
rect 22204 8634 22232 9318
rect 22388 8974 22416 10406
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22480 9178 22508 9998
rect 22468 9172 22520 9178
rect 22468 9114 22520 9120
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22192 8628 22244 8634
rect 22192 8570 22244 8576
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21719 8188 22027 8197
rect 21719 8186 21725 8188
rect 21781 8186 21805 8188
rect 21861 8186 21885 8188
rect 21941 8186 21965 8188
rect 22021 8186 22027 8188
rect 21781 8134 21783 8186
rect 21963 8134 21965 8186
rect 21719 8132 21725 8134
rect 21781 8132 21805 8134
rect 21861 8132 21885 8134
rect 21941 8132 21965 8134
rect 22021 8132 22027 8134
rect 21719 8123 22027 8132
rect 22296 7868 22324 8910
rect 22468 8560 22520 8566
rect 22468 8502 22520 8508
rect 22480 8430 22508 8502
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22468 8084 22520 8090
rect 22468 8026 22520 8032
rect 22376 7880 22428 7886
rect 22296 7840 22376 7868
rect 22376 7822 22428 7828
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 21719 7100 22027 7109
rect 21719 7098 21725 7100
rect 21781 7098 21805 7100
rect 21861 7098 21885 7100
rect 21941 7098 21965 7100
rect 22021 7098 22027 7100
rect 21781 7046 21783 7098
rect 21963 7046 21965 7098
rect 21719 7044 21725 7046
rect 21781 7044 21805 7046
rect 21861 7044 21885 7046
rect 21941 7044 21965 7046
rect 22021 7044 22027 7046
rect 21719 7035 22027 7044
rect 22112 6984 22140 7278
rect 22296 7002 22324 7686
rect 21836 6956 22140 6984
rect 22192 6996 22244 7002
rect 21836 6769 21864 6956
rect 22192 6938 22244 6944
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22204 6882 22232 6938
rect 22204 6854 22324 6882
rect 21916 6792 21968 6798
rect 21822 6760 21878 6769
rect 22192 6792 22244 6798
rect 21968 6752 22140 6780
rect 21916 6734 21968 6740
rect 21822 6695 21878 6704
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21468 6322 21496 6394
rect 21364 6316 21416 6322
rect 21284 6276 21364 6304
rect 21284 6118 21312 6276
rect 21364 6258 21416 6264
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21362 6216 21418 6225
rect 21362 6151 21418 6160
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 21376 5914 21404 6151
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 21180 5908 21232 5914
rect 21180 5850 21232 5856
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21008 5766 21312 5794
rect 20996 5704 21048 5710
rect 21048 5664 21128 5692
rect 20996 5646 21048 5652
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 4622 20944 5510
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21008 4690 21036 5102
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20902 4040 20958 4049
rect 20902 3975 20958 3984
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 20810 3632 20866 3641
rect 20916 3602 20944 3975
rect 20810 3567 20866 3576
rect 20904 3596 20956 3602
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20718 2952 20774 2961
rect 20824 2922 20852 3567
rect 20904 3538 20956 3544
rect 20916 3194 20944 3538
rect 20996 3460 21048 3466
rect 20996 3402 21048 3408
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20718 2887 20720 2896
rect 20772 2887 20774 2896
rect 20812 2916 20864 2922
rect 20720 2858 20772 2864
rect 20812 2858 20864 2864
rect 20718 2816 20774 2825
rect 20718 2751 20774 2760
rect 20732 2446 20760 2751
rect 20916 2446 20944 3130
rect 21008 3126 21036 3402
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20904 1964 20956 1970
rect 20904 1906 20956 1912
rect 20628 1760 20680 1766
rect 20628 1702 20680 1708
rect 20536 1556 20588 1562
rect 20536 1498 20588 1504
rect 20536 1352 20588 1358
rect 20536 1294 20588 1300
rect 20548 746 20576 1294
rect 20536 740 20588 746
rect 20536 682 20588 688
rect 20442 640 20498 649
rect 20442 575 20498 584
rect 20640 160 20668 1702
rect 20916 160 20944 1906
rect 21100 1329 21128 5664
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21192 4826 21220 5170
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21284 4706 21312 5766
rect 21468 5624 21496 6258
rect 21836 6254 21864 6695
rect 21824 6248 21876 6254
rect 21914 6216 21970 6225
rect 21876 6196 21914 6202
rect 21824 6190 21914 6196
rect 21836 6174 21914 6190
rect 21914 6151 21970 6160
rect 21640 6112 21692 6118
rect 21560 6089 21640 6100
rect 21546 6080 21640 6089
rect 21602 6072 21640 6080
rect 21640 6054 21692 6060
rect 21546 6015 21602 6024
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 22112 5817 22140 6752
rect 22192 6734 22244 6740
rect 22204 6458 22232 6734
rect 22296 6730 22324 6854
rect 22284 6724 22336 6730
rect 22284 6666 22336 6672
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22282 6216 22338 6225
rect 22282 6151 22338 6160
rect 22098 5808 22154 5817
rect 22098 5743 22154 5752
rect 21824 5636 21876 5642
rect 21468 5596 21824 5624
rect 21824 5578 21876 5584
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21928 5234 21956 5306
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 21192 4678 21312 4706
rect 21192 3380 21220 4678
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21284 3505 21312 4218
rect 21270 3496 21326 3505
rect 21270 3431 21326 3440
rect 21192 3352 21312 3380
rect 21284 3074 21312 3352
rect 21376 3194 21404 4966
rect 21468 4049 21496 5102
rect 21560 4826 21588 5170
rect 22020 5137 22048 5170
rect 22006 5128 22062 5137
rect 22006 5063 22062 5072
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 22112 4826 22140 5578
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 21546 4720 21602 4729
rect 21546 4655 21602 4664
rect 21454 4040 21510 4049
rect 21454 3975 21510 3984
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21468 3534 21496 3878
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21180 3052 21232 3058
rect 21284 3046 21404 3074
rect 21180 2994 21232 3000
rect 21192 2774 21220 2994
rect 21192 2746 21312 2774
rect 21284 1902 21312 2746
rect 21376 2038 21404 3046
rect 21560 2990 21588 4655
rect 21640 4616 21692 4622
rect 21640 4558 21692 4564
rect 21652 4282 21680 4558
rect 21732 4480 21784 4486
rect 21732 4422 21784 4428
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21744 3924 21772 4422
rect 22204 4162 22232 5510
rect 22296 4622 22324 6151
rect 22388 5710 22416 7822
rect 22480 6322 22508 8026
rect 22572 7478 22600 12543
rect 22664 11234 22692 12582
rect 22940 12434 22968 16374
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23124 14074 23152 14214
rect 23020 14068 23072 14074
rect 23020 14010 23072 14016
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23032 13954 23060 14010
rect 23032 13938 23152 13954
rect 23032 13932 23164 13938
rect 23032 13926 23112 13932
rect 23112 13874 23164 13880
rect 23216 13818 23244 17478
rect 23492 16250 23520 17818
rect 23584 16590 23612 18022
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23480 16244 23532 16250
rect 23480 16186 23532 16192
rect 23676 16046 23704 18770
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23860 16250 23888 17138
rect 23952 16810 23980 19230
rect 24228 18442 24256 20198
rect 24320 18834 24348 24618
rect 24400 24608 24452 24614
rect 24398 24576 24400 24585
rect 24452 24576 24454 24585
rect 24398 24511 24454 24520
rect 24400 23520 24452 23526
rect 24398 23488 24400 23497
rect 24452 23488 24454 23497
rect 24398 23423 24454 23432
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24412 19334 24440 23258
rect 24504 22710 24532 26454
rect 24492 22704 24544 22710
rect 24492 22646 24544 22652
rect 24490 22400 24546 22409
rect 24490 22335 24546 22344
rect 24504 21690 24532 22335
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24412 19306 24532 19334
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24136 18414 24256 18442
rect 24136 17082 24164 18414
rect 24400 18080 24452 18086
rect 24398 18048 24400 18057
rect 24452 18048 24454 18057
rect 24398 17983 24454 17992
rect 24504 17898 24532 19306
rect 24412 17870 24532 17898
rect 24308 17672 24360 17678
rect 24308 17614 24360 17620
rect 24136 17054 24256 17082
rect 24124 16992 24176 16998
rect 24122 16960 24124 16969
rect 24176 16960 24178 16969
rect 24122 16895 24178 16904
rect 23952 16782 24072 16810
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23952 16561 23980 16594
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 23664 16040 23716 16046
rect 23664 15982 23716 15988
rect 23664 15904 23716 15910
rect 23664 15846 23716 15852
rect 23676 15026 23704 15846
rect 23848 15700 23900 15706
rect 23848 15642 23900 15648
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23768 14482 23796 15302
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23124 13790 23244 13818
rect 23018 12608 23074 12617
rect 23124 12594 23152 13790
rect 23308 13546 23336 13874
rect 23388 13864 23440 13870
rect 23388 13806 23440 13812
rect 23216 13530 23336 13546
rect 23204 13524 23336 13530
rect 23256 13518 23336 13524
rect 23204 13466 23256 13472
rect 23204 13252 23256 13258
rect 23204 13194 23256 13200
rect 23074 12566 23152 12594
rect 23018 12543 23074 12552
rect 23216 12434 23244 13194
rect 23400 12986 23428 13806
rect 23480 13796 23532 13802
rect 23480 13738 23532 13744
rect 23492 13433 23520 13738
rect 23478 13424 23534 13433
rect 23478 13359 23534 13368
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 22940 12406 23060 12434
rect 23216 12406 23336 12434
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 22756 11898 22784 12174
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22848 11898 22876 12038
rect 22744 11892 22796 11898
rect 22744 11834 22796 11840
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 23032 11370 23060 12406
rect 23112 12096 23164 12102
rect 23112 12038 23164 12044
rect 23124 11898 23152 12038
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23204 11756 23256 11762
rect 23308 11744 23336 12406
rect 23492 11898 23520 13262
rect 23860 12238 23888 15642
rect 24044 14906 24072 16782
rect 24122 15872 24178 15881
rect 24122 15807 24178 15816
rect 24136 15706 24164 15807
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24228 15162 24256 17054
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24044 14878 24164 14906
rect 24032 14816 24084 14822
rect 24030 14784 24032 14793
rect 24084 14784 24086 14793
rect 24030 14719 24086 14728
rect 24136 14346 24164 14878
rect 24124 14340 24176 14346
rect 24124 14282 24176 14288
rect 24228 14278 24256 14962
rect 24216 14272 24268 14278
rect 24216 14214 24268 14220
rect 24216 12640 24268 12646
rect 24214 12608 24216 12617
rect 24268 12608 24270 12617
rect 24214 12543 24270 12552
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23256 11716 23336 11744
rect 23480 11756 23532 11762
rect 23204 11698 23256 11704
rect 23480 11698 23532 11704
rect 23032 11342 23152 11370
rect 23216 11354 23244 11698
rect 23492 11354 23520 11698
rect 23848 11552 23900 11558
rect 23846 11520 23848 11529
rect 23900 11520 23902 11529
rect 23846 11455 23902 11464
rect 22664 11206 23060 11234
rect 22652 11144 22704 11150
rect 22928 11144 22980 11150
rect 22704 11092 22928 11098
rect 22652 11086 22980 11092
rect 22664 11070 22968 11086
rect 22744 11008 22796 11014
rect 22744 10950 22796 10956
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22560 5704 22612 5710
rect 22560 5646 22612 5652
rect 22572 5098 22600 5646
rect 22664 5642 22692 10746
rect 22756 10606 22784 10950
rect 22744 10600 22796 10606
rect 22744 10542 22796 10548
rect 22756 10062 22784 10542
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22756 9518 22784 9998
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22756 8566 22784 9046
rect 22848 8838 22876 9590
rect 22836 8832 22888 8838
rect 22836 8774 22888 8780
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22744 8288 22796 8294
rect 22744 8230 22796 8236
rect 22756 8022 22784 8230
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22940 7970 22968 11070
rect 23032 10062 23060 11206
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23032 8090 23060 8434
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 22940 7942 23060 7970
rect 22744 6928 22796 6934
rect 22744 6870 22796 6876
rect 22756 6458 22784 6870
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22928 6656 22980 6662
rect 22928 6598 22980 6604
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22848 6322 22876 6598
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22742 5536 22798 5545
rect 22742 5471 22798 5480
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22296 4282 22324 4558
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22204 4134 22324 4162
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21652 3896 21772 3924
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 21548 2440 21600 2446
rect 21468 2400 21548 2428
rect 21364 2032 21416 2038
rect 21364 1974 21416 1980
rect 21272 1896 21324 1902
rect 21272 1838 21324 1844
rect 21362 1456 21418 1465
rect 21362 1391 21364 1400
rect 21416 1391 21418 1400
rect 21364 1362 21416 1368
rect 21086 1320 21142 1329
rect 20996 1284 21048 1290
rect 21086 1255 21142 1264
rect 21180 1284 21232 1290
rect 20996 1226 21048 1232
rect 21180 1226 21232 1232
rect 21008 678 21036 1226
rect 21088 1216 21140 1222
rect 21088 1158 21140 1164
rect 21100 950 21128 1158
rect 21192 1018 21220 1226
rect 21272 1216 21324 1222
rect 21272 1158 21324 1164
rect 21180 1012 21232 1018
rect 21180 954 21232 960
rect 21088 944 21140 950
rect 21088 886 21140 892
rect 21284 882 21312 1158
rect 21272 876 21324 882
rect 21272 818 21324 824
rect 20996 672 21048 678
rect 20996 614 21048 620
rect 21180 468 21232 474
rect 21180 410 21232 416
rect 21192 160 21220 410
rect 21468 160 21496 2400
rect 21548 2382 21600 2388
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21560 2038 21588 2246
rect 21548 2032 21600 2038
rect 21548 1974 21600 1980
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 19798 54 20024 82
rect 19798 0 19854 54
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20626 0 20682 160
rect 20902 0 20958 160
rect 21178 0 21234 160
rect 21454 0 21510 160
rect 21560 82 21588 1838
rect 21652 1358 21680 3896
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 22112 3398 22140 4014
rect 22100 3392 22152 3398
rect 22100 3334 22152 3340
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21836 1902 21864 2382
rect 21824 1896 21876 1902
rect 21824 1838 21876 1844
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 22112 1494 22140 3334
rect 22100 1488 22152 1494
rect 22100 1430 22152 1436
rect 21640 1352 21692 1358
rect 21640 1294 21692 1300
rect 21916 1284 21968 1290
rect 21916 1226 21968 1232
rect 22100 1284 22152 1290
rect 22100 1226 22152 1232
rect 21928 610 21956 1226
rect 22112 814 22140 1226
rect 22204 1222 22232 4014
rect 22296 3942 22324 4134
rect 22284 3936 22336 3942
rect 22284 3878 22336 3884
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22192 1216 22244 1222
rect 22192 1158 22244 1164
rect 22100 808 22152 814
rect 22100 750 22152 756
rect 22008 672 22060 678
rect 22008 614 22060 620
rect 21916 604 21968 610
rect 21916 546 21968 552
rect 22020 160 22048 614
rect 22296 160 22324 3470
rect 22388 1562 22416 4966
rect 22480 4146 22508 4966
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 22572 2972 22600 5034
rect 22664 4185 22692 5170
rect 22756 4622 22784 5471
rect 22940 5234 22968 6598
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22836 4480 22888 4486
rect 22836 4422 22888 4428
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22650 4176 22706 4185
rect 22650 4111 22706 4120
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22652 4004 22704 4010
rect 22652 3946 22704 3952
rect 22664 3097 22692 3946
rect 22650 3088 22706 3097
rect 22650 3023 22706 3032
rect 22572 2944 22692 2972
rect 22468 2508 22520 2514
rect 22468 2450 22520 2456
rect 22480 1562 22508 2450
rect 22664 2446 22692 2944
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22376 1556 22428 1562
rect 22376 1498 22428 1504
rect 22468 1556 22520 1562
rect 22468 1498 22520 1504
rect 22468 1352 22520 1358
rect 22468 1294 22520 1300
rect 22480 474 22508 1294
rect 22468 468 22520 474
rect 22468 410 22520 416
rect 21730 82 21786 160
rect 21560 54 21786 82
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 0 22338 160
rect 22558 82 22614 160
rect 22756 82 22784 4082
rect 22848 2106 22876 4422
rect 22836 2100 22888 2106
rect 22836 2042 22888 2048
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22848 160 22876 1498
rect 22940 1290 22968 4422
rect 23032 3058 23060 7942
rect 23124 3670 23152 11342
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23386 10432 23442 10441
rect 23386 10367 23442 10376
rect 23400 9178 23428 10367
rect 23756 9920 23808 9926
rect 23756 9862 23808 9868
rect 23388 9172 23440 9178
rect 23388 9114 23440 9120
rect 23572 8968 23624 8974
rect 23570 8936 23572 8945
rect 23624 8936 23626 8945
rect 23570 8871 23626 8880
rect 23768 8634 23796 9862
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24124 9376 24176 9382
rect 24030 9344 24086 9353
rect 24124 9318 24176 9324
rect 24030 9279 24086 9288
rect 24044 9178 24072 9279
rect 24136 9178 24164 9318
rect 24032 9172 24084 9178
rect 24032 9114 24084 9120
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 23296 8628 23348 8634
rect 23296 8570 23348 8576
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23204 6792 23256 6798
rect 23202 6760 23204 6769
rect 23256 6760 23258 6769
rect 23202 6695 23258 6704
rect 23204 6656 23256 6662
rect 23204 6598 23256 6604
rect 23216 4826 23244 6598
rect 23308 6118 23336 8570
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23572 8424 23624 8430
rect 23572 8366 23624 8372
rect 23584 7546 23612 8366
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23676 7546 23704 7822
rect 23940 7812 23992 7818
rect 23940 7754 23992 7760
rect 23952 7546 23980 7754
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23664 7540 23716 7546
rect 23664 7482 23716 7488
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23584 6798 23612 7482
rect 23754 7168 23810 7177
rect 23754 7103 23810 7112
rect 23662 6896 23718 6905
rect 23662 6831 23718 6840
rect 23388 6792 23440 6798
rect 23572 6792 23624 6798
rect 23440 6752 23520 6780
rect 23388 6734 23440 6740
rect 23386 6488 23442 6497
rect 23386 6423 23388 6432
rect 23440 6423 23442 6432
rect 23388 6394 23440 6400
rect 23386 6352 23442 6361
rect 23386 6287 23442 6296
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23308 4486 23336 5646
rect 23400 5642 23428 6287
rect 23388 5636 23440 5642
rect 23388 5578 23440 5584
rect 23386 5536 23442 5545
rect 23386 5471 23442 5480
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 23216 3738 23244 4218
rect 23400 4146 23428 5471
rect 23492 5114 23520 6752
rect 23572 6734 23624 6740
rect 23572 6112 23624 6118
rect 23676 6089 23704 6831
rect 23768 6322 23796 7103
rect 24044 6866 24072 8434
rect 24228 7290 24256 9454
rect 24320 9217 24348 17614
rect 24412 17082 24440 17870
rect 24596 17678 24624 30534
rect 24686 30492 24994 30501
rect 24686 30490 24692 30492
rect 24748 30490 24772 30492
rect 24828 30490 24852 30492
rect 24908 30490 24932 30492
rect 24988 30490 24994 30492
rect 24748 30438 24750 30490
rect 24930 30438 24932 30490
rect 24686 30436 24692 30438
rect 24748 30436 24772 30438
rect 24828 30436 24852 30438
rect 24908 30436 24932 30438
rect 24988 30436 24994 30438
rect 24686 30427 24994 30436
rect 24686 29404 24994 29413
rect 24686 29402 24692 29404
rect 24748 29402 24772 29404
rect 24828 29402 24852 29404
rect 24908 29402 24932 29404
rect 24988 29402 24994 29404
rect 24748 29350 24750 29402
rect 24930 29350 24932 29402
rect 24686 29348 24692 29350
rect 24748 29348 24772 29350
rect 24828 29348 24852 29350
rect 24908 29348 24932 29350
rect 24988 29348 24994 29350
rect 24686 29339 24994 29348
rect 24686 28316 24994 28325
rect 24686 28314 24692 28316
rect 24748 28314 24772 28316
rect 24828 28314 24852 28316
rect 24908 28314 24932 28316
rect 24988 28314 24994 28316
rect 24748 28262 24750 28314
rect 24930 28262 24932 28314
rect 24686 28260 24692 28262
rect 24748 28260 24772 28262
rect 24828 28260 24852 28262
rect 24908 28260 24932 28262
rect 24988 28260 24994 28262
rect 24686 28251 24994 28260
rect 24686 27228 24994 27237
rect 24686 27226 24692 27228
rect 24748 27226 24772 27228
rect 24828 27226 24852 27228
rect 24908 27226 24932 27228
rect 24988 27226 24994 27228
rect 24748 27174 24750 27226
rect 24930 27174 24932 27226
rect 24686 27172 24692 27174
rect 24748 27172 24772 27174
rect 24828 27172 24852 27174
rect 24908 27172 24932 27174
rect 24988 27172 24994 27174
rect 24686 27163 24994 27172
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 24872 26518 24900 26930
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 24686 26140 24994 26149
rect 24686 26138 24692 26140
rect 24748 26138 24772 26140
rect 24828 26138 24852 26140
rect 24908 26138 24932 26140
rect 24988 26138 24994 26140
rect 24748 26086 24750 26138
rect 24930 26086 24932 26138
rect 24686 26084 24692 26086
rect 24748 26084 24772 26086
rect 24828 26084 24852 26086
rect 24908 26084 24932 26086
rect 24988 26084 24994 26086
rect 24686 26075 24994 26084
rect 24686 25052 24994 25061
rect 24686 25050 24692 25052
rect 24748 25050 24772 25052
rect 24828 25050 24852 25052
rect 24908 25050 24932 25052
rect 24988 25050 24994 25052
rect 24748 24998 24750 25050
rect 24930 24998 24932 25050
rect 24686 24996 24692 24998
rect 24748 24996 24772 24998
rect 24828 24996 24852 24998
rect 24908 24996 24932 24998
rect 24988 24996 24994 24998
rect 24686 24987 24994 24996
rect 24686 23964 24994 23973
rect 24686 23962 24692 23964
rect 24748 23962 24772 23964
rect 24828 23962 24852 23964
rect 24908 23962 24932 23964
rect 24988 23962 24994 23964
rect 24748 23910 24750 23962
rect 24930 23910 24932 23962
rect 24686 23908 24692 23910
rect 24748 23908 24772 23910
rect 24828 23908 24852 23910
rect 24908 23908 24932 23910
rect 24988 23908 24994 23910
rect 24686 23899 24994 23908
rect 24686 22876 24994 22885
rect 24686 22874 24692 22876
rect 24748 22874 24772 22876
rect 24828 22874 24852 22876
rect 24908 22874 24932 22876
rect 24988 22874 24994 22876
rect 24748 22822 24750 22874
rect 24930 22822 24932 22874
rect 24686 22820 24692 22822
rect 24748 22820 24772 22822
rect 24828 22820 24852 22822
rect 24908 22820 24932 22822
rect 24988 22820 24994 22822
rect 24686 22811 24994 22820
rect 24686 21788 24994 21797
rect 24686 21786 24692 21788
rect 24748 21786 24772 21788
rect 24828 21786 24852 21788
rect 24908 21786 24932 21788
rect 24988 21786 24994 21788
rect 24748 21734 24750 21786
rect 24930 21734 24932 21786
rect 24686 21732 24692 21734
rect 24748 21732 24772 21734
rect 24828 21732 24852 21734
rect 24908 21732 24932 21734
rect 24988 21732 24994 21734
rect 24686 21723 24994 21732
rect 24686 20700 24994 20709
rect 24686 20698 24692 20700
rect 24748 20698 24772 20700
rect 24828 20698 24852 20700
rect 24908 20698 24932 20700
rect 24988 20698 24994 20700
rect 24748 20646 24750 20698
rect 24930 20646 24932 20698
rect 24686 20644 24692 20646
rect 24748 20644 24772 20646
rect 24828 20644 24852 20646
rect 24908 20644 24932 20646
rect 24988 20644 24994 20646
rect 24686 20635 24994 20644
rect 24686 19612 24994 19621
rect 24686 19610 24692 19612
rect 24748 19610 24772 19612
rect 24828 19610 24852 19612
rect 24908 19610 24932 19612
rect 24988 19610 24994 19612
rect 24748 19558 24750 19610
rect 24930 19558 24932 19610
rect 24686 19556 24692 19558
rect 24748 19556 24772 19558
rect 24828 19556 24852 19558
rect 24908 19556 24932 19558
rect 24988 19556 24994 19558
rect 24686 19547 24994 19556
rect 24686 18524 24994 18533
rect 24686 18522 24692 18524
rect 24748 18522 24772 18524
rect 24828 18522 24852 18524
rect 24908 18522 24932 18524
rect 24988 18522 24994 18524
rect 24748 18470 24750 18522
rect 24930 18470 24932 18522
rect 24686 18468 24692 18470
rect 24748 18468 24772 18470
rect 24828 18468 24852 18470
rect 24908 18468 24932 18470
rect 24988 18468 24994 18470
rect 24686 18459 24994 18468
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 25056 17524 25084 32778
rect 25148 32586 25176 35702
rect 25228 34944 25280 34950
rect 25226 34912 25228 34921
rect 25280 34912 25282 34921
rect 25226 34847 25282 34856
rect 25228 33856 25280 33862
rect 25226 33824 25228 33833
rect 25280 33824 25282 33833
rect 25226 33759 25282 33768
rect 25228 32768 25280 32774
rect 25226 32736 25228 32745
rect 25280 32736 25282 32745
rect 25226 32671 25282 32680
rect 25148 32558 25268 32586
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25148 31657 25176 31758
rect 25134 31648 25190 31657
rect 25134 31583 25190 31592
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 25148 30569 25176 30602
rect 25134 30560 25190 30569
rect 25134 30495 25190 30504
rect 25136 29504 25188 29510
rect 25134 29472 25136 29481
rect 25188 29472 25190 29481
rect 25134 29407 25190 29416
rect 25136 28416 25188 28422
rect 25134 28384 25136 28393
rect 25188 28384 25190 28393
rect 25134 28319 25190 28328
rect 25136 27328 25188 27334
rect 25134 27296 25136 27305
rect 25188 27296 25190 27305
rect 25134 27231 25190 27240
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25148 26217 25176 26250
rect 25134 26208 25190 26217
rect 25134 26143 25190 26152
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25148 25129 25176 25162
rect 25134 25120 25190 25129
rect 25134 25055 25190 25064
rect 25136 24064 25188 24070
rect 25134 24032 25136 24041
rect 25188 24032 25190 24041
rect 25134 23967 25190 23976
rect 25136 22976 25188 22982
rect 25134 22944 25136 22953
rect 25188 22944 25190 22953
rect 25134 22879 25190 22888
rect 25136 21956 25188 21962
rect 25136 21898 25188 21904
rect 25148 21865 25176 21898
rect 25134 21856 25190 21865
rect 25134 21791 25190 21800
rect 25134 20768 25190 20777
rect 25134 20703 25190 20712
rect 25148 19310 25176 20703
rect 25136 19304 25188 19310
rect 25136 19246 25188 19252
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25148 18601 25176 18838
rect 25134 18592 25190 18601
rect 25134 18527 25190 18536
rect 24596 17496 25084 17524
rect 25134 17504 25190 17513
rect 24412 17054 24532 17082
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24412 16114 24440 16934
rect 24400 16108 24452 16114
rect 24400 16050 24452 16056
rect 24400 13728 24452 13734
rect 24398 13696 24400 13705
rect 24452 13696 24454 13705
rect 24398 13631 24454 13640
rect 24400 12912 24452 12918
rect 24504 12900 24532 17054
rect 24452 12872 24532 12900
rect 24400 12854 24452 12860
rect 24490 12744 24546 12753
rect 24490 12679 24546 12688
rect 24306 9208 24362 9217
rect 24306 9143 24362 9152
rect 24504 8378 24532 12679
rect 24596 8514 24624 17496
rect 24686 17436 24994 17445
rect 25134 17439 25190 17448
rect 24686 17434 24692 17436
rect 24748 17434 24772 17436
rect 24828 17434 24852 17436
rect 24908 17434 24932 17436
rect 24988 17434 24994 17436
rect 24748 17382 24750 17434
rect 24930 17382 24932 17434
rect 24686 17380 24692 17382
rect 24748 17380 24772 17382
rect 24828 17380 24852 17382
rect 24908 17380 24932 17382
rect 24988 17380 24994 17382
rect 24686 17371 24994 17380
rect 25148 17338 25176 17439
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25240 17218 25268 32558
rect 25056 17190 25268 17218
rect 24686 16348 24994 16357
rect 24686 16346 24692 16348
rect 24748 16346 24772 16348
rect 24828 16346 24852 16348
rect 24908 16346 24932 16348
rect 24988 16346 24994 16348
rect 24748 16294 24750 16346
rect 24930 16294 24932 16346
rect 24686 16292 24692 16294
rect 24748 16292 24772 16294
rect 24828 16292 24852 16294
rect 24908 16292 24932 16294
rect 24988 16292 24994 16294
rect 24686 16283 24994 16292
rect 24686 15260 24994 15269
rect 24686 15258 24692 15260
rect 24748 15258 24772 15260
rect 24828 15258 24852 15260
rect 24908 15258 24932 15260
rect 24988 15258 24994 15260
rect 24748 15206 24750 15258
rect 24930 15206 24932 15258
rect 24686 15204 24692 15206
rect 24748 15204 24772 15206
rect 24828 15204 24852 15206
rect 24908 15204 24932 15206
rect 24988 15204 24994 15206
rect 24686 15195 24994 15204
rect 24686 14172 24994 14181
rect 24686 14170 24692 14172
rect 24748 14170 24772 14172
rect 24828 14170 24852 14172
rect 24908 14170 24932 14172
rect 24988 14170 24994 14172
rect 24748 14118 24750 14170
rect 24930 14118 24932 14170
rect 24686 14116 24692 14118
rect 24748 14116 24772 14118
rect 24828 14116 24852 14118
rect 24908 14116 24932 14118
rect 24988 14116 24994 14118
rect 24686 14107 24994 14116
rect 24686 13084 24994 13093
rect 24686 13082 24692 13084
rect 24748 13082 24772 13084
rect 24828 13082 24852 13084
rect 24908 13082 24932 13084
rect 24988 13082 24994 13084
rect 24748 13030 24750 13082
rect 24930 13030 24932 13082
rect 24686 13028 24692 13030
rect 24748 13028 24772 13030
rect 24828 13028 24852 13030
rect 24908 13028 24932 13030
rect 24988 13028 24994 13030
rect 24686 13019 24994 13028
rect 24686 11996 24994 12005
rect 24686 11994 24692 11996
rect 24748 11994 24772 11996
rect 24828 11994 24852 11996
rect 24908 11994 24932 11996
rect 24988 11994 24994 11996
rect 24748 11942 24750 11994
rect 24930 11942 24932 11994
rect 24686 11940 24692 11942
rect 24748 11940 24772 11942
rect 24828 11940 24852 11942
rect 24908 11940 24932 11942
rect 24988 11940 24994 11942
rect 24686 11931 24994 11940
rect 24686 10908 24994 10917
rect 24686 10906 24692 10908
rect 24748 10906 24772 10908
rect 24828 10906 24852 10908
rect 24908 10906 24932 10908
rect 24988 10906 24994 10908
rect 24748 10854 24750 10906
rect 24930 10854 24932 10906
rect 24686 10852 24692 10854
rect 24748 10852 24772 10854
rect 24828 10852 24852 10854
rect 24908 10852 24932 10854
rect 24988 10852 24994 10854
rect 24686 10843 24994 10852
rect 24686 9820 24994 9829
rect 24686 9818 24692 9820
rect 24748 9818 24772 9820
rect 24828 9818 24852 9820
rect 24908 9818 24932 9820
rect 24988 9818 24994 9820
rect 24748 9766 24750 9818
rect 24930 9766 24932 9818
rect 24686 9764 24692 9766
rect 24748 9764 24772 9766
rect 24828 9764 24852 9766
rect 24908 9764 24932 9766
rect 24988 9764 24994 9766
rect 24686 9755 24994 9764
rect 25056 9674 25084 17190
rect 25136 14544 25188 14550
rect 25136 14486 25188 14492
rect 25148 14249 25176 14486
rect 25134 14240 25190 14249
rect 25134 14175 25190 14184
rect 25134 12744 25190 12753
rect 25134 12679 25190 12688
rect 25148 12442 25176 12679
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25228 12368 25280 12374
rect 25228 12310 25280 12316
rect 25240 12073 25268 12310
rect 25226 12064 25282 12073
rect 25226 11999 25282 12008
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25240 10985 25268 11494
rect 25226 10976 25282 10985
rect 25226 10911 25282 10920
rect 25332 10010 25360 40598
rect 25412 37664 25464 37670
rect 25412 37606 25464 37612
rect 25424 23322 25452 37606
rect 25596 36780 25648 36786
rect 25596 36722 25648 36728
rect 25504 31816 25556 31822
rect 25504 31758 25556 31764
rect 25412 23316 25464 23322
rect 25412 23258 25464 23264
rect 25516 22094 25544 31758
rect 25608 26994 25636 36722
rect 25688 32972 25740 32978
rect 25688 32914 25740 32920
rect 25596 26988 25648 26994
rect 25596 26930 25648 26936
rect 25700 26874 25728 32914
rect 25424 22066 25544 22094
rect 25608 26846 25728 26874
rect 25424 12434 25452 22066
rect 25502 19680 25558 19689
rect 25502 19615 25558 19624
rect 25516 18766 25544 19615
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25502 15328 25558 15337
rect 25502 15263 25558 15272
rect 25516 14754 25544 15263
rect 25504 14748 25556 14754
rect 25504 14690 25556 14696
rect 25424 12406 25544 12434
rect 25332 9982 25452 10010
rect 25318 9888 25374 9897
rect 25318 9823 25374 9832
rect 25056 9646 25176 9674
rect 24686 8732 24994 8741
rect 24686 8730 24692 8732
rect 24748 8730 24772 8732
rect 24828 8730 24852 8732
rect 24908 8730 24932 8732
rect 24988 8730 24994 8732
rect 24748 8678 24750 8730
rect 24930 8678 24932 8730
rect 24686 8676 24692 8678
rect 24748 8676 24772 8678
rect 24828 8676 24852 8678
rect 24908 8676 24932 8678
rect 24988 8676 24994 8678
rect 24686 8667 24994 8676
rect 24596 8486 24716 8514
rect 24504 8350 24624 8378
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24490 8256 24546 8265
rect 24320 7478 24348 8230
rect 24490 8191 24546 8200
rect 24308 7472 24360 7478
rect 24308 7414 24360 7420
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24228 7262 24348 7290
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24032 6656 24084 6662
rect 24032 6598 24084 6604
rect 23756 6316 23808 6322
rect 23756 6258 23808 6264
rect 23572 6054 23624 6060
rect 23662 6080 23718 6089
rect 23584 5914 23612 6054
rect 23662 6015 23718 6024
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 24044 5794 24072 6598
rect 23860 5766 24072 5794
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23662 5400 23718 5409
rect 23662 5335 23718 5344
rect 23492 5086 23612 5114
rect 23388 4140 23440 4146
rect 23388 4082 23440 4088
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 23112 3664 23164 3670
rect 23112 3606 23164 3612
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 23020 2032 23072 2038
rect 23020 1974 23072 1980
rect 23032 1766 23060 1974
rect 23020 1760 23072 1766
rect 23020 1702 23072 1708
rect 22928 1284 22980 1290
rect 22928 1226 22980 1232
rect 23124 160 23152 3470
rect 23584 2650 23612 5086
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23492 2310 23520 2586
rect 23480 2304 23532 2310
rect 23480 2246 23532 2252
rect 23676 1970 23704 5335
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 23768 1358 23796 5646
rect 23860 3058 23888 5766
rect 24216 4548 24268 4554
rect 24216 4490 24268 4496
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23952 2938 23980 3878
rect 24044 3126 24072 4082
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 23952 2910 24072 2938
rect 23756 1352 23808 1358
rect 23756 1294 23808 1300
rect 23204 740 23256 746
rect 23204 682 23256 688
rect 22558 54 22784 82
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23216 82 23244 682
rect 23756 604 23808 610
rect 23756 546 23808 552
rect 23386 82 23442 160
rect 23216 54 23442 82
rect 23386 0 23442 54
rect 23662 82 23718 160
rect 23768 82 23796 546
rect 23662 54 23796 82
rect 23938 82 23994 160
rect 24044 82 24072 2910
rect 24228 950 24256 4490
rect 24320 4010 24348 7262
rect 24412 6458 24440 7346
rect 24400 6452 24452 6458
rect 24400 6394 24452 6400
rect 24504 6322 24532 8191
rect 24596 7426 24624 8350
rect 24688 8294 24716 8486
rect 24676 8288 24728 8294
rect 24676 8230 24728 8236
rect 24686 7644 24994 7653
rect 24686 7642 24692 7644
rect 24748 7642 24772 7644
rect 24828 7642 24852 7644
rect 24908 7642 24932 7644
rect 24988 7642 24994 7644
rect 24748 7590 24750 7642
rect 24930 7590 24932 7642
rect 24686 7588 24692 7590
rect 24748 7588 24772 7590
rect 24828 7588 24852 7590
rect 24908 7588 24932 7590
rect 24988 7588 24994 7590
rect 24686 7579 24994 7588
rect 24596 7398 25084 7426
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24492 6316 24544 6322
rect 24492 6258 24544 6264
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24584 4208 24636 4214
rect 24584 4150 24636 4156
rect 24308 4004 24360 4010
rect 24308 3946 24360 3952
rect 24492 3460 24544 3466
rect 24492 3402 24544 3408
rect 24216 944 24268 950
rect 24216 886 24268 892
rect 24216 536 24268 542
rect 24216 478 24268 484
rect 24228 160 24256 478
rect 24504 160 24532 3402
rect 23938 54 24072 82
rect 23662 0 23718 54
rect 23938 0 23994 54
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24596 82 24624 4150
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 24872 1306 24900 1702
rect 25056 1426 25084 7398
rect 25148 2122 25176 9646
rect 25226 7712 25282 7721
rect 25226 7647 25282 7656
rect 25240 6390 25268 7647
rect 25332 7342 25360 9823
rect 25320 7336 25372 7342
rect 25320 7278 25372 7284
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 25424 4826 25452 9982
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25228 4616 25280 4622
rect 25228 4558 25280 4564
rect 25240 4457 25268 4558
rect 25226 4448 25282 4457
rect 25226 4383 25282 4392
rect 25148 2094 25268 2122
rect 25136 2032 25188 2038
rect 25136 1974 25188 1980
rect 25044 1420 25096 1426
rect 25044 1362 25096 1368
rect 24872 1278 25084 1306
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 25056 160 25084 1278
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24766 0 24822 54
rect 25042 0 25098 160
rect 25148 82 25176 1974
rect 25240 814 25268 2094
rect 25516 882 25544 12406
rect 25608 2417 25636 26846
rect 25686 25256 25742 25265
rect 25686 25191 25742 25200
rect 25700 12306 25728 25191
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 25686 5808 25742 5817
rect 25686 5743 25742 5752
rect 25700 5545 25728 5743
rect 25686 5536 25742 5545
rect 25686 5471 25742 5480
rect 25686 3224 25742 3233
rect 25792 3210 25820 41550
rect 25872 30728 25924 30734
rect 25872 30670 25924 30676
rect 25884 17241 25912 30670
rect 25870 17232 25926 17241
rect 25870 17167 25926 17176
rect 25742 3182 25820 3210
rect 25686 3159 25742 3168
rect 25594 2408 25650 2417
rect 25594 2343 25650 2352
rect 25596 2304 25648 2310
rect 25686 2272 25742 2281
rect 25648 2252 25686 2258
rect 25596 2246 25686 2252
rect 25608 2230 25686 2246
rect 25686 2207 25742 2216
rect 25596 1012 25648 1018
rect 25596 954 25648 960
rect 25504 876 25556 882
rect 25504 818 25556 824
rect 25228 808 25280 814
rect 25228 750 25280 756
rect 25608 160 25636 954
rect 25318 82 25374 160
rect 25148 54 25374 82
rect 25318 0 25374 54
rect 25594 0 25650 160
<< via2 >>
rect 294 36896 350 36952
rect 938 40160 994 40216
rect 662 40024 718 40080
rect 754 37848 810 37904
rect 754 34584 810 34640
rect 846 31728 902 31784
rect 570 29280 626 29336
rect 386 24656 442 24712
rect 754 28328 810 28384
rect 754 27784 810 27840
rect 754 23432 810 23488
rect 386 22208 442 22264
rect 294 20032 350 20088
rect 386 4256 442 4312
rect 938 29688 994 29744
rect 1214 38156 1216 38176
rect 1216 38156 1268 38176
rect 1268 38156 1270 38176
rect 1214 38120 1270 38156
rect 1214 33496 1270 33552
rect 1214 32408 1270 32464
rect 1122 32136 1178 32192
rect 1214 31864 1270 31920
rect 1490 42064 1546 42120
rect 1490 39480 1546 39536
rect 1398 39344 1454 39400
rect 1398 34856 1454 34912
rect 2226 39344 2282 39400
rect 1674 37848 1730 37904
rect 2226 38276 2282 38312
rect 2226 38256 2228 38276
rect 2228 38256 2280 38276
rect 2280 38256 2282 38276
rect 1766 36644 1822 36680
rect 1766 36624 1768 36644
rect 1768 36624 1820 36644
rect 1820 36624 1822 36644
rect 1674 36216 1730 36272
rect 1582 35400 1638 35456
rect 1490 32952 1546 33008
rect 1674 32836 1730 32872
rect 1674 32816 1676 32836
rect 1676 32816 1728 32836
rect 1728 32816 1730 32836
rect 1490 31864 1546 31920
rect 1398 31320 1454 31376
rect 1306 30776 1362 30832
rect 1306 29416 1362 29472
rect 1950 36488 2006 36544
rect 2318 36524 2320 36544
rect 2320 36524 2372 36544
rect 2372 36524 2374 36544
rect 2318 36488 2374 36524
rect 2226 36080 2282 36136
rect 2042 34604 2098 34640
rect 2042 34584 2044 34604
rect 2044 34584 2096 34604
rect 2096 34584 2098 34604
rect 1858 32408 1914 32464
rect 1490 30096 1546 30152
rect 1582 29416 1638 29472
rect 1490 28736 1546 28792
rect 3054 42608 3110 42664
rect 3923 43002 3979 43004
rect 4003 43002 4059 43004
rect 4083 43002 4139 43004
rect 4163 43002 4219 43004
rect 3923 42950 3969 43002
rect 3969 42950 3979 43002
rect 4003 42950 4033 43002
rect 4033 42950 4045 43002
rect 4045 42950 4059 43002
rect 4083 42950 4097 43002
rect 4097 42950 4109 43002
rect 4109 42950 4139 43002
rect 4163 42950 4173 43002
rect 4173 42950 4219 43002
rect 3923 42948 3979 42950
rect 4003 42948 4059 42950
rect 4083 42948 4139 42950
rect 4163 42948 4219 42950
rect 3923 41914 3979 41916
rect 4003 41914 4059 41916
rect 4083 41914 4139 41916
rect 4163 41914 4219 41916
rect 3923 41862 3969 41914
rect 3969 41862 3979 41914
rect 4003 41862 4033 41914
rect 4033 41862 4045 41914
rect 4045 41862 4059 41914
rect 4083 41862 4097 41914
rect 4097 41862 4109 41914
rect 4109 41862 4139 41914
rect 4163 41862 4173 41914
rect 4173 41862 4219 41914
rect 3923 41860 3979 41862
rect 4003 41860 4059 41862
rect 4083 41860 4139 41862
rect 4163 41860 4219 41862
rect 3422 41384 3478 41440
rect 4158 41540 4214 41576
rect 4158 41520 4160 41540
rect 4160 41520 4212 41540
rect 4212 41520 4214 41540
rect 3238 40024 3294 40080
rect 2778 38936 2834 38992
rect 3054 38392 3110 38448
rect 3054 38120 3110 38176
rect 2962 37440 3018 37496
rect 2778 37188 2834 37224
rect 2778 37168 2780 37188
rect 2780 37168 2832 37188
rect 2832 37168 2834 37188
rect 2778 35672 2834 35728
rect 3146 36760 3202 36816
rect 2686 33904 2742 33960
rect 2686 33768 2742 33824
rect 2502 32544 2558 32600
rect 2134 30096 2190 30152
rect 1214 26424 1270 26480
rect 1122 26288 1178 26344
rect 1306 25336 1362 25392
rect 1214 25200 1270 25256
rect 938 24112 994 24168
rect 1122 24520 1178 24576
rect 1030 23704 1086 23760
rect 1766 27376 1822 27432
rect 1582 26832 1638 26888
rect 1766 26832 1822 26888
rect 1582 25744 1638 25800
rect 1398 23976 1454 24032
rect 1306 23568 1362 23624
rect 1950 28600 2006 28656
rect 1858 25336 1914 25392
rect 1858 25200 1914 25256
rect 2042 27648 2098 27704
rect 2042 26016 2098 26072
rect 2410 30776 2466 30832
rect 2318 28328 2374 28384
rect 2318 27512 2374 27568
rect 2226 26968 2282 27024
rect 3422 37984 3478 38040
rect 3606 35980 3608 36000
rect 3608 35980 3660 36000
rect 3660 35980 3662 36000
rect 3606 35944 3662 35980
rect 3422 34040 3478 34096
rect 2870 33224 2926 33280
rect 2778 32680 2834 32736
rect 2778 31048 2834 31104
rect 2594 30676 2596 30696
rect 2596 30676 2648 30696
rect 2648 30676 2650 30696
rect 2594 30640 2650 30676
rect 2594 28500 2596 28520
rect 2596 28500 2648 28520
rect 2648 28500 2650 28520
rect 2594 28464 2650 28500
rect 3146 30368 3202 30424
rect 2686 27512 2742 27568
rect 2594 26560 2650 26616
rect 1674 24248 1730 24304
rect 1766 23704 1822 23760
rect 1306 22888 1362 22944
rect 754 20168 810 20224
rect 846 19896 902 19952
rect 662 12552 718 12608
rect 1030 17040 1086 17096
rect 1030 16904 1086 16960
rect 846 9288 902 9344
rect 1030 9288 1086 9344
rect 1030 9016 1086 9072
rect 1030 6568 1086 6624
rect 938 1944 994 2000
rect 1306 21800 1362 21856
rect 1214 21528 1270 21584
rect 1582 23160 1638 23216
rect 1490 22344 1546 22400
rect 2134 24792 2190 24848
rect 2134 23432 2190 23488
rect 1766 21956 1822 21992
rect 1766 21936 1768 21956
rect 1768 21936 1820 21956
rect 1820 21936 1822 21956
rect 1214 21256 1270 21312
rect 1306 20984 1362 21040
rect 1214 20848 1270 20904
rect 1306 20712 1362 20768
rect 1398 20440 1454 20496
rect 1306 19624 1362 19680
rect 1674 21664 1730 21720
rect 1858 20848 1914 20904
rect 1582 19760 1638 19816
rect 1766 19352 1822 19408
rect 1674 19252 1676 19272
rect 1676 19252 1728 19272
rect 1728 19252 1730 19272
rect 1674 19216 1730 19252
rect 1398 18808 1454 18864
rect 1306 18264 1362 18320
rect 1214 17992 1270 18048
rect 1490 18536 1546 18592
rect 1582 17720 1638 17776
rect 1214 13096 1270 13152
rect 1398 13912 1454 13968
rect 1766 17448 1822 17504
rect 2778 26832 2834 26888
rect 2962 27376 3018 27432
rect 2962 27276 2964 27296
rect 2964 27276 3016 27296
rect 3016 27276 3018 27296
rect 2962 27240 3018 27276
rect 3238 29280 3294 29336
rect 3330 29144 3386 29200
rect 3146 28056 3202 28112
rect 3606 34040 3662 34096
rect 3923 40826 3979 40828
rect 4003 40826 4059 40828
rect 4083 40826 4139 40828
rect 4163 40826 4219 40828
rect 3923 40774 3969 40826
rect 3969 40774 3979 40826
rect 4003 40774 4033 40826
rect 4033 40774 4045 40826
rect 4045 40774 4059 40826
rect 4083 40774 4097 40826
rect 4097 40774 4109 40826
rect 4109 40774 4139 40826
rect 4163 40774 4173 40826
rect 4173 40774 4219 40826
rect 3923 40772 3979 40774
rect 4003 40772 4059 40774
rect 4083 40772 4139 40774
rect 4163 40772 4219 40774
rect 3790 40432 3846 40488
rect 4618 41556 4620 41576
rect 4620 41556 4672 41576
rect 4672 41556 4674 41576
rect 4618 41520 4674 41556
rect 4250 40160 4306 40216
rect 3923 39738 3979 39740
rect 4003 39738 4059 39740
rect 4083 39738 4139 39740
rect 4163 39738 4219 39740
rect 3923 39686 3969 39738
rect 3969 39686 3979 39738
rect 4003 39686 4033 39738
rect 4033 39686 4045 39738
rect 4045 39686 4059 39738
rect 4083 39686 4097 39738
rect 4097 39686 4109 39738
rect 4109 39686 4139 39738
rect 4163 39686 4173 39738
rect 4173 39686 4219 39738
rect 3923 39684 3979 39686
rect 4003 39684 4059 39686
rect 4083 39684 4139 39686
rect 4163 39684 4219 39686
rect 3882 38836 3884 38856
rect 3884 38836 3936 38856
rect 3936 38836 3938 38856
rect 3882 38800 3938 38836
rect 3923 38650 3979 38652
rect 4003 38650 4059 38652
rect 4083 38650 4139 38652
rect 4163 38650 4219 38652
rect 3923 38598 3969 38650
rect 3969 38598 3979 38650
rect 4003 38598 4033 38650
rect 4033 38598 4045 38650
rect 4045 38598 4059 38650
rect 4083 38598 4097 38650
rect 4097 38598 4109 38650
rect 4109 38598 4139 38650
rect 4163 38598 4173 38650
rect 4173 38598 4219 38650
rect 3923 38596 3979 38598
rect 4003 38596 4059 38598
rect 4083 38596 4139 38598
rect 4163 38596 4219 38598
rect 3923 37562 3979 37564
rect 4003 37562 4059 37564
rect 4083 37562 4139 37564
rect 4163 37562 4219 37564
rect 3923 37510 3969 37562
rect 3969 37510 3979 37562
rect 4003 37510 4033 37562
rect 4033 37510 4045 37562
rect 4045 37510 4059 37562
rect 4083 37510 4097 37562
rect 4097 37510 4109 37562
rect 4109 37510 4139 37562
rect 4163 37510 4173 37562
rect 4173 37510 4219 37562
rect 3923 37508 3979 37510
rect 4003 37508 4059 37510
rect 4083 37508 4139 37510
rect 4163 37508 4219 37510
rect 3882 37032 3938 37088
rect 4066 36760 4122 36816
rect 3790 36488 3846 36544
rect 3923 36474 3979 36476
rect 4003 36474 4059 36476
rect 4083 36474 4139 36476
rect 4163 36474 4219 36476
rect 3923 36422 3969 36474
rect 3969 36422 3979 36474
rect 4003 36422 4033 36474
rect 4033 36422 4045 36474
rect 4045 36422 4059 36474
rect 4083 36422 4097 36474
rect 4097 36422 4109 36474
rect 4109 36422 4139 36474
rect 4163 36422 4173 36474
rect 4173 36422 4219 36474
rect 3923 36420 3979 36422
rect 4003 36420 4059 36422
rect 4083 36420 4139 36422
rect 4163 36420 4219 36422
rect 4066 35944 4122 36000
rect 3923 35386 3979 35388
rect 4003 35386 4059 35388
rect 4083 35386 4139 35388
rect 4163 35386 4219 35388
rect 3923 35334 3969 35386
rect 3969 35334 3979 35386
rect 4003 35334 4033 35386
rect 4033 35334 4045 35386
rect 4045 35334 4059 35386
rect 4083 35334 4097 35386
rect 4097 35334 4109 35386
rect 4109 35334 4139 35386
rect 4163 35334 4173 35386
rect 4173 35334 4219 35386
rect 3923 35332 3979 35334
rect 4003 35332 4059 35334
rect 4083 35332 4139 35334
rect 4163 35332 4219 35334
rect 3790 35128 3846 35184
rect 4342 36896 4398 36952
rect 4250 34856 4306 34912
rect 4066 34448 4122 34504
rect 3923 34298 3979 34300
rect 4003 34298 4059 34300
rect 4083 34298 4139 34300
rect 4163 34298 4219 34300
rect 3923 34246 3969 34298
rect 3969 34246 3979 34298
rect 4003 34246 4033 34298
rect 4033 34246 4045 34298
rect 4045 34246 4059 34298
rect 4083 34246 4097 34298
rect 4097 34246 4109 34298
rect 4109 34246 4139 34298
rect 4163 34246 4173 34298
rect 4173 34246 4219 34298
rect 3923 34244 3979 34246
rect 4003 34244 4059 34246
rect 4083 34244 4139 34246
rect 4163 34244 4219 34246
rect 3923 33210 3979 33212
rect 4003 33210 4059 33212
rect 4083 33210 4139 33212
rect 4163 33210 4219 33212
rect 3923 33158 3969 33210
rect 3969 33158 3979 33210
rect 4003 33158 4033 33210
rect 4033 33158 4045 33210
rect 4045 33158 4059 33210
rect 4083 33158 4097 33210
rect 4097 33158 4109 33210
rect 4109 33158 4139 33210
rect 4163 33158 4173 33210
rect 4173 33158 4219 33210
rect 3923 33156 3979 33158
rect 4003 33156 4059 33158
rect 4083 33156 4139 33158
rect 4163 33156 4219 33158
rect 4342 33632 4398 33688
rect 3923 32122 3979 32124
rect 4003 32122 4059 32124
rect 4083 32122 4139 32124
rect 4163 32122 4219 32124
rect 3923 32070 3969 32122
rect 3969 32070 3979 32122
rect 4003 32070 4033 32122
rect 4033 32070 4045 32122
rect 4045 32070 4059 32122
rect 4083 32070 4097 32122
rect 4097 32070 4109 32122
rect 4109 32070 4139 32122
rect 4163 32070 4173 32122
rect 4173 32070 4219 32122
rect 3923 32068 3979 32070
rect 4003 32068 4059 32070
rect 4083 32068 4139 32070
rect 4163 32068 4219 32070
rect 3790 31592 3846 31648
rect 3923 31034 3979 31036
rect 4003 31034 4059 31036
rect 4083 31034 4139 31036
rect 4163 31034 4219 31036
rect 3923 30982 3969 31034
rect 3969 30982 3979 31034
rect 4003 30982 4033 31034
rect 4033 30982 4045 31034
rect 4045 30982 4059 31034
rect 4083 30982 4097 31034
rect 4097 30982 4109 31034
rect 4109 30982 4139 31034
rect 4163 30982 4173 31034
rect 4173 30982 4219 31034
rect 3923 30980 3979 30982
rect 4003 30980 4059 30982
rect 4083 30980 4139 30982
rect 4163 30980 4219 30982
rect 3698 30504 3754 30560
rect 3882 30368 3938 30424
rect 3790 30232 3846 30288
rect 4710 38664 4766 38720
rect 4894 37304 4950 37360
rect 4618 32308 4620 32328
rect 4620 32308 4672 32328
rect 4672 32308 4674 32328
rect 4618 32272 4674 32308
rect 4434 31456 4490 31512
rect 4434 31184 4490 31240
rect 3923 29946 3979 29948
rect 4003 29946 4059 29948
rect 4083 29946 4139 29948
rect 4163 29946 4219 29948
rect 3923 29894 3969 29946
rect 3969 29894 3979 29946
rect 4003 29894 4033 29946
rect 4033 29894 4045 29946
rect 4045 29894 4059 29946
rect 4083 29894 4097 29946
rect 4097 29894 4109 29946
rect 4109 29894 4139 29946
rect 4163 29894 4173 29946
rect 4173 29894 4219 29946
rect 3923 29892 3979 29894
rect 4003 29892 4059 29894
rect 4083 29892 4139 29894
rect 4163 29892 4219 29894
rect 3606 28872 3662 28928
rect 3923 28858 3979 28860
rect 4003 28858 4059 28860
rect 4083 28858 4139 28860
rect 4163 28858 4219 28860
rect 3923 28806 3969 28858
rect 3969 28806 3979 28858
rect 4003 28806 4033 28858
rect 4033 28806 4045 28858
rect 4045 28806 4059 28858
rect 4083 28806 4097 28858
rect 4097 28806 4109 28858
rect 4109 28806 4139 28858
rect 4163 28806 4173 28858
rect 4173 28806 4219 28858
rect 3923 28804 3979 28806
rect 4003 28804 4059 28806
rect 4083 28804 4139 28806
rect 4163 28804 4219 28806
rect 4158 28500 4160 28520
rect 4160 28500 4212 28520
rect 4212 28500 4214 28520
rect 2778 26016 2834 26072
rect 2870 25608 2926 25664
rect 2870 24656 2926 24712
rect 2778 23840 2834 23896
rect 2870 22616 2926 22672
rect 2134 21392 2190 21448
rect 2594 20984 2650 21040
rect 2318 20712 2374 20768
rect 2042 20440 2098 20496
rect 1950 19352 2006 19408
rect 1858 16768 1914 16824
rect 1674 15816 1730 15872
rect 1858 14592 1914 14648
rect 1766 14320 1822 14376
rect 1766 14184 1822 14240
rect 1398 12008 1454 12064
rect 1214 9560 1270 9616
rect 1950 14184 2006 14240
rect 1858 11464 1914 11520
rect 1674 10920 1730 10976
rect 1582 9424 1638 9480
rect 1766 9832 1822 9888
rect 1582 8744 1638 8800
rect 1306 8472 1362 8528
rect 1398 8200 1454 8256
rect 1214 6840 1270 6896
rect 1306 6296 1362 6352
rect 1306 5752 1362 5808
rect 1398 4936 1454 4992
rect 1674 7656 1730 7712
rect 1582 6024 1638 6080
rect 3146 22616 3202 22672
rect 2962 20168 3018 20224
rect 3054 19760 3110 19816
rect 2318 15136 2374 15192
rect 2594 18400 2650 18456
rect 2594 18264 2650 18320
rect 2686 16396 2688 16416
rect 2688 16396 2740 16416
rect 2740 16396 2742 16416
rect 2686 16360 2742 16396
rect 2870 16632 2926 16688
rect 3054 16088 3110 16144
rect 3054 15544 3110 15600
rect 3238 22072 3294 22128
rect 3238 21800 3294 21856
rect 4158 28464 4214 28500
rect 4066 28056 4122 28112
rect 4250 27920 4306 27976
rect 3923 27770 3979 27772
rect 4003 27770 4059 27772
rect 4083 27770 4139 27772
rect 4163 27770 4219 27772
rect 3923 27718 3969 27770
rect 3969 27718 3979 27770
rect 4003 27718 4033 27770
rect 4033 27718 4045 27770
rect 4045 27718 4059 27770
rect 4083 27718 4097 27770
rect 4097 27718 4109 27770
rect 4109 27718 4139 27770
rect 4163 27718 4173 27770
rect 4173 27718 4219 27770
rect 3923 27716 3979 27718
rect 4003 27716 4059 27718
rect 4083 27716 4139 27718
rect 4163 27716 4219 27718
rect 3422 25880 3478 25936
rect 3923 26682 3979 26684
rect 4003 26682 4059 26684
rect 4083 26682 4139 26684
rect 4163 26682 4219 26684
rect 3923 26630 3969 26682
rect 3969 26630 3979 26682
rect 4003 26630 4033 26682
rect 4033 26630 4045 26682
rect 4045 26630 4059 26682
rect 4083 26630 4097 26682
rect 4097 26630 4109 26682
rect 4109 26630 4139 26682
rect 4163 26630 4173 26682
rect 4173 26630 4219 26682
rect 3923 26628 3979 26630
rect 4003 26628 4059 26630
rect 4083 26628 4139 26630
rect 4163 26628 4219 26630
rect 3790 26152 3846 26208
rect 4434 27784 4490 27840
rect 3923 25594 3979 25596
rect 4003 25594 4059 25596
rect 4083 25594 4139 25596
rect 4163 25594 4219 25596
rect 3923 25542 3969 25594
rect 3969 25542 3979 25594
rect 4003 25542 4033 25594
rect 4033 25542 4045 25594
rect 4045 25542 4059 25594
rect 4083 25542 4097 25594
rect 4097 25542 4109 25594
rect 4109 25542 4139 25594
rect 4163 25542 4173 25594
rect 4173 25542 4219 25594
rect 3923 25540 3979 25542
rect 4003 25540 4059 25542
rect 4083 25540 4139 25542
rect 4163 25540 4219 25542
rect 3923 24506 3979 24508
rect 4003 24506 4059 24508
rect 4083 24506 4139 24508
rect 4163 24506 4219 24508
rect 3923 24454 3969 24506
rect 3969 24454 3979 24506
rect 4003 24454 4033 24506
rect 4033 24454 4045 24506
rect 4045 24454 4059 24506
rect 4083 24454 4097 24506
rect 4097 24454 4109 24506
rect 4109 24454 4139 24506
rect 4163 24454 4173 24506
rect 4173 24454 4219 24506
rect 3923 24452 3979 24454
rect 4003 24452 4059 24454
rect 4083 24452 4139 24454
rect 4163 24452 4219 24454
rect 3422 21664 3478 21720
rect 4066 24112 4122 24168
rect 3923 23418 3979 23420
rect 4003 23418 4059 23420
rect 4083 23418 4139 23420
rect 4163 23418 4219 23420
rect 3923 23366 3969 23418
rect 3969 23366 3979 23418
rect 4003 23366 4033 23418
rect 4033 23366 4045 23418
rect 4045 23366 4059 23418
rect 4083 23366 4097 23418
rect 4097 23366 4109 23418
rect 4109 23366 4139 23418
rect 4163 23366 4173 23418
rect 4173 23366 4219 23418
rect 3923 23364 3979 23366
rect 4003 23364 4059 23366
rect 4083 23364 4139 23366
rect 4163 23364 4219 23366
rect 3974 22888 4030 22944
rect 4710 29688 4766 29744
rect 4986 34856 5042 34912
rect 5078 34604 5134 34640
rect 5078 34584 5080 34604
rect 5080 34584 5132 34604
rect 5132 34584 5134 34604
rect 4894 31048 4950 31104
rect 4894 30368 4950 30424
rect 6890 43546 6946 43548
rect 6970 43546 7026 43548
rect 7050 43546 7106 43548
rect 7130 43546 7186 43548
rect 6890 43494 6936 43546
rect 6936 43494 6946 43546
rect 6970 43494 7000 43546
rect 7000 43494 7012 43546
rect 7012 43494 7026 43546
rect 7050 43494 7064 43546
rect 7064 43494 7076 43546
rect 7076 43494 7106 43546
rect 7130 43494 7140 43546
rect 7140 43494 7186 43546
rect 6890 43492 6946 43494
rect 6970 43492 7026 43494
rect 7050 43492 7106 43494
rect 7130 43492 7186 43494
rect 6890 42458 6946 42460
rect 6970 42458 7026 42460
rect 7050 42458 7106 42460
rect 7130 42458 7186 42460
rect 6890 42406 6936 42458
rect 6936 42406 6946 42458
rect 6970 42406 7000 42458
rect 7000 42406 7012 42458
rect 7012 42406 7026 42458
rect 7050 42406 7064 42458
rect 7064 42406 7076 42458
rect 7076 42406 7106 42458
rect 7130 42406 7140 42458
rect 7140 42406 7186 42458
rect 6890 42404 6946 42406
rect 6970 42404 7026 42406
rect 7050 42404 7106 42406
rect 7130 42404 7186 42406
rect 6182 41792 6238 41848
rect 6550 41656 6606 41712
rect 6734 41556 6736 41576
rect 6736 41556 6788 41576
rect 6788 41556 6790 41576
rect 6734 41520 6790 41556
rect 7378 42064 7434 42120
rect 7654 41792 7710 41848
rect 5262 39072 5318 39128
rect 5630 38256 5686 38312
rect 5814 40568 5870 40624
rect 5814 37848 5870 37904
rect 5538 37304 5594 37360
rect 6890 41370 6946 41372
rect 6970 41370 7026 41372
rect 7050 41370 7106 41372
rect 7130 41370 7186 41372
rect 6890 41318 6936 41370
rect 6936 41318 6946 41370
rect 6970 41318 7000 41370
rect 7000 41318 7012 41370
rect 7012 41318 7026 41370
rect 7050 41318 7064 41370
rect 7064 41318 7076 41370
rect 7076 41318 7106 41370
rect 7130 41318 7140 41370
rect 7140 41318 7186 41370
rect 6890 41316 6946 41318
rect 6970 41316 7026 41318
rect 7050 41316 7106 41318
rect 7130 41316 7186 41318
rect 6826 40468 6828 40488
rect 6828 40468 6880 40488
rect 6880 40468 6882 40488
rect 6826 40432 6882 40468
rect 6890 40282 6946 40284
rect 6970 40282 7026 40284
rect 7050 40282 7106 40284
rect 7130 40282 7186 40284
rect 6890 40230 6936 40282
rect 6936 40230 6946 40282
rect 6970 40230 7000 40282
rect 7000 40230 7012 40282
rect 7012 40230 7026 40282
rect 7050 40230 7064 40282
rect 7064 40230 7076 40282
rect 7076 40230 7106 40282
rect 7130 40230 7140 40282
rect 7140 40230 7186 40282
rect 6890 40228 6946 40230
rect 6970 40228 7026 40230
rect 7050 40228 7106 40230
rect 7130 40228 7186 40230
rect 5446 35164 5448 35184
rect 5448 35164 5500 35184
rect 5500 35164 5502 35184
rect 5446 35128 5502 35164
rect 5630 35536 5686 35592
rect 5538 34448 5594 34504
rect 5906 34992 5962 35048
rect 5906 31728 5962 31784
rect 6182 33904 6238 33960
rect 6274 33224 6330 33280
rect 5446 31356 5448 31376
rect 5448 31356 5500 31376
rect 5500 31356 5502 31376
rect 5446 31320 5502 31356
rect 5446 30776 5502 30832
rect 4986 28736 5042 28792
rect 4986 28464 5042 28520
rect 3923 22330 3979 22332
rect 4003 22330 4059 22332
rect 4083 22330 4139 22332
rect 4163 22330 4219 22332
rect 3923 22278 3969 22330
rect 3969 22278 3979 22330
rect 4003 22278 4033 22330
rect 4033 22278 4045 22330
rect 4045 22278 4059 22330
rect 4083 22278 4097 22330
rect 4097 22278 4109 22330
rect 4109 22278 4139 22330
rect 4163 22278 4173 22330
rect 4173 22278 4219 22330
rect 3923 22276 3979 22278
rect 4003 22276 4059 22278
rect 4083 22276 4139 22278
rect 4163 22276 4219 22278
rect 3974 22072 4030 22128
rect 3923 21242 3979 21244
rect 4003 21242 4059 21244
rect 4083 21242 4139 21244
rect 4163 21242 4219 21244
rect 3923 21190 3969 21242
rect 3969 21190 3979 21242
rect 4003 21190 4033 21242
rect 4033 21190 4045 21242
rect 4045 21190 4059 21242
rect 4083 21190 4097 21242
rect 4097 21190 4109 21242
rect 4109 21190 4139 21242
rect 4163 21190 4173 21242
rect 4173 21190 4219 21242
rect 3923 21188 3979 21190
rect 4003 21188 4059 21190
rect 4083 21188 4139 21190
rect 4163 21188 4219 21190
rect 4158 20712 4214 20768
rect 3330 19080 3386 19136
rect 3923 20154 3979 20156
rect 4003 20154 4059 20156
rect 4083 20154 4139 20156
rect 4163 20154 4219 20156
rect 3923 20102 3969 20154
rect 3969 20102 3979 20154
rect 4003 20102 4033 20154
rect 4033 20102 4045 20154
rect 4045 20102 4059 20154
rect 4083 20102 4097 20154
rect 4097 20102 4109 20154
rect 4109 20102 4139 20154
rect 4163 20102 4173 20154
rect 4173 20102 4219 20154
rect 3923 20100 3979 20102
rect 4003 20100 4059 20102
rect 4083 20100 4139 20102
rect 4163 20100 4219 20102
rect 3923 19066 3979 19068
rect 4003 19066 4059 19068
rect 4083 19066 4139 19068
rect 4163 19066 4219 19068
rect 3923 19014 3969 19066
rect 3969 19014 3979 19066
rect 4003 19014 4033 19066
rect 4033 19014 4045 19066
rect 4045 19014 4059 19066
rect 4083 19014 4097 19066
rect 4097 19014 4109 19066
rect 4109 19014 4139 19066
rect 4163 19014 4173 19066
rect 4173 19014 4219 19066
rect 3923 19012 3979 19014
rect 4003 19012 4059 19014
rect 4083 19012 4139 19014
rect 4163 19012 4219 19014
rect 3974 18808 4030 18864
rect 3974 18164 3976 18184
rect 3976 18164 4028 18184
rect 4028 18164 4030 18184
rect 3974 18128 4030 18164
rect 4158 18400 4214 18456
rect 3923 17978 3979 17980
rect 4003 17978 4059 17980
rect 4083 17978 4139 17980
rect 4163 17978 4219 17980
rect 3923 17926 3969 17978
rect 3969 17926 3979 17978
rect 4003 17926 4033 17978
rect 4033 17926 4045 17978
rect 4045 17926 4059 17978
rect 4083 17926 4097 17978
rect 4097 17926 4109 17978
rect 4109 17926 4139 17978
rect 4163 17926 4173 17978
rect 4173 17926 4219 17978
rect 3923 17924 3979 17926
rect 4003 17924 4059 17926
rect 4083 17924 4139 17926
rect 4163 17924 4219 17926
rect 3330 17176 3386 17232
rect 3330 16224 3386 16280
rect 2778 14456 2834 14512
rect 2318 12824 2374 12880
rect 2042 11056 2098 11112
rect 2042 9968 2098 10024
rect 2042 9288 2098 9344
rect 1766 7384 1822 7440
rect 1766 5344 1822 5400
rect 1858 3032 1914 3088
rect 1122 2216 1178 2272
rect 2134 7828 2136 7848
rect 2136 7828 2188 7848
rect 2188 7828 2190 7848
rect 2134 7792 2190 7828
rect 2318 8336 2374 8392
rect 3330 13232 3386 13288
rect 2962 12144 3018 12200
rect 2870 12008 2926 12064
rect 2778 11872 2834 11928
rect 2686 9968 2742 10024
rect 2594 6724 2650 6760
rect 2594 6704 2596 6724
rect 2596 6704 2648 6724
rect 2648 6704 2650 6724
rect 2134 4392 2190 4448
rect 2318 5652 2320 5672
rect 2320 5652 2372 5672
rect 2372 5652 2374 5672
rect 2318 5616 2374 5652
rect 2134 2644 2190 2680
rect 2134 2624 2136 2644
rect 2136 2624 2188 2644
rect 2188 2624 2190 2644
rect 3146 11736 3202 11792
rect 3330 11600 3386 11656
rect 3238 11464 3294 11520
rect 3054 10104 3110 10160
rect 2870 5208 2926 5264
rect 3974 17720 4030 17776
rect 3923 16890 3979 16892
rect 4003 16890 4059 16892
rect 4083 16890 4139 16892
rect 4163 16890 4219 16892
rect 3923 16838 3969 16890
rect 3969 16838 3979 16890
rect 4003 16838 4033 16890
rect 4033 16838 4045 16890
rect 4045 16838 4059 16890
rect 4083 16838 4097 16890
rect 4097 16838 4109 16890
rect 4109 16838 4139 16890
rect 4163 16838 4173 16890
rect 4173 16838 4219 16890
rect 3923 16836 3979 16838
rect 4003 16836 4059 16838
rect 4083 16836 4139 16838
rect 4163 16836 4219 16838
rect 3514 15544 3570 15600
rect 3923 15802 3979 15804
rect 4003 15802 4059 15804
rect 4083 15802 4139 15804
rect 4163 15802 4219 15804
rect 3923 15750 3969 15802
rect 3969 15750 3979 15802
rect 4003 15750 4033 15802
rect 4033 15750 4045 15802
rect 4045 15750 4059 15802
rect 4083 15750 4097 15802
rect 4097 15750 4109 15802
rect 4109 15750 4139 15802
rect 4163 15750 4173 15802
rect 4173 15750 4219 15802
rect 3923 15748 3979 15750
rect 4003 15748 4059 15750
rect 4083 15748 4139 15750
rect 4163 15748 4219 15750
rect 3974 15408 4030 15464
rect 3923 14714 3979 14716
rect 4003 14714 4059 14716
rect 4083 14714 4139 14716
rect 4163 14714 4219 14716
rect 3923 14662 3969 14714
rect 3969 14662 3979 14714
rect 4003 14662 4033 14714
rect 4033 14662 4045 14714
rect 4045 14662 4059 14714
rect 4083 14662 4097 14714
rect 4097 14662 4109 14714
rect 4109 14662 4139 14714
rect 4163 14662 4173 14714
rect 4173 14662 4219 14714
rect 3923 14660 3979 14662
rect 4003 14660 4059 14662
rect 4083 14660 4139 14662
rect 4163 14660 4219 14662
rect 4434 21120 4490 21176
rect 4342 16088 4398 16144
rect 4618 22752 4674 22808
rect 4618 22208 4674 22264
rect 4986 25608 5042 25664
rect 5170 29008 5226 29064
rect 5630 29008 5686 29064
rect 5538 28192 5594 28248
rect 5262 28056 5318 28112
rect 5630 27956 5632 27976
rect 5632 27956 5684 27976
rect 5684 27956 5686 27976
rect 5630 27920 5686 27956
rect 5078 24248 5134 24304
rect 4986 23432 5042 23488
rect 4618 21528 4674 21584
rect 4618 20032 4674 20088
rect 4894 21256 4950 21312
rect 4894 20848 4950 20904
rect 4250 14456 4306 14512
rect 5262 22072 5318 22128
rect 5078 21120 5134 21176
rect 5538 26152 5594 26208
rect 5446 23160 5502 23216
rect 5722 24656 5778 24712
rect 5630 24248 5686 24304
rect 6182 30912 6238 30968
rect 6090 29552 6146 29608
rect 6090 29008 6146 29064
rect 6090 27920 6146 27976
rect 6890 39194 6946 39196
rect 6970 39194 7026 39196
rect 7050 39194 7106 39196
rect 7130 39194 7186 39196
rect 6890 39142 6936 39194
rect 6936 39142 6946 39194
rect 6970 39142 7000 39194
rect 7000 39142 7012 39194
rect 7012 39142 7026 39194
rect 7050 39142 7064 39194
rect 7064 39142 7076 39194
rect 7076 39142 7106 39194
rect 7130 39142 7140 39194
rect 7140 39142 7186 39194
rect 6890 39140 6946 39142
rect 6970 39140 7026 39142
rect 7050 39140 7106 39142
rect 7130 39140 7186 39142
rect 6890 38106 6946 38108
rect 6970 38106 7026 38108
rect 7050 38106 7106 38108
rect 7130 38106 7186 38108
rect 6890 38054 6936 38106
rect 6936 38054 6946 38106
rect 6970 38054 7000 38106
rect 7000 38054 7012 38106
rect 7012 38054 7026 38106
rect 7050 38054 7064 38106
rect 7064 38054 7076 38106
rect 7076 38054 7106 38106
rect 7130 38054 7140 38106
rect 7140 38054 7186 38106
rect 6890 38052 6946 38054
rect 6970 38052 7026 38054
rect 7050 38052 7106 38054
rect 7130 38052 7186 38054
rect 6890 37018 6946 37020
rect 6970 37018 7026 37020
rect 7050 37018 7106 37020
rect 7130 37018 7186 37020
rect 6890 36966 6936 37018
rect 6936 36966 6946 37018
rect 6970 36966 7000 37018
rect 7000 36966 7012 37018
rect 7012 36966 7026 37018
rect 7050 36966 7064 37018
rect 7064 36966 7076 37018
rect 7076 36966 7106 37018
rect 7130 36966 7140 37018
rect 7140 36966 7186 37018
rect 6890 36964 6946 36966
rect 6970 36964 7026 36966
rect 7050 36964 7106 36966
rect 7130 36964 7186 36966
rect 6890 35930 6946 35932
rect 6970 35930 7026 35932
rect 7050 35930 7106 35932
rect 7130 35930 7186 35932
rect 6890 35878 6936 35930
rect 6936 35878 6946 35930
rect 6970 35878 7000 35930
rect 7000 35878 7012 35930
rect 7012 35878 7026 35930
rect 7050 35878 7064 35930
rect 7064 35878 7076 35930
rect 7076 35878 7106 35930
rect 7130 35878 7140 35930
rect 7140 35878 7186 35930
rect 6890 35876 6946 35878
rect 6970 35876 7026 35878
rect 7050 35876 7106 35878
rect 7130 35876 7186 35878
rect 6890 34842 6946 34844
rect 6970 34842 7026 34844
rect 7050 34842 7106 34844
rect 7130 34842 7186 34844
rect 6890 34790 6936 34842
rect 6936 34790 6946 34842
rect 6970 34790 7000 34842
rect 7000 34790 7012 34842
rect 7012 34790 7026 34842
rect 7050 34790 7064 34842
rect 7064 34790 7076 34842
rect 7076 34790 7106 34842
rect 7130 34790 7140 34842
rect 7140 34790 7186 34842
rect 6890 34788 6946 34790
rect 6970 34788 7026 34790
rect 7050 34788 7106 34790
rect 7130 34788 7186 34790
rect 6890 33754 6946 33756
rect 6970 33754 7026 33756
rect 7050 33754 7106 33756
rect 7130 33754 7186 33756
rect 6890 33702 6936 33754
rect 6936 33702 6946 33754
rect 6970 33702 7000 33754
rect 7000 33702 7012 33754
rect 7012 33702 7026 33754
rect 7050 33702 7064 33754
rect 7064 33702 7076 33754
rect 7076 33702 7106 33754
rect 7130 33702 7140 33754
rect 7140 33702 7186 33754
rect 6890 33700 6946 33702
rect 6970 33700 7026 33702
rect 7050 33700 7106 33702
rect 7130 33700 7186 33702
rect 6642 32544 6698 32600
rect 6918 33360 6974 33416
rect 7194 33396 7196 33416
rect 7196 33396 7248 33416
rect 7248 33396 7250 33416
rect 7194 33360 7250 33396
rect 6890 32666 6946 32668
rect 6970 32666 7026 32668
rect 7050 32666 7106 32668
rect 7130 32666 7186 32668
rect 6890 32614 6936 32666
rect 6936 32614 6946 32666
rect 6970 32614 7000 32666
rect 7000 32614 7012 32666
rect 7012 32614 7026 32666
rect 7050 32614 7064 32666
rect 7064 32614 7076 32666
rect 7076 32614 7106 32666
rect 7130 32614 7140 32666
rect 7140 32614 7186 32666
rect 6890 32612 6946 32614
rect 6970 32612 7026 32614
rect 7050 32612 7106 32614
rect 7130 32612 7186 32614
rect 6642 31864 6698 31920
rect 6458 29416 6514 29472
rect 5354 19216 5410 19272
rect 5354 19116 5356 19136
rect 5356 19116 5408 19136
rect 5408 19116 5410 19136
rect 5354 19080 5410 19116
rect 4986 18128 5042 18184
rect 5170 16904 5226 16960
rect 4618 15156 4674 15192
rect 4618 15136 4620 15156
rect 4620 15136 4672 15156
rect 4672 15136 4674 15156
rect 3514 12960 3570 13016
rect 3514 11756 3570 11792
rect 3514 11736 3516 11756
rect 3516 11736 3568 11756
rect 3568 11736 3570 11756
rect 3790 13676 3792 13696
rect 3792 13676 3844 13696
rect 3844 13676 3846 13696
rect 3790 13640 3846 13676
rect 3923 13626 3979 13628
rect 4003 13626 4059 13628
rect 4083 13626 4139 13628
rect 4163 13626 4219 13628
rect 3923 13574 3969 13626
rect 3969 13574 3979 13626
rect 4003 13574 4033 13626
rect 4033 13574 4045 13626
rect 4045 13574 4059 13626
rect 4083 13574 4097 13626
rect 4097 13574 4109 13626
rect 4109 13574 4139 13626
rect 4163 13574 4173 13626
rect 4173 13574 4219 13626
rect 3923 13572 3979 13574
rect 4003 13572 4059 13574
rect 4083 13572 4139 13574
rect 4163 13572 4219 13574
rect 3790 13388 3846 13424
rect 3790 13368 3792 13388
rect 3792 13368 3844 13388
rect 3844 13368 3846 13388
rect 4066 13268 4068 13288
rect 4068 13268 4120 13288
rect 4120 13268 4122 13288
rect 4066 13232 4122 13268
rect 3882 12860 3884 12880
rect 3884 12860 3936 12880
rect 3936 12860 3938 12880
rect 3882 12824 3938 12860
rect 4066 12724 4068 12744
rect 4068 12724 4120 12744
rect 4120 12724 4122 12744
rect 4066 12688 4122 12724
rect 3923 12538 3979 12540
rect 4003 12538 4059 12540
rect 4083 12538 4139 12540
rect 4163 12538 4219 12540
rect 3923 12486 3969 12538
rect 3969 12486 3979 12538
rect 4003 12486 4033 12538
rect 4033 12486 4045 12538
rect 4045 12486 4059 12538
rect 4083 12486 4097 12538
rect 4097 12486 4109 12538
rect 4109 12486 4139 12538
rect 4163 12486 4173 12538
rect 4173 12486 4219 12538
rect 3923 12484 3979 12486
rect 4003 12484 4059 12486
rect 4083 12484 4139 12486
rect 4163 12484 4219 12486
rect 3698 12280 3754 12336
rect 3606 11464 3662 11520
rect 3606 11192 3662 11248
rect 3330 10376 3386 10432
rect 3330 9560 3386 9616
rect 2686 3476 2688 3496
rect 2688 3476 2740 3496
rect 2740 3476 2742 3496
rect 2686 3440 2742 3476
rect 3330 7928 3386 7984
rect 3882 12144 3938 12200
rect 4250 12280 4306 12336
rect 4158 12008 4214 12064
rect 3923 11450 3979 11452
rect 4003 11450 4059 11452
rect 4083 11450 4139 11452
rect 4163 11450 4219 11452
rect 3923 11398 3969 11450
rect 3969 11398 3979 11450
rect 4003 11398 4033 11450
rect 4033 11398 4045 11450
rect 4045 11398 4059 11450
rect 4083 11398 4097 11450
rect 4097 11398 4109 11450
rect 4109 11398 4139 11450
rect 4163 11398 4173 11450
rect 4173 11398 4219 11450
rect 3923 11396 3979 11398
rect 4003 11396 4059 11398
rect 4083 11396 4139 11398
rect 4163 11396 4219 11398
rect 4802 13368 4858 13424
rect 3974 10648 4030 10704
rect 4066 10548 4068 10568
rect 4068 10548 4120 10568
rect 4120 10548 4122 10568
rect 4066 10512 4122 10548
rect 3923 10362 3979 10364
rect 4003 10362 4059 10364
rect 4083 10362 4139 10364
rect 4163 10362 4219 10364
rect 3923 10310 3969 10362
rect 3969 10310 3979 10362
rect 4003 10310 4033 10362
rect 4033 10310 4045 10362
rect 4045 10310 4059 10362
rect 4083 10310 4097 10362
rect 4097 10310 4109 10362
rect 4109 10310 4139 10362
rect 4163 10310 4173 10362
rect 4173 10310 4219 10362
rect 3923 10308 3979 10310
rect 4003 10308 4059 10310
rect 4083 10308 4139 10310
rect 4163 10308 4219 10310
rect 3974 10104 4030 10160
rect 3974 10004 3976 10024
rect 3976 10004 4028 10024
rect 4028 10004 4030 10024
rect 3974 9968 4030 10004
rect 3923 9274 3979 9276
rect 4003 9274 4059 9276
rect 4083 9274 4139 9276
rect 4163 9274 4219 9276
rect 3923 9222 3969 9274
rect 3969 9222 3979 9274
rect 4003 9222 4033 9274
rect 4033 9222 4045 9274
rect 4045 9222 4059 9274
rect 4083 9222 4097 9274
rect 4097 9222 4109 9274
rect 4109 9222 4139 9274
rect 4163 9222 4173 9274
rect 4173 9222 4219 9274
rect 3923 9220 3979 9222
rect 4003 9220 4059 9222
rect 4083 9220 4139 9222
rect 4163 9220 4219 9222
rect 3238 6332 3240 6352
rect 3240 6332 3292 6352
rect 3292 6332 3294 6352
rect 3238 6296 3294 6332
rect 3514 7112 3570 7168
rect 3330 3984 3386 4040
rect 3923 8186 3979 8188
rect 4003 8186 4059 8188
rect 4083 8186 4139 8188
rect 4163 8186 4219 8188
rect 3923 8134 3969 8186
rect 3969 8134 3979 8186
rect 4003 8134 4033 8186
rect 4033 8134 4045 8186
rect 4045 8134 4059 8186
rect 4083 8134 4097 8186
rect 4097 8134 4109 8186
rect 4109 8134 4139 8186
rect 4163 8134 4173 8186
rect 4173 8134 4219 8186
rect 3923 8132 3979 8134
rect 4003 8132 4059 8134
rect 4083 8132 4139 8134
rect 4163 8132 4219 8134
rect 3923 7098 3979 7100
rect 4003 7098 4059 7100
rect 4083 7098 4139 7100
rect 4163 7098 4219 7100
rect 3923 7046 3969 7098
rect 3969 7046 3979 7098
rect 4003 7046 4033 7098
rect 4033 7046 4045 7098
rect 4045 7046 4059 7098
rect 4083 7046 4097 7098
rect 4097 7046 4109 7098
rect 4109 7046 4139 7098
rect 4163 7046 4173 7098
rect 4173 7046 4219 7098
rect 3923 7044 3979 7046
rect 4003 7044 4059 7046
rect 4083 7044 4139 7046
rect 4163 7044 4219 7046
rect 4250 6840 4306 6896
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 4066 5752 4122 5808
rect 4802 12416 4858 12472
rect 4710 11736 4766 11792
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 3974 4564 3976 4584
rect 3976 4564 4028 4584
rect 4028 4564 4030 4584
rect 3974 4528 4030 4564
rect 4526 4936 4582 4992
rect 5078 12552 5134 12608
rect 4894 8336 4950 8392
rect 4894 5208 4950 5264
rect 4434 4256 4490 4312
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 4066 2932 4068 2952
rect 4068 2932 4120 2952
rect 4120 2932 4122 2952
rect 4066 2896 4122 2932
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 3974 1264 4030 1320
rect 4066 1128 4122 1184
rect 5078 3712 5134 3768
rect 4894 3340 4896 3360
rect 4896 3340 4948 3360
rect 4948 3340 4950 3360
rect 4894 3304 4950 3340
rect 5354 18400 5410 18456
rect 6182 21800 6238 21856
rect 6090 21392 6146 21448
rect 5630 14592 5686 14648
rect 5998 19216 6054 19272
rect 5998 17756 6000 17776
rect 6000 17756 6052 17776
rect 6052 17756 6054 17776
rect 5998 17720 6054 17756
rect 5814 14728 5870 14784
rect 5354 14320 5410 14376
rect 5262 11756 5318 11792
rect 5262 11736 5264 11756
rect 5264 11736 5316 11756
rect 5316 11736 5318 11756
rect 5446 14048 5502 14104
rect 5906 14048 5962 14104
rect 5630 13912 5686 13968
rect 5446 11192 5502 11248
rect 5906 13504 5962 13560
rect 6458 23024 6514 23080
rect 6366 18264 6422 18320
rect 7102 31864 7158 31920
rect 7930 41656 7986 41712
rect 8390 42744 8446 42800
rect 7470 40180 7526 40216
rect 7470 40160 7472 40180
rect 7472 40160 7524 40180
rect 7524 40160 7526 40180
rect 7378 36116 7380 36136
rect 7380 36116 7432 36136
rect 7432 36116 7434 36136
rect 7378 36080 7434 36116
rect 7746 36780 7802 36816
rect 7746 36760 7748 36780
rect 7748 36760 7800 36780
rect 7800 36760 7802 36780
rect 7838 34856 7894 34912
rect 7838 33632 7894 33688
rect 6890 31578 6946 31580
rect 6970 31578 7026 31580
rect 7050 31578 7106 31580
rect 7130 31578 7186 31580
rect 6890 31526 6936 31578
rect 6936 31526 6946 31578
rect 6970 31526 7000 31578
rect 7000 31526 7012 31578
rect 7012 31526 7026 31578
rect 7050 31526 7064 31578
rect 7064 31526 7076 31578
rect 7076 31526 7106 31578
rect 7130 31526 7140 31578
rect 7140 31526 7186 31578
rect 6890 31524 6946 31526
rect 6970 31524 7026 31526
rect 7050 31524 7106 31526
rect 7130 31524 7186 31526
rect 6890 30490 6946 30492
rect 6970 30490 7026 30492
rect 7050 30490 7106 30492
rect 7130 30490 7186 30492
rect 6890 30438 6936 30490
rect 6936 30438 6946 30490
rect 6970 30438 7000 30490
rect 7000 30438 7012 30490
rect 7012 30438 7026 30490
rect 7050 30438 7064 30490
rect 7064 30438 7076 30490
rect 7076 30438 7106 30490
rect 7130 30438 7140 30490
rect 7140 30438 7186 30490
rect 6890 30436 6946 30438
rect 6970 30436 7026 30438
rect 7050 30436 7106 30438
rect 7130 30436 7186 30438
rect 7102 29588 7104 29608
rect 7104 29588 7156 29608
rect 7156 29588 7158 29608
rect 7102 29552 7158 29588
rect 6890 29402 6946 29404
rect 6970 29402 7026 29404
rect 7050 29402 7106 29404
rect 7130 29402 7186 29404
rect 6890 29350 6936 29402
rect 6936 29350 6946 29402
rect 6970 29350 7000 29402
rect 7000 29350 7012 29402
rect 7012 29350 7026 29402
rect 7050 29350 7064 29402
rect 7064 29350 7076 29402
rect 7076 29350 7106 29402
rect 7130 29350 7140 29402
rect 7140 29350 7186 29402
rect 6890 29348 6946 29350
rect 6970 29348 7026 29350
rect 7050 29348 7106 29350
rect 7130 29348 7186 29350
rect 6734 29280 6790 29336
rect 7102 29028 7158 29064
rect 7102 29008 7104 29028
rect 7104 29008 7156 29028
rect 7156 29008 7158 29028
rect 6890 28314 6946 28316
rect 6970 28314 7026 28316
rect 7050 28314 7106 28316
rect 7130 28314 7186 28316
rect 6890 28262 6936 28314
rect 6936 28262 6946 28314
rect 6970 28262 7000 28314
rect 7000 28262 7012 28314
rect 7012 28262 7026 28314
rect 7050 28262 7064 28314
rect 7064 28262 7076 28314
rect 7076 28262 7106 28314
rect 7130 28262 7140 28314
rect 7140 28262 7186 28314
rect 6890 28260 6946 28262
rect 6970 28260 7026 28262
rect 7050 28260 7106 28262
rect 7130 28260 7186 28262
rect 6826 28056 6882 28112
rect 7194 27784 7250 27840
rect 7102 27512 7158 27568
rect 6734 27240 6790 27296
rect 6890 27226 6946 27228
rect 6970 27226 7026 27228
rect 7050 27226 7106 27228
rect 7130 27226 7186 27228
rect 6890 27174 6936 27226
rect 6936 27174 6946 27226
rect 6970 27174 7000 27226
rect 7000 27174 7012 27226
rect 7012 27174 7026 27226
rect 7050 27174 7064 27226
rect 7064 27174 7076 27226
rect 7076 27174 7106 27226
rect 7130 27174 7140 27226
rect 7140 27174 7186 27226
rect 6890 27172 6946 27174
rect 6970 27172 7026 27174
rect 7050 27172 7106 27174
rect 7130 27172 7186 27174
rect 7286 26832 7342 26888
rect 6734 26424 6790 26480
rect 6890 26138 6946 26140
rect 6970 26138 7026 26140
rect 7050 26138 7106 26140
rect 7130 26138 7186 26140
rect 6890 26086 6936 26138
rect 6936 26086 6946 26138
rect 6970 26086 7000 26138
rect 7000 26086 7012 26138
rect 7012 26086 7026 26138
rect 7050 26086 7064 26138
rect 7064 26086 7076 26138
rect 7076 26086 7106 26138
rect 7130 26086 7140 26138
rect 7140 26086 7186 26138
rect 6890 26084 6946 26086
rect 6970 26084 7026 26086
rect 7050 26084 7106 26086
rect 7130 26084 7186 26086
rect 6826 25472 6882 25528
rect 6826 25200 6882 25256
rect 7010 25236 7012 25256
rect 7012 25236 7064 25256
rect 7064 25236 7066 25256
rect 7010 25200 7066 25236
rect 6890 25050 6946 25052
rect 6970 25050 7026 25052
rect 7050 25050 7106 25052
rect 7130 25050 7186 25052
rect 6890 24998 6936 25050
rect 6936 24998 6946 25050
rect 6970 24998 7000 25050
rect 7000 24998 7012 25050
rect 7012 24998 7026 25050
rect 7050 24998 7064 25050
rect 7064 24998 7076 25050
rect 7076 24998 7106 25050
rect 7130 24998 7140 25050
rect 7140 24998 7186 25050
rect 6890 24996 6946 24998
rect 6970 24996 7026 24998
rect 7050 24996 7106 24998
rect 7130 24996 7186 24998
rect 6890 23962 6946 23964
rect 6970 23962 7026 23964
rect 7050 23962 7106 23964
rect 7130 23962 7186 23964
rect 6890 23910 6936 23962
rect 6936 23910 6946 23962
rect 6970 23910 7000 23962
rect 7000 23910 7012 23962
rect 7012 23910 7026 23962
rect 7050 23910 7064 23962
rect 7064 23910 7076 23962
rect 7076 23910 7106 23962
rect 7130 23910 7140 23962
rect 7140 23910 7186 23962
rect 6890 23908 6946 23910
rect 6970 23908 7026 23910
rect 7050 23908 7106 23910
rect 7130 23908 7186 23910
rect 6890 22874 6946 22876
rect 6970 22874 7026 22876
rect 7050 22874 7106 22876
rect 7130 22874 7186 22876
rect 6890 22822 6936 22874
rect 6936 22822 6946 22874
rect 6970 22822 7000 22874
rect 7000 22822 7012 22874
rect 7012 22822 7026 22874
rect 7050 22822 7064 22874
rect 7064 22822 7076 22874
rect 7076 22822 7106 22874
rect 7130 22822 7140 22874
rect 7140 22822 7186 22874
rect 6890 22820 6946 22822
rect 6970 22820 7026 22822
rect 7050 22820 7106 22822
rect 7130 22820 7186 22822
rect 6826 22072 6882 22128
rect 7562 29416 7618 29472
rect 7470 28464 7526 28520
rect 7470 28192 7526 28248
rect 7470 27376 7526 27432
rect 7470 26968 7526 27024
rect 7654 29164 7710 29200
rect 7654 29144 7656 29164
rect 7656 29144 7708 29164
rect 7708 29144 7710 29164
rect 7838 31204 7894 31240
rect 7838 31184 7840 31204
rect 7840 31184 7892 31204
rect 7892 31184 7894 31204
rect 8298 41928 8354 41984
rect 8206 37304 8262 37360
rect 8666 39344 8722 39400
rect 8298 34584 8354 34640
rect 8114 33632 8170 33688
rect 8206 32408 8262 32464
rect 8022 31320 8078 31376
rect 8022 30912 8078 30968
rect 7654 26288 7710 26344
rect 7654 25916 7656 25936
rect 7656 25916 7708 25936
rect 7708 25916 7710 25936
rect 7654 25880 7710 25916
rect 6890 21786 6946 21788
rect 6970 21786 7026 21788
rect 7050 21786 7106 21788
rect 7130 21786 7186 21788
rect 6890 21734 6936 21786
rect 6936 21734 6946 21786
rect 6970 21734 7000 21786
rect 7000 21734 7012 21786
rect 7012 21734 7026 21786
rect 7050 21734 7064 21786
rect 7064 21734 7076 21786
rect 7076 21734 7106 21786
rect 7130 21734 7140 21786
rect 7140 21734 7186 21786
rect 6890 21732 6946 21734
rect 6970 21732 7026 21734
rect 7050 21732 7106 21734
rect 7130 21732 7186 21734
rect 7194 20848 7250 20904
rect 6890 20698 6946 20700
rect 6970 20698 7026 20700
rect 7050 20698 7106 20700
rect 7130 20698 7186 20700
rect 6890 20646 6936 20698
rect 6936 20646 6946 20698
rect 6970 20646 7000 20698
rect 7000 20646 7012 20698
rect 7012 20646 7026 20698
rect 7050 20646 7064 20698
rect 7064 20646 7076 20698
rect 7076 20646 7106 20698
rect 7130 20646 7140 20698
rect 7140 20646 7186 20698
rect 6890 20644 6946 20646
rect 6970 20644 7026 20646
rect 7050 20644 7106 20646
rect 7130 20644 7186 20646
rect 6826 19760 6882 19816
rect 6890 19610 6946 19612
rect 6970 19610 7026 19612
rect 7050 19610 7106 19612
rect 7130 19610 7186 19612
rect 6890 19558 6936 19610
rect 6936 19558 6946 19610
rect 6970 19558 7000 19610
rect 7000 19558 7012 19610
rect 7012 19558 7026 19610
rect 7050 19558 7064 19610
rect 7064 19558 7076 19610
rect 7076 19558 7106 19610
rect 7130 19558 7140 19610
rect 7140 19558 7186 19610
rect 6890 19556 6946 19558
rect 6970 19556 7026 19558
rect 7050 19556 7106 19558
rect 7130 19556 7186 19558
rect 8298 29008 8354 29064
rect 8758 35400 8814 35456
rect 8758 34060 8814 34096
rect 8758 34040 8760 34060
rect 8760 34040 8812 34060
rect 8812 34040 8814 34060
rect 8574 31456 8630 31512
rect 8114 25200 8170 25256
rect 8206 24928 8262 24984
rect 8114 23044 8170 23080
rect 8114 23024 8116 23044
rect 8116 23024 8168 23044
rect 8168 23024 8170 23044
rect 7654 21800 7710 21856
rect 6890 18522 6946 18524
rect 6970 18522 7026 18524
rect 7050 18522 7106 18524
rect 7130 18522 7186 18524
rect 6890 18470 6936 18522
rect 6936 18470 6946 18522
rect 6970 18470 7000 18522
rect 7000 18470 7012 18522
rect 7012 18470 7026 18522
rect 7050 18470 7064 18522
rect 7064 18470 7076 18522
rect 7076 18470 7106 18522
rect 7130 18470 7140 18522
rect 7140 18470 7186 18522
rect 6890 18468 6946 18470
rect 6970 18468 7026 18470
rect 7050 18468 7106 18470
rect 7130 18468 7186 18470
rect 6734 18264 6790 18320
rect 6550 17212 6552 17232
rect 6552 17212 6604 17232
rect 6604 17212 6606 17232
rect 6550 17176 6606 17212
rect 6182 16088 6238 16144
rect 6090 13368 6146 13424
rect 5906 12300 5962 12336
rect 5906 12280 5908 12300
rect 5908 12280 5960 12300
rect 5960 12280 5962 12300
rect 5998 10648 6054 10704
rect 5998 9424 6054 9480
rect 6274 12844 6330 12880
rect 6274 12824 6276 12844
rect 6276 12824 6328 12844
rect 6328 12824 6330 12844
rect 5906 5072 5962 5128
rect 5998 4972 6000 4992
rect 6000 4972 6052 4992
rect 6052 4972 6054 4992
rect 5998 4936 6054 4972
rect 5538 1808 5594 1864
rect 6182 2352 6238 2408
rect 5538 1300 5540 1320
rect 5540 1300 5592 1320
rect 5592 1300 5594 1320
rect 5538 1264 5594 1300
rect 6550 15000 6606 15056
rect 6890 17434 6946 17436
rect 6970 17434 7026 17436
rect 7050 17434 7106 17436
rect 7130 17434 7186 17436
rect 6890 17382 6936 17434
rect 6936 17382 6946 17434
rect 6970 17382 7000 17434
rect 7000 17382 7012 17434
rect 7012 17382 7026 17434
rect 7050 17382 7064 17434
rect 7064 17382 7076 17434
rect 7076 17382 7106 17434
rect 7130 17382 7140 17434
rect 7140 17382 7186 17434
rect 6890 17380 6946 17382
rect 6970 17380 7026 17382
rect 7050 17380 7106 17382
rect 7130 17380 7186 17382
rect 6918 17040 6974 17096
rect 7838 21412 7894 21448
rect 7838 21392 7840 21412
rect 7840 21392 7892 21412
rect 7892 21392 7894 21412
rect 7838 21256 7894 21312
rect 7838 20884 7840 20904
rect 7840 20884 7892 20904
rect 7892 20884 7894 20904
rect 7838 20848 7894 20884
rect 7746 19760 7802 19816
rect 7562 18808 7618 18864
rect 7470 16904 7526 16960
rect 6890 16346 6946 16348
rect 6970 16346 7026 16348
rect 7050 16346 7106 16348
rect 7130 16346 7186 16348
rect 6890 16294 6936 16346
rect 6936 16294 6946 16346
rect 6970 16294 7000 16346
rect 7000 16294 7012 16346
rect 7012 16294 7026 16346
rect 7050 16294 7064 16346
rect 7064 16294 7076 16346
rect 7076 16294 7106 16346
rect 7130 16294 7140 16346
rect 7140 16294 7186 16346
rect 6890 16292 6946 16294
rect 6970 16292 7026 16294
rect 7050 16292 7106 16294
rect 7130 16292 7186 16294
rect 6890 15258 6946 15260
rect 6970 15258 7026 15260
rect 7050 15258 7106 15260
rect 7130 15258 7186 15260
rect 6890 15206 6936 15258
rect 6936 15206 6946 15258
rect 6970 15206 7000 15258
rect 7000 15206 7012 15258
rect 7012 15206 7026 15258
rect 7050 15206 7064 15258
rect 7064 15206 7076 15258
rect 7076 15206 7106 15258
rect 7130 15206 7140 15258
rect 7140 15206 7186 15258
rect 6890 15204 6946 15206
rect 6970 15204 7026 15206
rect 7050 15204 7106 15206
rect 7130 15204 7186 15206
rect 7378 16496 7434 16552
rect 6826 15000 6882 15056
rect 6826 14320 6882 14376
rect 6890 14170 6946 14172
rect 6970 14170 7026 14172
rect 7050 14170 7106 14172
rect 7130 14170 7186 14172
rect 6890 14118 6936 14170
rect 6936 14118 6946 14170
rect 6970 14118 7000 14170
rect 7000 14118 7012 14170
rect 7012 14118 7026 14170
rect 7050 14118 7064 14170
rect 7064 14118 7076 14170
rect 7076 14118 7106 14170
rect 7130 14118 7140 14170
rect 7140 14118 7186 14170
rect 6890 14116 6946 14118
rect 6970 14116 7026 14118
rect 7050 14116 7106 14118
rect 7130 14116 7186 14118
rect 6642 13368 6698 13424
rect 6890 13082 6946 13084
rect 6970 13082 7026 13084
rect 7050 13082 7106 13084
rect 7130 13082 7186 13084
rect 6890 13030 6936 13082
rect 6936 13030 6946 13082
rect 6970 13030 7000 13082
rect 7000 13030 7012 13082
rect 7012 13030 7026 13082
rect 7050 13030 7064 13082
rect 7064 13030 7076 13082
rect 7076 13030 7106 13082
rect 7130 13030 7140 13082
rect 7140 13030 7186 13082
rect 6890 13028 6946 13030
rect 6970 13028 7026 13030
rect 7050 13028 7106 13030
rect 7130 13028 7186 13030
rect 6890 11994 6946 11996
rect 6970 11994 7026 11996
rect 7050 11994 7106 11996
rect 7130 11994 7186 11996
rect 6890 11942 6936 11994
rect 6936 11942 6946 11994
rect 6970 11942 7000 11994
rect 7000 11942 7012 11994
rect 7012 11942 7026 11994
rect 7050 11942 7064 11994
rect 7064 11942 7076 11994
rect 7076 11942 7106 11994
rect 7130 11942 7140 11994
rect 7140 11942 7186 11994
rect 6890 11940 6946 11942
rect 6970 11940 7026 11942
rect 7050 11940 7106 11942
rect 7130 11940 7186 11942
rect 7010 11192 7066 11248
rect 6890 10906 6946 10908
rect 6970 10906 7026 10908
rect 7050 10906 7106 10908
rect 7130 10906 7186 10908
rect 6890 10854 6936 10906
rect 6936 10854 6946 10906
rect 6970 10854 7000 10906
rect 7000 10854 7012 10906
rect 7012 10854 7026 10906
rect 7050 10854 7064 10906
rect 7064 10854 7076 10906
rect 7076 10854 7106 10906
rect 7130 10854 7140 10906
rect 7140 10854 7186 10906
rect 6890 10852 6946 10854
rect 6970 10852 7026 10854
rect 7050 10852 7106 10854
rect 7130 10852 7186 10854
rect 6826 10512 6882 10568
rect 6550 3576 6606 3632
rect 6890 9818 6946 9820
rect 6970 9818 7026 9820
rect 7050 9818 7106 9820
rect 7130 9818 7186 9820
rect 6890 9766 6936 9818
rect 6936 9766 6946 9818
rect 6970 9766 7000 9818
rect 7000 9766 7012 9818
rect 7012 9766 7026 9818
rect 7050 9766 7064 9818
rect 7064 9766 7076 9818
rect 7076 9766 7106 9818
rect 7130 9766 7140 9818
rect 7140 9766 7186 9818
rect 6890 9764 6946 9766
rect 6970 9764 7026 9766
rect 7050 9764 7106 9766
rect 7130 9764 7186 9766
rect 7838 16108 7894 16144
rect 7838 16088 7840 16108
rect 7840 16088 7892 16108
rect 7892 16088 7894 16108
rect 8482 22208 8538 22264
rect 8298 21120 8354 21176
rect 8114 20748 8116 20768
rect 8116 20748 8168 20768
rect 8168 20748 8170 20768
rect 8114 20712 8170 20748
rect 8022 19080 8078 19136
rect 8206 19388 8208 19408
rect 8208 19388 8260 19408
rect 8260 19388 8262 19408
rect 8206 19352 8262 19388
rect 8758 30232 8814 30288
rect 8942 40160 8998 40216
rect 9126 42608 9182 42664
rect 9126 40160 9182 40216
rect 9857 43002 9913 43004
rect 9937 43002 9993 43004
rect 10017 43002 10073 43004
rect 10097 43002 10153 43004
rect 9857 42950 9903 43002
rect 9903 42950 9913 43002
rect 9937 42950 9967 43002
rect 9967 42950 9979 43002
rect 9979 42950 9993 43002
rect 10017 42950 10031 43002
rect 10031 42950 10043 43002
rect 10043 42950 10073 43002
rect 10097 42950 10107 43002
rect 10107 42950 10153 43002
rect 9857 42948 9913 42950
rect 9937 42948 9993 42950
rect 10017 42948 10073 42950
rect 10097 42948 10153 42950
rect 9402 42744 9458 42800
rect 9402 41792 9458 41848
rect 9862 42064 9918 42120
rect 9857 41914 9913 41916
rect 9937 41914 9993 41916
rect 10017 41914 10073 41916
rect 10097 41914 10153 41916
rect 9857 41862 9903 41914
rect 9903 41862 9913 41914
rect 9937 41862 9967 41914
rect 9967 41862 9979 41914
rect 9979 41862 9993 41914
rect 10017 41862 10031 41914
rect 10031 41862 10043 41914
rect 10043 41862 10073 41914
rect 10097 41862 10107 41914
rect 10107 41862 10153 41914
rect 9857 41860 9913 41862
rect 9937 41860 9993 41862
rect 10017 41860 10073 41862
rect 10097 41860 10153 41862
rect 8942 36080 8998 36136
rect 9034 34584 9090 34640
rect 9857 40826 9913 40828
rect 9937 40826 9993 40828
rect 10017 40826 10073 40828
rect 10097 40826 10153 40828
rect 9857 40774 9903 40826
rect 9903 40774 9913 40826
rect 9937 40774 9967 40826
rect 9967 40774 9979 40826
rect 9979 40774 9993 40826
rect 10017 40774 10031 40826
rect 10031 40774 10043 40826
rect 10043 40774 10073 40826
rect 10097 40774 10107 40826
rect 10107 40774 10153 40826
rect 9857 40772 9913 40774
rect 9937 40772 9993 40774
rect 10017 40772 10073 40774
rect 10097 40772 10153 40774
rect 9857 39738 9913 39740
rect 9937 39738 9993 39740
rect 10017 39738 10073 39740
rect 10097 39738 10153 39740
rect 9857 39686 9903 39738
rect 9903 39686 9913 39738
rect 9937 39686 9967 39738
rect 9967 39686 9979 39738
rect 9979 39686 9993 39738
rect 10017 39686 10031 39738
rect 10031 39686 10043 39738
rect 10043 39686 10073 39738
rect 10097 39686 10107 39738
rect 10107 39686 10153 39738
rect 9857 39684 9913 39686
rect 9937 39684 9993 39686
rect 10017 39684 10073 39686
rect 10097 39684 10153 39686
rect 9857 38650 9913 38652
rect 9937 38650 9993 38652
rect 10017 38650 10073 38652
rect 10097 38650 10153 38652
rect 9857 38598 9903 38650
rect 9903 38598 9913 38650
rect 9937 38598 9967 38650
rect 9967 38598 9979 38650
rect 9979 38598 9993 38650
rect 10017 38598 10031 38650
rect 10031 38598 10043 38650
rect 10043 38598 10073 38650
rect 10097 38598 10107 38650
rect 10107 38598 10153 38650
rect 9857 38596 9913 38598
rect 9937 38596 9993 38598
rect 10017 38596 10073 38598
rect 10097 38596 10153 38598
rect 9857 37562 9913 37564
rect 9937 37562 9993 37564
rect 10017 37562 10073 37564
rect 10097 37562 10153 37564
rect 9857 37510 9903 37562
rect 9903 37510 9913 37562
rect 9937 37510 9967 37562
rect 9967 37510 9979 37562
rect 9979 37510 9993 37562
rect 10017 37510 10031 37562
rect 10031 37510 10043 37562
rect 10043 37510 10073 37562
rect 10097 37510 10107 37562
rect 10107 37510 10153 37562
rect 9857 37508 9913 37510
rect 9937 37508 9993 37510
rect 10017 37508 10073 37510
rect 10097 37508 10153 37510
rect 9402 36080 9458 36136
rect 9857 36474 9913 36476
rect 9937 36474 9993 36476
rect 10017 36474 10073 36476
rect 10097 36474 10153 36476
rect 9857 36422 9903 36474
rect 9903 36422 9913 36474
rect 9937 36422 9967 36474
rect 9967 36422 9979 36474
rect 9979 36422 9993 36474
rect 10017 36422 10031 36474
rect 10031 36422 10043 36474
rect 10043 36422 10073 36474
rect 10097 36422 10107 36474
rect 10107 36422 10153 36474
rect 9857 36420 9913 36422
rect 9937 36420 9993 36422
rect 10017 36420 10073 36422
rect 10097 36420 10153 36422
rect 9218 34856 9274 34912
rect 9586 34856 9642 34912
rect 9126 34312 9182 34368
rect 8942 33940 8944 33960
rect 8944 33940 8996 33960
rect 8996 33940 8998 33960
rect 8942 33904 8998 33940
rect 9494 34348 9496 34368
rect 9496 34348 9548 34368
rect 9548 34348 9550 34368
rect 9494 34312 9550 34348
rect 9857 35386 9913 35388
rect 9937 35386 9993 35388
rect 10017 35386 10073 35388
rect 10097 35386 10153 35388
rect 9857 35334 9903 35386
rect 9903 35334 9913 35386
rect 9937 35334 9967 35386
rect 9967 35334 9979 35386
rect 9979 35334 9993 35386
rect 10017 35334 10031 35386
rect 10031 35334 10043 35386
rect 10043 35334 10073 35386
rect 10097 35334 10107 35386
rect 10107 35334 10153 35386
rect 9857 35332 9913 35334
rect 9937 35332 9993 35334
rect 10017 35332 10073 35334
rect 10097 35332 10153 35334
rect 10046 35128 10102 35184
rect 10414 35808 10470 35864
rect 10414 35264 10470 35320
rect 9857 34298 9913 34300
rect 9937 34298 9993 34300
rect 10017 34298 10073 34300
rect 10097 34298 10153 34300
rect 9857 34246 9903 34298
rect 9903 34246 9913 34298
rect 9937 34246 9967 34298
rect 9967 34246 9979 34298
rect 9979 34246 9993 34298
rect 10017 34246 10031 34298
rect 10031 34246 10043 34298
rect 10043 34246 10073 34298
rect 10097 34246 10107 34298
rect 10107 34246 10153 34298
rect 9857 34244 9913 34246
rect 9937 34244 9993 34246
rect 10017 34244 10073 34246
rect 10097 34244 10153 34246
rect 9402 33224 9458 33280
rect 8666 26152 8722 26208
rect 8758 25780 8760 25800
rect 8760 25780 8812 25800
rect 8812 25780 8814 25800
rect 8758 25744 8814 25780
rect 8758 25472 8814 25528
rect 8942 29008 8998 29064
rect 8942 25880 8998 25936
rect 9862 33360 9918 33416
rect 9857 33210 9913 33212
rect 9937 33210 9993 33212
rect 10017 33210 10073 33212
rect 10097 33210 10153 33212
rect 9857 33158 9903 33210
rect 9903 33158 9913 33210
rect 9937 33158 9967 33210
rect 9967 33158 9979 33210
rect 9979 33158 9993 33210
rect 10017 33158 10031 33210
rect 10031 33158 10043 33210
rect 10043 33158 10073 33210
rect 10097 33158 10107 33210
rect 10107 33158 10153 33210
rect 9857 33156 9913 33158
rect 9937 33156 9993 33158
rect 10017 33156 10073 33158
rect 10097 33156 10153 33158
rect 10138 32272 10194 32328
rect 9857 32122 9913 32124
rect 9937 32122 9993 32124
rect 10017 32122 10073 32124
rect 10097 32122 10153 32124
rect 9857 32070 9903 32122
rect 9903 32070 9913 32122
rect 9937 32070 9967 32122
rect 9967 32070 9979 32122
rect 9979 32070 9993 32122
rect 10017 32070 10031 32122
rect 10031 32070 10043 32122
rect 10043 32070 10073 32122
rect 10097 32070 10107 32122
rect 10107 32070 10153 32122
rect 9857 32068 9913 32070
rect 9937 32068 9993 32070
rect 10017 32068 10073 32070
rect 10097 32068 10153 32070
rect 9678 31048 9734 31104
rect 9857 31034 9913 31036
rect 9937 31034 9993 31036
rect 10017 31034 10073 31036
rect 10097 31034 10153 31036
rect 9857 30982 9903 31034
rect 9903 30982 9913 31034
rect 9937 30982 9967 31034
rect 9967 30982 9979 31034
rect 9979 30982 9993 31034
rect 10017 30982 10031 31034
rect 10031 30982 10043 31034
rect 10043 30982 10073 31034
rect 10097 30982 10107 31034
rect 10107 30982 10153 31034
rect 9857 30980 9913 30982
rect 9937 30980 9993 30982
rect 10017 30980 10073 30982
rect 10097 30980 10153 30982
rect 10138 30640 10194 30696
rect 11702 42880 11758 42936
rect 12824 43546 12880 43548
rect 12904 43546 12960 43548
rect 12984 43546 13040 43548
rect 13064 43546 13120 43548
rect 12824 43494 12870 43546
rect 12870 43494 12880 43546
rect 12904 43494 12934 43546
rect 12934 43494 12946 43546
rect 12946 43494 12960 43546
rect 12984 43494 12998 43546
rect 12998 43494 13010 43546
rect 13010 43494 13040 43546
rect 13064 43494 13074 43546
rect 13074 43494 13120 43546
rect 12824 43492 12880 43494
rect 12904 43492 12960 43494
rect 12984 43492 13040 43494
rect 13064 43492 13120 43494
rect 12254 42880 12310 42936
rect 12530 42880 12586 42936
rect 11794 42200 11850 42256
rect 10690 34620 10692 34640
rect 10692 34620 10744 34640
rect 10744 34620 10746 34640
rect 10690 34584 10746 34620
rect 11242 33904 11298 33960
rect 10874 31864 10930 31920
rect 9857 29946 9913 29948
rect 9937 29946 9993 29948
rect 10017 29946 10073 29948
rect 10097 29946 10153 29948
rect 9857 29894 9903 29946
rect 9903 29894 9913 29946
rect 9937 29894 9967 29946
rect 9967 29894 9979 29946
rect 9979 29894 9993 29946
rect 10017 29894 10031 29946
rect 10031 29894 10043 29946
rect 10043 29894 10073 29946
rect 10097 29894 10107 29946
rect 10107 29894 10153 29946
rect 9857 29892 9913 29894
rect 9937 29892 9993 29894
rect 10017 29892 10073 29894
rect 10097 29892 10153 29894
rect 9402 28736 9458 28792
rect 9402 28464 9458 28520
rect 8298 17992 8354 18048
rect 7838 12300 7894 12336
rect 7838 12280 7840 12300
rect 7840 12280 7892 12300
rect 7892 12280 7894 12300
rect 7562 11736 7618 11792
rect 7562 10920 7618 10976
rect 6890 8730 6946 8732
rect 6970 8730 7026 8732
rect 7050 8730 7106 8732
rect 7130 8730 7186 8732
rect 6890 8678 6936 8730
rect 6936 8678 6946 8730
rect 6970 8678 7000 8730
rect 7000 8678 7012 8730
rect 7012 8678 7026 8730
rect 7050 8678 7064 8730
rect 7064 8678 7076 8730
rect 7076 8678 7106 8730
rect 7130 8678 7140 8730
rect 7140 8678 7186 8730
rect 6890 8676 6946 8678
rect 6970 8676 7026 8678
rect 7050 8676 7106 8678
rect 7130 8676 7186 8678
rect 7194 8084 7250 8120
rect 7194 8064 7196 8084
rect 7196 8064 7248 8084
rect 7248 8064 7250 8084
rect 6890 7642 6946 7644
rect 6970 7642 7026 7644
rect 7050 7642 7106 7644
rect 7130 7642 7186 7644
rect 6890 7590 6936 7642
rect 6936 7590 6946 7642
rect 6970 7590 7000 7642
rect 7000 7590 7012 7642
rect 7012 7590 7026 7642
rect 7050 7590 7064 7642
rect 7064 7590 7076 7642
rect 7076 7590 7106 7642
rect 7130 7590 7140 7642
rect 7140 7590 7186 7642
rect 6890 7588 6946 7590
rect 6970 7588 7026 7590
rect 7050 7588 7106 7590
rect 7130 7588 7186 7590
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 6918 5616 6974 5672
rect 7470 5752 7526 5808
rect 7286 5616 7342 5672
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 6826 4548 6882 4584
rect 6826 4528 6828 4548
rect 6828 4528 6880 4548
rect 6880 4528 6882 4548
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 7930 9968 7986 10024
rect 7838 6840 7894 6896
rect 6550 2488 6606 2544
rect 7194 2352 7250 2408
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 8666 18572 8668 18592
rect 8668 18572 8720 18592
rect 8720 18572 8722 18592
rect 8666 18536 8722 18572
rect 8850 20168 8906 20224
rect 8298 8064 8354 8120
rect 8298 7792 8354 7848
rect 9126 20032 9182 20088
rect 8206 6160 8262 6216
rect 9586 28328 9642 28384
rect 9857 28858 9913 28860
rect 9937 28858 9993 28860
rect 10017 28858 10073 28860
rect 10097 28858 10153 28860
rect 9857 28806 9903 28858
rect 9903 28806 9913 28858
rect 9937 28806 9967 28858
rect 9967 28806 9979 28858
rect 9979 28806 9993 28858
rect 10017 28806 10031 28858
rect 10031 28806 10043 28858
rect 10043 28806 10073 28858
rect 10097 28806 10107 28858
rect 10107 28806 10153 28858
rect 9857 28804 9913 28806
rect 9937 28804 9993 28806
rect 10017 28804 10073 28806
rect 10097 28804 10153 28806
rect 9857 27770 9913 27772
rect 9937 27770 9993 27772
rect 10017 27770 10073 27772
rect 10097 27770 10153 27772
rect 9857 27718 9903 27770
rect 9903 27718 9913 27770
rect 9937 27718 9967 27770
rect 9967 27718 9979 27770
rect 9979 27718 9993 27770
rect 10017 27718 10031 27770
rect 10031 27718 10043 27770
rect 10043 27718 10073 27770
rect 10097 27718 10107 27770
rect 10107 27718 10153 27770
rect 9857 27716 9913 27718
rect 9937 27716 9993 27718
rect 10017 27716 10073 27718
rect 10097 27716 10153 27718
rect 10506 27920 10562 27976
rect 10414 27548 10416 27568
rect 10416 27548 10468 27568
rect 10468 27548 10470 27568
rect 10414 27512 10470 27548
rect 9857 26682 9913 26684
rect 9937 26682 9993 26684
rect 10017 26682 10073 26684
rect 10097 26682 10153 26684
rect 9857 26630 9903 26682
rect 9903 26630 9913 26682
rect 9937 26630 9967 26682
rect 9967 26630 9979 26682
rect 9979 26630 9993 26682
rect 10017 26630 10031 26682
rect 10031 26630 10043 26682
rect 10043 26630 10073 26682
rect 10097 26630 10107 26682
rect 10107 26630 10153 26682
rect 9857 26628 9913 26630
rect 9937 26628 9993 26630
rect 10017 26628 10073 26630
rect 10097 26628 10153 26630
rect 10046 26016 10102 26072
rect 9494 24792 9550 24848
rect 9862 25744 9918 25800
rect 10322 26288 10378 26344
rect 9857 25594 9913 25596
rect 9937 25594 9993 25596
rect 10017 25594 10073 25596
rect 10097 25594 10153 25596
rect 9857 25542 9903 25594
rect 9903 25542 9913 25594
rect 9937 25542 9967 25594
rect 9967 25542 9979 25594
rect 9979 25542 9993 25594
rect 10017 25542 10031 25594
rect 10031 25542 10043 25594
rect 10043 25542 10073 25594
rect 10097 25542 10107 25594
rect 10107 25542 10153 25594
rect 9857 25540 9913 25542
rect 9937 25540 9993 25542
rect 10017 25540 10073 25542
rect 10097 25540 10153 25542
rect 9857 24506 9913 24508
rect 9937 24506 9993 24508
rect 10017 24506 10073 24508
rect 10097 24506 10153 24508
rect 9857 24454 9903 24506
rect 9903 24454 9913 24506
rect 9937 24454 9967 24506
rect 9967 24454 9979 24506
rect 9979 24454 9993 24506
rect 10017 24454 10031 24506
rect 10031 24454 10043 24506
rect 10043 24454 10073 24506
rect 10097 24454 10107 24506
rect 10107 24454 10153 24506
rect 9857 24452 9913 24454
rect 9937 24452 9993 24454
rect 10017 24452 10073 24454
rect 10097 24452 10153 24454
rect 10322 25336 10378 25392
rect 9586 23976 9642 24032
rect 9586 23724 9642 23760
rect 9586 23704 9588 23724
rect 9588 23704 9640 23724
rect 9640 23704 9642 23724
rect 9770 23860 9826 23896
rect 9770 23840 9772 23860
rect 9772 23840 9824 23860
rect 9824 23840 9826 23860
rect 9770 23724 9826 23760
rect 9770 23704 9772 23724
rect 9772 23704 9824 23724
rect 9824 23704 9826 23724
rect 10138 23588 10194 23624
rect 9678 23432 9734 23488
rect 9586 22208 9642 22264
rect 10138 23568 10140 23588
rect 10140 23568 10192 23588
rect 10192 23568 10194 23588
rect 9857 23418 9913 23420
rect 9937 23418 9993 23420
rect 10017 23418 10073 23420
rect 10097 23418 10153 23420
rect 9857 23366 9903 23418
rect 9903 23366 9913 23418
rect 9937 23366 9967 23418
rect 9967 23366 9979 23418
rect 9979 23366 9993 23418
rect 10017 23366 10031 23418
rect 10031 23366 10043 23418
rect 10043 23366 10073 23418
rect 10097 23366 10107 23418
rect 10107 23366 10153 23418
rect 9857 23364 9913 23366
rect 9937 23364 9993 23366
rect 10017 23364 10073 23366
rect 10097 23364 10153 23366
rect 10138 23160 10194 23216
rect 9857 22330 9913 22332
rect 9937 22330 9993 22332
rect 10017 22330 10073 22332
rect 10097 22330 10153 22332
rect 9857 22278 9903 22330
rect 9903 22278 9913 22330
rect 9937 22278 9967 22330
rect 9967 22278 9979 22330
rect 9979 22278 9993 22330
rect 10017 22278 10031 22330
rect 10031 22278 10043 22330
rect 10043 22278 10073 22330
rect 10097 22278 10107 22330
rect 10107 22278 10153 22330
rect 9857 22276 9913 22278
rect 9937 22276 9993 22278
rect 10017 22276 10073 22278
rect 10097 22276 10153 22278
rect 9862 21528 9918 21584
rect 9586 21120 9642 21176
rect 9857 21242 9913 21244
rect 9937 21242 9993 21244
rect 10017 21242 10073 21244
rect 10097 21242 10153 21244
rect 9857 21190 9903 21242
rect 9903 21190 9913 21242
rect 9937 21190 9967 21242
rect 9967 21190 9979 21242
rect 9979 21190 9993 21242
rect 10017 21190 10031 21242
rect 10031 21190 10043 21242
rect 10043 21190 10073 21242
rect 10097 21190 10107 21242
rect 10107 21190 10153 21242
rect 9857 21188 9913 21190
rect 9937 21188 9993 21190
rect 10017 21188 10073 21190
rect 10097 21188 10153 21190
rect 9770 20576 9826 20632
rect 8942 12688 8998 12744
rect 9857 20154 9913 20156
rect 9937 20154 9993 20156
rect 10017 20154 10073 20156
rect 10097 20154 10153 20156
rect 9857 20102 9903 20154
rect 9903 20102 9913 20154
rect 9937 20102 9967 20154
rect 9967 20102 9979 20154
rect 9979 20102 9993 20154
rect 10017 20102 10031 20154
rect 10031 20102 10043 20154
rect 10043 20102 10073 20154
rect 10097 20102 10107 20154
rect 10107 20102 10153 20154
rect 9857 20100 9913 20102
rect 9937 20100 9993 20102
rect 10017 20100 10073 20102
rect 10097 20100 10153 20102
rect 9494 18264 9550 18320
rect 9857 19066 9913 19068
rect 9937 19066 9993 19068
rect 10017 19066 10073 19068
rect 10097 19066 10153 19068
rect 9857 19014 9903 19066
rect 9903 19014 9913 19066
rect 9937 19014 9967 19066
rect 9967 19014 9979 19066
rect 9979 19014 9993 19066
rect 10017 19014 10031 19066
rect 10031 19014 10043 19066
rect 10043 19014 10073 19066
rect 10097 19014 10107 19066
rect 10107 19014 10153 19066
rect 9857 19012 9913 19014
rect 9937 19012 9993 19014
rect 10017 19012 10073 19014
rect 10097 19012 10153 19014
rect 9862 18808 9918 18864
rect 10046 18536 10102 18592
rect 10690 29300 10746 29336
rect 10690 29280 10692 29300
rect 10692 29280 10744 29300
rect 10744 29280 10746 29300
rect 10690 24656 10746 24712
rect 10598 20984 10654 21040
rect 10322 19372 10378 19408
rect 10322 19352 10324 19372
rect 10324 19352 10376 19372
rect 10376 19352 10378 19372
rect 9857 17978 9913 17980
rect 9937 17978 9993 17980
rect 10017 17978 10073 17980
rect 10097 17978 10153 17980
rect 9857 17926 9903 17978
rect 9903 17926 9913 17978
rect 9937 17926 9967 17978
rect 9967 17926 9979 17978
rect 9979 17926 9993 17978
rect 10017 17926 10031 17978
rect 10031 17926 10043 17978
rect 10043 17926 10073 17978
rect 10097 17926 10107 17978
rect 10107 17926 10153 17978
rect 9857 17924 9913 17926
rect 9937 17924 9993 17926
rect 10017 17924 10073 17926
rect 10097 17924 10153 17926
rect 10598 18672 10654 18728
rect 9857 16890 9913 16892
rect 9937 16890 9993 16892
rect 10017 16890 10073 16892
rect 10097 16890 10153 16892
rect 9857 16838 9903 16890
rect 9903 16838 9913 16890
rect 9937 16838 9967 16890
rect 9967 16838 9979 16890
rect 9979 16838 9993 16890
rect 10017 16838 10031 16890
rect 10031 16838 10043 16890
rect 10043 16838 10073 16890
rect 10097 16838 10107 16890
rect 10107 16838 10153 16890
rect 9857 16836 9913 16838
rect 9937 16836 9993 16838
rect 10017 16836 10073 16838
rect 10097 16836 10153 16838
rect 9770 16496 9826 16552
rect 9034 11056 9090 11112
rect 9857 15802 9913 15804
rect 9937 15802 9993 15804
rect 10017 15802 10073 15804
rect 10097 15802 10153 15804
rect 9857 15750 9903 15802
rect 9903 15750 9913 15802
rect 9937 15750 9967 15802
rect 9967 15750 9979 15802
rect 9979 15750 9993 15802
rect 10017 15750 10031 15802
rect 10031 15750 10043 15802
rect 10043 15750 10073 15802
rect 10097 15750 10107 15802
rect 10107 15750 10153 15802
rect 9857 15748 9913 15750
rect 9937 15748 9993 15750
rect 10017 15748 10073 15750
rect 10097 15748 10153 15750
rect 9862 15544 9918 15600
rect 9857 14714 9913 14716
rect 9937 14714 9993 14716
rect 10017 14714 10073 14716
rect 10097 14714 10153 14716
rect 9857 14662 9903 14714
rect 9903 14662 9913 14714
rect 9937 14662 9967 14714
rect 9967 14662 9979 14714
rect 9979 14662 9993 14714
rect 10017 14662 10031 14714
rect 10031 14662 10043 14714
rect 10043 14662 10073 14714
rect 10097 14662 10107 14714
rect 10107 14662 10153 14714
rect 9857 14660 9913 14662
rect 9937 14660 9993 14662
rect 10017 14660 10073 14662
rect 10097 14660 10153 14662
rect 9857 13626 9913 13628
rect 9937 13626 9993 13628
rect 10017 13626 10073 13628
rect 10097 13626 10153 13628
rect 9857 13574 9903 13626
rect 9903 13574 9913 13626
rect 9937 13574 9967 13626
rect 9967 13574 9979 13626
rect 9979 13574 9993 13626
rect 10017 13574 10031 13626
rect 10031 13574 10043 13626
rect 10043 13574 10073 13626
rect 10097 13574 10107 13626
rect 10107 13574 10153 13626
rect 9857 13572 9913 13574
rect 9937 13572 9993 13574
rect 10017 13572 10073 13574
rect 10097 13572 10153 13574
rect 10414 17040 10470 17096
rect 10598 13640 10654 13696
rect 9857 12538 9913 12540
rect 9937 12538 9993 12540
rect 10017 12538 10073 12540
rect 10097 12538 10153 12540
rect 9857 12486 9903 12538
rect 9903 12486 9913 12538
rect 9937 12486 9967 12538
rect 9967 12486 9979 12538
rect 9979 12486 9993 12538
rect 10017 12486 10031 12538
rect 10031 12486 10043 12538
rect 10043 12486 10073 12538
rect 10097 12486 10107 12538
rect 10107 12486 10153 12538
rect 9857 12484 9913 12486
rect 9937 12484 9993 12486
rect 10017 12484 10073 12486
rect 10097 12484 10153 12486
rect 9857 11450 9913 11452
rect 9937 11450 9993 11452
rect 10017 11450 10073 11452
rect 10097 11450 10153 11452
rect 9857 11398 9903 11450
rect 9903 11398 9913 11450
rect 9937 11398 9967 11450
rect 9967 11398 9979 11450
rect 9979 11398 9993 11450
rect 10017 11398 10031 11450
rect 10031 11398 10043 11450
rect 10043 11398 10073 11450
rect 10097 11398 10107 11450
rect 10107 11398 10153 11450
rect 9857 11396 9913 11398
rect 9937 11396 9993 11398
rect 10017 11396 10073 11398
rect 10097 11396 10153 11398
rect 9494 10920 9550 10976
rect 9310 6704 9366 6760
rect 10046 11056 10102 11112
rect 9310 5888 9366 5944
rect 9678 8472 9734 8528
rect 9857 10362 9913 10364
rect 9937 10362 9993 10364
rect 10017 10362 10073 10364
rect 10097 10362 10153 10364
rect 9857 10310 9903 10362
rect 9903 10310 9913 10362
rect 9937 10310 9967 10362
rect 9967 10310 9979 10362
rect 9979 10310 9993 10362
rect 10017 10310 10031 10362
rect 10031 10310 10043 10362
rect 10043 10310 10073 10362
rect 10097 10310 10107 10362
rect 10107 10310 10153 10362
rect 9857 10308 9913 10310
rect 9937 10308 9993 10310
rect 10017 10308 10073 10310
rect 10097 10308 10153 10310
rect 10414 12688 10470 12744
rect 11242 32952 11298 33008
rect 11242 31048 11298 31104
rect 11058 29416 11114 29472
rect 11610 35284 11666 35320
rect 11610 35264 11612 35284
rect 11612 35264 11664 35284
rect 11664 35264 11666 35284
rect 11610 34448 11666 34504
rect 11794 35536 11850 35592
rect 11794 34856 11850 34912
rect 11702 34040 11758 34096
rect 11518 32680 11574 32736
rect 10874 29008 10930 29064
rect 11058 29008 11114 29064
rect 11150 28328 11206 28384
rect 10966 25880 11022 25936
rect 10874 24248 10930 24304
rect 11518 28192 11574 28248
rect 11518 27648 11574 27704
rect 10874 21528 10930 21584
rect 10874 14864 10930 14920
rect 10966 14592 11022 14648
rect 9857 9274 9913 9276
rect 9937 9274 9993 9276
rect 10017 9274 10073 9276
rect 10097 9274 10153 9276
rect 9857 9222 9903 9274
rect 9903 9222 9913 9274
rect 9937 9222 9967 9274
rect 9967 9222 9979 9274
rect 9979 9222 9993 9274
rect 10017 9222 10031 9274
rect 10031 9222 10043 9274
rect 10043 9222 10073 9274
rect 10097 9222 10107 9274
rect 10107 9222 10153 9274
rect 9857 9220 9913 9222
rect 9937 9220 9993 9222
rect 10017 9220 10073 9222
rect 10097 9220 10153 9222
rect 9857 8186 9913 8188
rect 9937 8186 9993 8188
rect 10017 8186 10073 8188
rect 10097 8186 10153 8188
rect 9857 8134 9903 8186
rect 9903 8134 9913 8186
rect 9937 8134 9967 8186
rect 9967 8134 9979 8186
rect 9979 8134 9993 8186
rect 10017 8134 10031 8186
rect 10031 8134 10043 8186
rect 10043 8134 10073 8186
rect 10097 8134 10107 8186
rect 10107 8134 10153 8186
rect 9857 8132 9913 8134
rect 9937 8132 9993 8134
rect 10017 8132 10073 8134
rect 10097 8132 10153 8134
rect 9857 7098 9913 7100
rect 9937 7098 9993 7100
rect 10017 7098 10073 7100
rect 10097 7098 10153 7100
rect 9857 7046 9903 7098
rect 9903 7046 9913 7098
rect 9937 7046 9967 7098
rect 9967 7046 9979 7098
rect 9979 7046 9993 7098
rect 10017 7046 10031 7098
rect 10031 7046 10043 7098
rect 10043 7046 10073 7098
rect 10097 7046 10107 7098
rect 10107 7046 10153 7098
rect 9857 7044 9913 7046
rect 9937 7044 9993 7046
rect 10017 7044 10073 7046
rect 10097 7044 10153 7046
rect 9310 5480 9366 5536
rect 9126 3304 9182 3360
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 10046 5652 10048 5672
rect 10048 5652 10100 5672
rect 10100 5652 10102 5672
rect 10046 5616 10102 5652
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 11058 8880 11114 8936
rect 10230 4120 10286 4176
rect 10138 3984 10194 4040
rect 9494 3732 9550 3768
rect 9494 3712 9496 3732
rect 9496 3712 9548 3732
rect 9548 3712 9550 3732
rect 6550 1264 6606 1320
rect 6734 1164 6736 1184
rect 6736 1164 6788 1184
rect 6788 1164 6790 1184
rect 6734 1128 6790 1164
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 7746 2216 7802 2272
rect 7654 2080 7710 2136
rect 7930 1300 7932 1320
rect 7932 1300 7984 1320
rect 7984 1300 7986 1320
rect 7930 1264 7986 1300
rect 8482 2352 8538 2408
rect 8114 2216 8170 2272
rect 8390 2216 8446 2272
rect 8666 1264 8722 1320
rect 8850 2216 8906 2272
rect 9218 2352 9274 2408
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 9770 3440 9826 3496
rect 9954 3168 10010 3224
rect 9494 2644 9550 2680
rect 9494 2624 9496 2644
rect 9496 2624 9548 2644
rect 9548 2624 9550 2644
rect 10138 3304 10194 3360
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 9678 1844 9680 1864
rect 9680 1844 9732 1864
rect 9732 1844 9734 1864
rect 9678 1808 9734 1844
rect 10966 7928 11022 7984
rect 12162 32852 12164 32872
rect 12164 32852 12216 32872
rect 12216 32852 12218 32872
rect 12162 32816 12218 32852
rect 12070 30640 12126 30696
rect 11886 28736 11942 28792
rect 11610 24928 11666 24984
rect 11702 23704 11758 23760
rect 11242 20032 11298 20088
rect 11426 20460 11482 20496
rect 11426 20440 11428 20460
rect 11428 20440 11480 20460
rect 11480 20440 11482 20460
rect 11794 22480 11850 22536
rect 11702 22072 11758 22128
rect 12346 37168 12402 37224
rect 12346 34856 12402 34912
rect 12824 42458 12880 42460
rect 12904 42458 12960 42460
rect 12984 42458 13040 42460
rect 13064 42458 13120 42460
rect 12824 42406 12870 42458
rect 12870 42406 12880 42458
rect 12904 42406 12934 42458
rect 12934 42406 12946 42458
rect 12946 42406 12960 42458
rect 12984 42406 12998 42458
rect 12998 42406 13010 42458
rect 13010 42406 13040 42458
rect 13064 42406 13074 42458
rect 13074 42406 13120 42458
rect 12824 42404 12880 42406
rect 12904 42404 12960 42406
rect 12984 42404 13040 42406
rect 13064 42404 13120 42406
rect 12824 41370 12880 41372
rect 12904 41370 12960 41372
rect 12984 41370 13040 41372
rect 13064 41370 13120 41372
rect 12824 41318 12870 41370
rect 12870 41318 12880 41370
rect 12904 41318 12934 41370
rect 12934 41318 12946 41370
rect 12946 41318 12960 41370
rect 12984 41318 12998 41370
rect 12998 41318 13010 41370
rect 13010 41318 13040 41370
rect 13064 41318 13074 41370
rect 13074 41318 13120 41370
rect 12824 41316 12880 41318
rect 12904 41316 12960 41318
rect 12984 41316 13040 41318
rect 13064 41316 13120 41318
rect 12824 40282 12880 40284
rect 12904 40282 12960 40284
rect 12984 40282 13040 40284
rect 13064 40282 13120 40284
rect 12824 40230 12870 40282
rect 12870 40230 12880 40282
rect 12904 40230 12934 40282
rect 12934 40230 12946 40282
rect 12946 40230 12960 40282
rect 12984 40230 12998 40282
rect 12998 40230 13010 40282
rect 13010 40230 13040 40282
rect 13064 40230 13074 40282
rect 13074 40230 13120 40282
rect 12824 40228 12880 40230
rect 12904 40228 12960 40230
rect 12984 40228 13040 40230
rect 13064 40228 13120 40230
rect 12824 39194 12880 39196
rect 12904 39194 12960 39196
rect 12984 39194 13040 39196
rect 13064 39194 13120 39196
rect 12824 39142 12870 39194
rect 12870 39142 12880 39194
rect 12904 39142 12934 39194
rect 12934 39142 12946 39194
rect 12946 39142 12960 39194
rect 12984 39142 12998 39194
rect 12998 39142 13010 39194
rect 13010 39142 13040 39194
rect 13064 39142 13074 39194
rect 13074 39142 13120 39194
rect 12824 39140 12880 39142
rect 12904 39140 12960 39142
rect 12984 39140 13040 39142
rect 13064 39140 13120 39142
rect 12622 33360 12678 33416
rect 12530 33224 12586 33280
rect 12824 38106 12880 38108
rect 12904 38106 12960 38108
rect 12984 38106 13040 38108
rect 13064 38106 13120 38108
rect 12824 38054 12870 38106
rect 12870 38054 12880 38106
rect 12904 38054 12934 38106
rect 12934 38054 12946 38106
rect 12946 38054 12960 38106
rect 12984 38054 12998 38106
rect 12998 38054 13010 38106
rect 13010 38054 13040 38106
rect 13064 38054 13074 38106
rect 13074 38054 13120 38106
rect 12824 38052 12880 38054
rect 12904 38052 12960 38054
rect 12984 38052 13040 38054
rect 13064 38052 13120 38054
rect 12824 37018 12880 37020
rect 12904 37018 12960 37020
rect 12984 37018 13040 37020
rect 13064 37018 13120 37020
rect 12824 36966 12870 37018
rect 12870 36966 12880 37018
rect 12904 36966 12934 37018
rect 12934 36966 12946 37018
rect 12946 36966 12960 37018
rect 12984 36966 12998 37018
rect 12998 36966 13010 37018
rect 13010 36966 13040 37018
rect 13064 36966 13074 37018
rect 13074 36966 13120 37018
rect 12824 36964 12880 36966
rect 12904 36964 12960 36966
rect 12984 36964 13040 36966
rect 13064 36964 13120 36966
rect 13818 42880 13874 42936
rect 14278 42880 14334 42936
rect 14922 42880 14978 42936
rect 14094 40568 14150 40624
rect 12824 35930 12880 35932
rect 12904 35930 12960 35932
rect 12984 35930 13040 35932
rect 13064 35930 13120 35932
rect 12824 35878 12870 35930
rect 12870 35878 12880 35930
rect 12904 35878 12934 35930
rect 12934 35878 12946 35930
rect 12946 35878 12960 35930
rect 12984 35878 12998 35930
rect 12998 35878 13010 35930
rect 13010 35878 13040 35930
rect 13064 35878 13074 35930
rect 13074 35878 13120 35930
rect 12824 35876 12880 35878
rect 12904 35876 12960 35878
rect 12984 35876 13040 35878
rect 13064 35876 13120 35878
rect 13174 35128 13230 35184
rect 12990 34992 13046 35048
rect 12824 34842 12880 34844
rect 12904 34842 12960 34844
rect 12984 34842 13040 34844
rect 13064 34842 13120 34844
rect 12824 34790 12870 34842
rect 12870 34790 12880 34842
rect 12904 34790 12934 34842
rect 12934 34790 12946 34842
rect 12946 34790 12960 34842
rect 12984 34790 12998 34842
rect 12998 34790 13010 34842
rect 13010 34790 13040 34842
rect 13064 34790 13074 34842
rect 13074 34790 13120 34842
rect 12824 34788 12880 34790
rect 12904 34788 12960 34790
rect 12984 34788 13040 34790
rect 13064 34788 13120 34790
rect 13266 34584 13322 34640
rect 12824 33754 12880 33756
rect 12904 33754 12960 33756
rect 12984 33754 13040 33756
rect 13064 33754 13120 33756
rect 12824 33702 12870 33754
rect 12870 33702 12880 33754
rect 12904 33702 12934 33754
rect 12934 33702 12946 33754
rect 12946 33702 12960 33754
rect 12984 33702 12998 33754
rect 12998 33702 13010 33754
rect 13010 33702 13040 33754
rect 13064 33702 13074 33754
rect 13074 33702 13120 33754
rect 12824 33700 12880 33702
rect 12904 33700 12960 33702
rect 12984 33700 13040 33702
rect 13064 33700 13120 33702
rect 12824 32666 12880 32668
rect 12904 32666 12960 32668
rect 12984 32666 13040 32668
rect 13064 32666 13120 32668
rect 12824 32614 12870 32666
rect 12870 32614 12880 32666
rect 12904 32614 12934 32666
rect 12934 32614 12946 32666
rect 12946 32614 12960 32666
rect 12984 32614 12998 32666
rect 12998 32614 13010 32666
rect 13010 32614 13040 32666
rect 13064 32614 13074 32666
rect 13074 32614 13120 32666
rect 12824 32612 12880 32614
rect 12904 32612 12960 32614
rect 12984 32612 13040 32614
rect 13064 32612 13120 32614
rect 12438 31456 12494 31512
rect 12346 27648 12402 27704
rect 12254 27512 12310 27568
rect 12346 23976 12402 24032
rect 12254 23432 12310 23488
rect 11610 18944 11666 19000
rect 11242 12824 11298 12880
rect 10506 3712 10562 3768
rect 10506 3440 10562 3496
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 10690 3984 10746 4040
rect 11058 5480 11114 5536
rect 10874 3168 10930 3224
rect 11058 2896 11114 2952
rect 11518 15136 11574 15192
rect 11886 18808 11942 18864
rect 11794 18300 11796 18320
rect 11796 18300 11848 18320
rect 11848 18300 11850 18320
rect 11794 18264 11850 18300
rect 11610 13912 11666 13968
rect 11886 14340 11942 14376
rect 11886 14320 11888 14340
rect 11888 14320 11940 14340
rect 11940 14320 11942 14340
rect 12254 17196 12310 17232
rect 12254 17176 12256 17196
rect 12256 17176 12308 17196
rect 12308 17176 12310 17196
rect 12622 31728 12678 31784
rect 12824 31578 12880 31580
rect 12904 31578 12960 31580
rect 12984 31578 13040 31580
rect 13064 31578 13120 31580
rect 12824 31526 12870 31578
rect 12870 31526 12880 31578
rect 12904 31526 12934 31578
rect 12934 31526 12946 31578
rect 12946 31526 12960 31578
rect 12984 31526 12998 31578
rect 12998 31526 13010 31578
rect 13010 31526 13040 31578
rect 13064 31526 13074 31578
rect 13074 31526 13120 31578
rect 12824 31524 12880 31526
rect 12904 31524 12960 31526
rect 12984 31524 13040 31526
rect 13064 31524 13120 31526
rect 12824 30490 12880 30492
rect 12904 30490 12960 30492
rect 12984 30490 13040 30492
rect 13064 30490 13120 30492
rect 12824 30438 12870 30490
rect 12870 30438 12880 30490
rect 12904 30438 12934 30490
rect 12934 30438 12946 30490
rect 12946 30438 12960 30490
rect 12984 30438 12998 30490
rect 12998 30438 13010 30490
rect 13010 30438 13040 30490
rect 13064 30438 13074 30490
rect 13074 30438 13120 30490
rect 12824 30436 12880 30438
rect 12904 30436 12960 30438
rect 12984 30436 13040 30438
rect 13064 30436 13120 30438
rect 12714 29588 12716 29608
rect 12716 29588 12768 29608
rect 12768 29588 12770 29608
rect 12714 29552 12770 29588
rect 12824 29402 12880 29404
rect 12904 29402 12960 29404
rect 12984 29402 13040 29404
rect 13064 29402 13120 29404
rect 12824 29350 12870 29402
rect 12870 29350 12880 29402
rect 12904 29350 12934 29402
rect 12934 29350 12946 29402
rect 12946 29350 12960 29402
rect 12984 29350 12998 29402
rect 12998 29350 13010 29402
rect 13010 29350 13040 29402
rect 13064 29350 13074 29402
rect 13074 29350 13120 29402
rect 12824 29348 12880 29350
rect 12904 29348 12960 29350
rect 12984 29348 13040 29350
rect 13064 29348 13120 29350
rect 12824 28314 12880 28316
rect 12904 28314 12960 28316
rect 12984 28314 13040 28316
rect 13064 28314 13120 28316
rect 12824 28262 12870 28314
rect 12870 28262 12880 28314
rect 12904 28262 12934 28314
rect 12934 28262 12946 28314
rect 12946 28262 12960 28314
rect 12984 28262 12998 28314
rect 12998 28262 13010 28314
rect 13010 28262 13040 28314
rect 13064 28262 13074 28314
rect 13074 28262 13120 28314
rect 12824 28260 12880 28262
rect 12904 28260 12960 28262
rect 12984 28260 13040 28262
rect 13064 28260 13120 28262
rect 12824 27226 12880 27228
rect 12904 27226 12960 27228
rect 12984 27226 13040 27228
rect 13064 27226 13120 27228
rect 12824 27174 12870 27226
rect 12870 27174 12880 27226
rect 12904 27174 12934 27226
rect 12934 27174 12946 27226
rect 12946 27174 12960 27226
rect 12984 27174 12998 27226
rect 12998 27174 13010 27226
rect 13010 27174 13040 27226
rect 13064 27174 13074 27226
rect 13074 27174 13120 27226
rect 12824 27172 12880 27174
rect 12904 27172 12960 27174
rect 12984 27172 13040 27174
rect 13064 27172 13120 27174
rect 13542 35400 13598 35456
rect 13726 33496 13782 33552
rect 13634 31864 13690 31920
rect 13266 26696 13322 26752
rect 12824 26138 12880 26140
rect 12904 26138 12960 26140
rect 12984 26138 13040 26140
rect 13064 26138 13120 26140
rect 12824 26086 12870 26138
rect 12870 26086 12880 26138
rect 12904 26086 12934 26138
rect 12934 26086 12946 26138
rect 12946 26086 12960 26138
rect 12984 26086 12998 26138
rect 12998 26086 13010 26138
rect 13010 26086 13040 26138
rect 13064 26086 13074 26138
rect 13074 26086 13120 26138
rect 12824 26084 12880 26086
rect 12904 26084 12960 26086
rect 12984 26084 13040 26086
rect 13064 26084 13120 26086
rect 12824 25050 12880 25052
rect 12904 25050 12960 25052
rect 12984 25050 13040 25052
rect 13064 25050 13120 25052
rect 12824 24998 12870 25050
rect 12870 24998 12880 25050
rect 12904 24998 12934 25050
rect 12934 24998 12946 25050
rect 12946 24998 12960 25050
rect 12984 24998 12998 25050
rect 12998 24998 13010 25050
rect 13010 24998 13040 25050
rect 13064 24998 13074 25050
rect 13074 24998 13120 25050
rect 12824 24996 12880 24998
rect 12904 24996 12960 24998
rect 12984 24996 13040 24998
rect 13064 24996 13120 24998
rect 12824 23962 12880 23964
rect 12904 23962 12960 23964
rect 12984 23962 13040 23964
rect 13064 23962 13120 23964
rect 12824 23910 12870 23962
rect 12870 23910 12880 23962
rect 12904 23910 12934 23962
rect 12934 23910 12946 23962
rect 12946 23910 12960 23962
rect 12984 23910 12998 23962
rect 12998 23910 13010 23962
rect 13010 23910 13040 23962
rect 13064 23910 13074 23962
rect 13074 23910 13120 23962
rect 12824 23908 12880 23910
rect 12904 23908 12960 23910
rect 12984 23908 13040 23910
rect 13064 23908 13120 23910
rect 12530 21120 12586 21176
rect 12438 17856 12494 17912
rect 12254 15408 12310 15464
rect 11886 12688 11942 12744
rect 12162 13776 12218 13832
rect 11702 10648 11758 10704
rect 11886 9424 11942 9480
rect 11794 8336 11850 8392
rect 11794 8200 11850 8256
rect 11518 5888 11574 5944
rect 11426 4528 11482 4584
rect 14370 35264 14426 35320
rect 14186 32544 14242 32600
rect 14094 29688 14150 29744
rect 13634 28056 13690 28112
rect 13818 28328 13874 28384
rect 13542 26424 13598 26480
rect 13450 25880 13506 25936
rect 12824 22874 12880 22876
rect 12904 22874 12960 22876
rect 12984 22874 13040 22876
rect 13064 22874 13120 22876
rect 12824 22822 12870 22874
rect 12870 22822 12880 22874
rect 12904 22822 12934 22874
rect 12934 22822 12946 22874
rect 12946 22822 12960 22874
rect 12984 22822 12998 22874
rect 12998 22822 13010 22874
rect 13010 22822 13040 22874
rect 13064 22822 13074 22874
rect 13074 22822 13120 22874
rect 12824 22820 12880 22822
rect 12904 22820 12960 22822
rect 12984 22820 13040 22822
rect 13064 22820 13120 22822
rect 12824 21786 12880 21788
rect 12904 21786 12960 21788
rect 12984 21786 13040 21788
rect 13064 21786 13120 21788
rect 12824 21734 12870 21786
rect 12870 21734 12880 21786
rect 12904 21734 12934 21786
rect 12934 21734 12946 21786
rect 12946 21734 12960 21786
rect 12984 21734 12998 21786
rect 12998 21734 13010 21786
rect 13010 21734 13040 21786
rect 13064 21734 13074 21786
rect 13074 21734 13120 21786
rect 12824 21732 12880 21734
rect 12904 21732 12960 21734
rect 12984 21732 13040 21734
rect 13064 21732 13120 21734
rect 12824 20698 12880 20700
rect 12904 20698 12960 20700
rect 12984 20698 13040 20700
rect 13064 20698 13120 20700
rect 12824 20646 12870 20698
rect 12870 20646 12880 20698
rect 12904 20646 12934 20698
rect 12934 20646 12946 20698
rect 12946 20646 12960 20698
rect 12984 20646 12998 20698
rect 12998 20646 13010 20698
rect 13010 20646 13040 20698
rect 13064 20646 13074 20698
rect 13074 20646 13120 20698
rect 12824 20644 12880 20646
rect 12904 20644 12960 20646
rect 12984 20644 13040 20646
rect 13064 20644 13120 20646
rect 12714 19796 12716 19816
rect 12716 19796 12768 19816
rect 12768 19796 12770 19816
rect 12714 19760 12770 19796
rect 12824 19610 12880 19612
rect 12904 19610 12960 19612
rect 12984 19610 13040 19612
rect 13064 19610 13120 19612
rect 12824 19558 12870 19610
rect 12870 19558 12880 19610
rect 12904 19558 12934 19610
rect 12934 19558 12946 19610
rect 12946 19558 12960 19610
rect 12984 19558 12998 19610
rect 12998 19558 13010 19610
rect 13010 19558 13040 19610
rect 13064 19558 13074 19610
rect 13074 19558 13120 19610
rect 12824 19556 12880 19558
rect 12904 19556 12960 19558
rect 12984 19556 13040 19558
rect 13064 19556 13120 19558
rect 12824 18522 12880 18524
rect 12904 18522 12960 18524
rect 12984 18522 13040 18524
rect 13064 18522 13120 18524
rect 12824 18470 12870 18522
rect 12870 18470 12880 18522
rect 12904 18470 12934 18522
rect 12934 18470 12946 18522
rect 12946 18470 12960 18522
rect 12984 18470 12998 18522
rect 12998 18470 13010 18522
rect 13010 18470 13040 18522
rect 13064 18470 13074 18522
rect 13074 18470 13120 18522
rect 12824 18468 12880 18470
rect 12904 18468 12960 18470
rect 12984 18468 13040 18470
rect 13064 18468 13120 18470
rect 12824 17434 12880 17436
rect 12904 17434 12960 17436
rect 12984 17434 13040 17436
rect 13064 17434 13120 17436
rect 12824 17382 12870 17434
rect 12870 17382 12880 17434
rect 12904 17382 12934 17434
rect 12934 17382 12946 17434
rect 12946 17382 12960 17434
rect 12984 17382 12998 17434
rect 12998 17382 13010 17434
rect 13010 17382 13040 17434
rect 13064 17382 13074 17434
rect 13074 17382 13120 17434
rect 12824 17380 12880 17382
rect 12904 17380 12960 17382
rect 12984 17380 13040 17382
rect 13064 17380 13120 17382
rect 12824 16346 12880 16348
rect 12904 16346 12960 16348
rect 12984 16346 13040 16348
rect 13064 16346 13120 16348
rect 12824 16294 12870 16346
rect 12870 16294 12880 16346
rect 12904 16294 12934 16346
rect 12934 16294 12946 16346
rect 12946 16294 12960 16346
rect 12984 16294 12998 16346
rect 12998 16294 13010 16346
rect 13010 16294 13040 16346
rect 13064 16294 13074 16346
rect 13074 16294 13120 16346
rect 12824 16292 12880 16294
rect 12904 16292 12960 16294
rect 12984 16292 13040 16294
rect 13064 16292 13120 16294
rect 12438 13232 12494 13288
rect 12824 15258 12880 15260
rect 12904 15258 12960 15260
rect 12984 15258 13040 15260
rect 13064 15258 13120 15260
rect 12824 15206 12870 15258
rect 12870 15206 12880 15258
rect 12904 15206 12934 15258
rect 12934 15206 12946 15258
rect 12946 15206 12960 15258
rect 12984 15206 12998 15258
rect 12998 15206 13010 15258
rect 13010 15206 13040 15258
rect 13064 15206 13074 15258
rect 13074 15206 13120 15258
rect 12824 15204 12880 15206
rect 12904 15204 12960 15206
rect 12984 15204 13040 15206
rect 13064 15204 13120 15206
rect 13542 23160 13598 23216
rect 13542 22888 13598 22944
rect 13450 21120 13506 21176
rect 13358 17856 13414 17912
rect 12824 14170 12880 14172
rect 12904 14170 12960 14172
rect 12984 14170 13040 14172
rect 13064 14170 13120 14172
rect 12824 14118 12870 14170
rect 12870 14118 12880 14170
rect 12904 14118 12934 14170
rect 12934 14118 12946 14170
rect 12946 14118 12960 14170
rect 12984 14118 12998 14170
rect 12998 14118 13010 14170
rect 13010 14118 13040 14170
rect 13064 14118 13074 14170
rect 13074 14118 13120 14170
rect 12824 14116 12880 14118
rect 12904 14116 12960 14118
rect 12984 14116 13040 14118
rect 13064 14116 13120 14118
rect 12824 13082 12880 13084
rect 12904 13082 12960 13084
rect 12984 13082 13040 13084
rect 13064 13082 13120 13084
rect 12824 13030 12870 13082
rect 12870 13030 12880 13082
rect 12904 13030 12934 13082
rect 12934 13030 12946 13082
rect 12946 13030 12960 13082
rect 12984 13030 12998 13082
rect 12998 13030 13010 13082
rect 13010 13030 13040 13082
rect 13064 13030 13074 13082
rect 13074 13030 13120 13082
rect 12824 13028 12880 13030
rect 12904 13028 12960 13030
rect 12984 13028 13040 13030
rect 13064 13028 13120 13030
rect 12254 9696 12310 9752
rect 12162 7248 12218 7304
rect 12162 5752 12218 5808
rect 12162 4936 12218 4992
rect 12824 11994 12880 11996
rect 12904 11994 12960 11996
rect 12984 11994 13040 11996
rect 13064 11994 13120 11996
rect 12824 11942 12870 11994
rect 12870 11942 12880 11994
rect 12904 11942 12934 11994
rect 12934 11942 12946 11994
rect 12946 11942 12960 11994
rect 12984 11942 12998 11994
rect 12998 11942 13010 11994
rect 13010 11942 13040 11994
rect 13064 11942 13074 11994
rect 13074 11942 13120 11994
rect 12824 11940 12880 11942
rect 12904 11940 12960 11942
rect 12984 11940 13040 11942
rect 13064 11940 13120 11942
rect 12824 10906 12880 10908
rect 12904 10906 12960 10908
rect 12984 10906 13040 10908
rect 13064 10906 13120 10908
rect 12824 10854 12870 10906
rect 12870 10854 12880 10906
rect 12904 10854 12934 10906
rect 12934 10854 12946 10906
rect 12946 10854 12960 10906
rect 12984 10854 12998 10906
rect 12998 10854 13010 10906
rect 13010 10854 13040 10906
rect 13064 10854 13074 10906
rect 13074 10854 13120 10906
rect 12824 10852 12880 10854
rect 12904 10852 12960 10854
rect 12984 10852 13040 10854
rect 13064 10852 13120 10854
rect 12824 9818 12880 9820
rect 12904 9818 12960 9820
rect 12984 9818 13040 9820
rect 13064 9818 13120 9820
rect 12824 9766 12870 9818
rect 12870 9766 12880 9818
rect 12904 9766 12934 9818
rect 12934 9766 12946 9818
rect 12946 9766 12960 9818
rect 12984 9766 12998 9818
rect 12998 9766 13010 9818
rect 13010 9766 13040 9818
rect 13064 9766 13074 9818
rect 13074 9766 13120 9818
rect 12824 9764 12880 9766
rect 12904 9764 12960 9766
rect 12984 9764 13040 9766
rect 13064 9764 13120 9766
rect 12824 8730 12880 8732
rect 12904 8730 12960 8732
rect 12984 8730 13040 8732
rect 13064 8730 13120 8732
rect 12824 8678 12870 8730
rect 12870 8678 12880 8730
rect 12904 8678 12934 8730
rect 12934 8678 12946 8730
rect 12946 8678 12960 8730
rect 12984 8678 12998 8730
rect 12998 8678 13010 8730
rect 13010 8678 13040 8730
rect 13064 8678 13074 8730
rect 13074 8678 13120 8730
rect 12824 8676 12880 8678
rect 12904 8676 12960 8678
rect 12984 8676 13040 8678
rect 13064 8676 13120 8678
rect 13542 19352 13598 19408
rect 13726 23296 13782 23352
rect 13634 18672 13690 18728
rect 15106 41112 15162 41168
rect 14738 28464 14794 28520
rect 14462 23432 14518 23488
rect 14186 20712 14242 20768
rect 12714 8336 12770 8392
rect 12824 7642 12880 7644
rect 12904 7642 12960 7644
rect 12984 7642 13040 7644
rect 13064 7642 13120 7644
rect 12824 7590 12870 7642
rect 12870 7590 12880 7642
rect 12904 7590 12934 7642
rect 12934 7590 12946 7642
rect 12946 7590 12960 7642
rect 12984 7590 12998 7642
rect 12998 7590 13010 7642
rect 13010 7590 13040 7642
rect 13064 7590 13074 7642
rect 13074 7590 13120 7642
rect 12824 7588 12880 7590
rect 12904 7588 12960 7590
rect 12984 7588 13040 7590
rect 13064 7588 13120 7590
rect 12806 6840 12862 6896
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 12254 3984 12310 4040
rect 12070 3576 12126 3632
rect 12162 3168 12218 3224
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 13818 12824 13874 12880
rect 13358 6024 13414 6080
rect 12622 5072 12678 5128
rect 13634 7520 13690 7576
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 13358 4120 13414 4176
rect 12622 3304 12678 3360
rect 11794 2352 11850 2408
rect 12070 1944 12126 2000
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 13726 3984 13782 4040
rect 12622 2080 12678 2136
rect 12898 2624 12954 2680
rect 13266 2388 13268 2408
rect 13268 2388 13320 2408
rect 13320 2388 13322 2408
rect 13266 2352 13322 2388
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 13542 1964 13598 2000
rect 13542 1944 13544 1964
rect 13544 1944 13596 1964
rect 13596 1944 13598 1964
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 14278 14592 14334 14648
rect 15791 43002 15847 43004
rect 15871 43002 15927 43004
rect 15951 43002 16007 43004
rect 16031 43002 16087 43004
rect 15791 42950 15837 43002
rect 15837 42950 15847 43002
rect 15871 42950 15901 43002
rect 15901 42950 15913 43002
rect 15913 42950 15927 43002
rect 15951 42950 15965 43002
rect 15965 42950 15977 43002
rect 15977 42950 16007 43002
rect 16031 42950 16041 43002
rect 16041 42950 16087 43002
rect 15791 42948 15847 42950
rect 15871 42948 15927 42950
rect 15951 42948 16007 42950
rect 16031 42948 16087 42950
rect 15658 42880 15714 42936
rect 15791 41914 15847 41916
rect 15871 41914 15927 41916
rect 15951 41914 16007 41916
rect 16031 41914 16087 41916
rect 15791 41862 15837 41914
rect 15837 41862 15847 41914
rect 15871 41862 15901 41914
rect 15901 41862 15913 41914
rect 15913 41862 15927 41914
rect 15951 41862 15965 41914
rect 15965 41862 15977 41914
rect 15977 41862 16007 41914
rect 16031 41862 16041 41914
rect 16041 41862 16087 41914
rect 15791 41860 15847 41862
rect 15871 41860 15927 41862
rect 15951 41860 16007 41862
rect 16031 41860 16087 41862
rect 15566 36624 15622 36680
rect 15474 33224 15530 33280
rect 15014 32544 15070 32600
rect 15198 31864 15254 31920
rect 15106 31048 15162 31104
rect 15014 27920 15070 27976
rect 15382 29280 15438 29336
rect 15566 29008 15622 29064
rect 15791 40826 15847 40828
rect 15871 40826 15927 40828
rect 15951 40826 16007 40828
rect 16031 40826 16087 40828
rect 15791 40774 15837 40826
rect 15837 40774 15847 40826
rect 15871 40774 15901 40826
rect 15901 40774 15913 40826
rect 15913 40774 15927 40826
rect 15951 40774 15965 40826
rect 15965 40774 15977 40826
rect 15977 40774 16007 40826
rect 16031 40774 16041 40826
rect 16041 40774 16087 40826
rect 15791 40772 15847 40774
rect 15871 40772 15927 40774
rect 15951 40772 16007 40774
rect 16031 40772 16087 40774
rect 15791 39738 15847 39740
rect 15871 39738 15927 39740
rect 15951 39738 16007 39740
rect 16031 39738 16087 39740
rect 15791 39686 15837 39738
rect 15837 39686 15847 39738
rect 15871 39686 15901 39738
rect 15901 39686 15913 39738
rect 15913 39686 15927 39738
rect 15951 39686 15965 39738
rect 15965 39686 15977 39738
rect 15977 39686 16007 39738
rect 16031 39686 16041 39738
rect 16041 39686 16087 39738
rect 15791 39684 15847 39686
rect 15871 39684 15927 39686
rect 15951 39684 16007 39686
rect 16031 39684 16087 39686
rect 15791 38650 15847 38652
rect 15871 38650 15927 38652
rect 15951 38650 16007 38652
rect 16031 38650 16087 38652
rect 15791 38598 15837 38650
rect 15837 38598 15847 38650
rect 15871 38598 15901 38650
rect 15901 38598 15913 38650
rect 15913 38598 15927 38650
rect 15951 38598 15965 38650
rect 15965 38598 15977 38650
rect 15977 38598 16007 38650
rect 16031 38598 16041 38650
rect 16041 38598 16087 38650
rect 15791 38596 15847 38598
rect 15871 38596 15927 38598
rect 15951 38596 16007 38598
rect 16031 38596 16087 38598
rect 15791 37562 15847 37564
rect 15871 37562 15927 37564
rect 15951 37562 16007 37564
rect 16031 37562 16087 37564
rect 15791 37510 15837 37562
rect 15837 37510 15847 37562
rect 15871 37510 15901 37562
rect 15901 37510 15913 37562
rect 15913 37510 15927 37562
rect 15951 37510 15965 37562
rect 15965 37510 15977 37562
rect 15977 37510 16007 37562
rect 16031 37510 16041 37562
rect 16041 37510 16087 37562
rect 15791 37508 15847 37510
rect 15871 37508 15927 37510
rect 15951 37508 16007 37510
rect 16031 37508 16087 37510
rect 15791 36474 15847 36476
rect 15871 36474 15927 36476
rect 15951 36474 16007 36476
rect 16031 36474 16087 36476
rect 15791 36422 15837 36474
rect 15837 36422 15847 36474
rect 15871 36422 15901 36474
rect 15901 36422 15913 36474
rect 15913 36422 15927 36474
rect 15951 36422 15965 36474
rect 15965 36422 15977 36474
rect 15977 36422 16007 36474
rect 16031 36422 16041 36474
rect 16041 36422 16087 36474
rect 15791 36420 15847 36422
rect 15871 36420 15927 36422
rect 15951 36420 16007 36422
rect 16031 36420 16087 36422
rect 15791 35386 15847 35388
rect 15871 35386 15927 35388
rect 15951 35386 16007 35388
rect 16031 35386 16087 35388
rect 15791 35334 15837 35386
rect 15837 35334 15847 35386
rect 15871 35334 15901 35386
rect 15901 35334 15913 35386
rect 15913 35334 15927 35386
rect 15951 35334 15965 35386
rect 15965 35334 15977 35386
rect 15977 35334 16007 35386
rect 16031 35334 16041 35386
rect 16041 35334 16087 35386
rect 15791 35332 15847 35334
rect 15871 35332 15927 35334
rect 15951 35332 16007 35334
rect 16031 35332 16087 35334
rect 15791 34298 15847 34300
rect 15871 34298 15927 34300
rect 15951 34298 16007 34300
rect 16031 34298 16087 34300
rect 15791 34246 15837 34298
rect 15837 34246 15847 34298
rect 15871 34246 15901 34298
rect 15901 34246 15913 34298
rect 15913 34246 15927 34298
rect 15951 34246 15965 34298
rect 15965 34246 15977 34298
rect 15977 34246 16007 34298
rect 16031 34246 16041 34298
rect 16041 34246 16087 34298
rect 15791 34244 15847 34246
rect 15871 34244 15927 34246
rect 15951 34244 16007 34246
rect 16031 34244 16087 34246
rect 15791 33210 15847 33212
rect 15871 33210 15927 33212
rect 15951 33210 16007 33212
rect 16031 33210 16087 33212
rect 15791 33158 15837 33210
rect 15837 33158 15847 33210
rect 15871 33158 15901 33210
rect 15901 33158 15913 33210
rect 15913 33158 15927 33210
rect 15951 33158 15965 33210
rect 15965 33158 15977 33210
rect 15977 33158 16007 33210
rect 16031 33158 16041 33210
rect 16041 33158 16087 33210
rect 15791 33156 15847 33158
rect 15871 33156 15927 33158
rect 15951 33156 16007 33158
rect 16031 33156 16087 33158
rect 16394 41656 16450 41712
rect 16026 32852 16028 32872
rect 16028 32852 16080 32872
rect 16080 32852 16082 32872
rect 16026 32816 16082 32852
rect 15791 32122 15847 32124
rect 15871 32122 15927 32124
rect 15951 32122 16007 32124
rect 16031 32122 16087 32124
rect 15791 32070 15837 32122
rect 15837 32070 15847 32122
rect 15871 32070 15901 32122
rect 15901 32070 15913 32122
rect 15913 32070 15927 32122
rect 15951 32070 15965 32122
rect 15965 32070 15977 32122
rect 15977 32070 16007 32122
rect 16031 32070 16041 32122
rect 16041 32070 16087 32122
rect 15791 32068 15847 32070
rect 15871 32068 15927 32070
rect 15951 32068 16007 32070
rect 16031 32068 16087 32070
rect 15791 31034 15847 31036
rect 15871 31034 15927 31036
rect 15951 31034 16007 31036
rect 16031 31034 16087 31036
rect 15791 30982 15837 31034
rect 15837 30982 15847 31034
rect 15871 30982 15901 31034
rect 15901 30982 15913 31034
rect 15913 30982 15927 31034
rect 15951 30982 15965 31034
rect 15965 30982 15977 31034
rect 15977 30982 16007 31034
rect 16031 30982 16041 31034
rect 16041 30982 16087 31034
rect 15791 30980 15847 30982
rect 15871 30980 15927 30982
rect 15951 30980 16007 30982
rect 16031 30980 16087 30982
rect 15791 29946 15847 29948
rect 15871 29946 15927 29948
rect 15951 29946 16007 29948
rect 16031 29946 16087 29948
rect 15791 29894 15837 29946
rect 15837 29894 15847 29946
rect 15871 29894 15901 29946
rect 15901 29894 15913 29946
rect 15913 29894 15927 29946
rect 15951 29894 15965 29946
rect 15965 29894 15977 29946
rect 15977 29894 16007 29946
rect 16031 29894 16041 29946
rect 16041 29894 16087 29946
rect 15791 29892 15847 29894
rect 15871 29892 15927 29894
rect 15951 29892 16007 29894
rect 16031 29892 16087 29894
rect 15750 29008 15806 29064
rect 15791 28858 15847 28860
rect 15871 28858 15927 28860
rect 15951 28858 16007 28860
rect 16031 28858 16087 28860
rect 15791 28806 15837 28858
rect 15837 28806 15847 28858
rect 15871 28806 15901 28858
rect 15901 28806 15913 28858
rect 15913 28806 15927 28858
rect 15951 28806 15965 28858
rect 15965 28806 15977 28858
rect 15977 28806 16007 28858
rect 16031 28806 16041 28858
rect 16041 28806 16087 28858
rect 15791 28804 15847 28806
rect 15871 28804 15927 28806
rect 15951 28804 16007 28806
rect 16031 28804 16087 28806
rect 16210 29280 16266 29336
rect 15791 27770 15847 27772
rect 15871 27770 15927 27772
rect 15951 27770 16007 27772
rect 16031 27770 16087 27772
rect 15791 27718 15837 27770
rect 15837 27718 15847 27770
rect 15871 27718 15901 27770
rect 15901 27718 15913 27770
rect 15913 27718 15927 27770
rect 15951 27718 15965 27770
rect 15965 27718 15977 27770
rect 15977 27718 16007 27770
rect 16031 27718 16041 27770
rect 16041 27718 16087 27770
rect 15791 27716 15847 27718
rect 15871 27716 15927 27718
rect 15951 27716 16007 27718
rect 16031 27716 16087 27718
rect 14738 20712 14794 20768
rect 14462 17040 14518 17096
rect 14738 11736 14794 11792
rect 15382 21140 15438 21176
rect 15382 21120 15384 21140
rect 15384 21120 15436 21140
rect 15436 21120 15438 21140
rect 14922 13932 14978 13968
rect 14922 13912 14924 13932
rect 14924 13912 14976 13932
rect 14976 13912 14978 13932
rect 15791 26682 15847 26684
rect 15871 26682 15927 26684
rect 15951 26682 16007 26684
rect 16031 26682 16087 26684
rect 15791 26630 15837 26682
rect 15837 26630 15847 26682
rect 15871 26630 15901 26682
rect 15901 26630 15913 26682
rect 15913 26630 15927 26682
rect 15951 26630 15965 26682
rect 15965 26630 15977 26682
rect 15977 26630 16007 26682
rect 16031 26630 16041 26682
rect 16041 26630 16087 26682
rect 15791 26628 15847 26630
rect 15871 26628 15927 26630
rect 15951 26628 16007 26630
rect 16031 26628 16087 26630
rect 15791 25594 15847 25596
rect 15871 25594 15927 25596
rect 15951 25594 16007 25596
rect 16031 25594 16087 25596
rect 15791 25542 15837 25594
rect 15837 25542 15847 25594
rect 15871 25542 15901 25594
rect 15901 25542 15913 25594
rect 15913 25542 15927 25594
rect 15951 25542 15965 25594
rect 15965 25542 15977 25594
rect 15977 25542 16007 25594
rect 16031 25542 16041 25594
rect 16041 25542 16087 25594
rect 15791 25540 15847 25542
rect 15871 25540 15927 25542
rect 15951 25540 16007 25542
rect 16031 25540 16087 25542
rect 15791 24506 15847 24508
rect 15871 24506 15927 24508
rect 15951 24506 16007 24508
rect 16031 24506 16087 24508
rect 15791 24454 15837 24506
rect 15837 24454 15847 24506
rect 15871 24454 15901 24506
rect 15901 24454 15913 24506
rect 15913 24454 15927 24506
rect 15951 24454 15965 24506
rect 15965 24454 15977 24506
rect 15977 24454 16007 24506
rect 16031 24454 16041 24506
rect 16041 24454 16087 24506
rect 15791 24452 15847 24454
rect 15871 24452 15927 24454
rect 15951 24452 16007 24454
rect 16031 24452 16087 24454
rect 16302 25200 16358 25256
rect 15791 23418 15847 23420
rect 15871 23418 15927 23420
rect 15951 23418 16007 23420
rect 16031 23418 16087 23420
rect 15791 23366 15837 23418
rect 15837 23366 15847 23418
rect 15871 23366 15901 23418
rect 15901 23366 15913 23418
rect 15913 23366 15927 23418
rect 15951 23366 15965 23418
rect 15965 23366 15977 23418
rect 15977 23366 16007 23418
rect 16031 23366 16041 23418
rect 16041 23366 16087 23418
rect 15791 23364 15847 23366
rect 15871 23364 15927 23366
rect 15951 23364 16007 23366
rect 16031 23364 16087 23366
rect 16118 22480 16174 22536
rect 15791 22330 15847 22332
rect 15871 22330 15927 22332
rect 15951 22330 16007 22332
rect 16031 22330 16087 22332
rect 15791 22278 15837 22330
rect 15837 22278 15847 22330
rect 15871 22278 15901 22330
rect 15901 22278 15913 22330
rect 15913 22278 15927 22330
rect 15951 22278 15965 22330
rect 15965 22278 15977 22330
rect 15977 22278 16007 22330
rect 16031 22278 16041 22330
rect 16041 22278 16087 22330
rect 15791 22276 15847 22278
rect 15871 22276 15927 22278
rect 15951 22276 16007 22278
rect 16031 22276 16087 22278
rect 15791 21242 15847 21244
rect 15871 21242 15927 21244
rect 15951 21242 16007 21244
rect 16031 21242 16087 21244
rect 15791 21190 15837 21242
rect 15837 21190 15847 21242
rect 15871 21190 15901 21242
rect 15901 21190 15913 21242
rect 15913 21190 15927 21242
rect 15951 21190 15965 21242
rect 15965 21190 15977 21242
rect 15977 21190 16007 21242
rect 16031 21190 16041 21242
rect 16041 21190 16087 21242
rect 15791 21188 15847 21190
rect 15871 21188 15927 21190
rect 15951 21188 16007 21190
rect 16031 21188 16087 21190
rect 15791 20154 15847 20156
rect 15871 20154 15927 20156
rect 15951 20154 16007 20156
rect 16031 20154 16087 20156
rect 15791 20102 15837 20154
rect 15837 20102 15847 20154
rect 15871 20102 15901 20154
rect 15901 20102 15913 20154
rect 15913 20102 15927 20154
rect 15951 20102 15965 20154
rect 15965 20102 15977 20154
rect 15977 20102 16007 20154
rect 16031 20102 16041 20154
rect 16041 20102 16087 20154
rect 15791 20100 15847 20102
rect 15871 20100 15927 20102
rect 15951 20100 16007 20102
rect 16031 20100 16087 20102
rect 15791 19066 15847 19068
rect 15871 19066 15927 19068
rect 15951 19066 16007 19068
rect 16031 19066 16087 19068
rect 15791 19014 15837 19066
rect 15837 19014 15847 19066
rect 15871 19014 15901 19066
rect 15901 19014 15913 19066
rect 15913 19014 15927 19066
rect 15951 19014 15965 19066
rect 15965 19014 15977 19066
rect 15977 19014 16007 19066
rect 16031 19014 16041 19066
rect 16041 19014 16087 19066
rect 15791 19012 15847 19014
rect 15871 19012 15927 19014
rect 15951 19012 16007 19014
rect 16031 19012 16087 19014
rect 16854 38936 16910 38992
rect 17314 41792 17370 41848
rect 17590 41656 17646 41712
rect 17774 41540 17830 41576
rect 17774 41520 17776 41540
rect 17776 41520 17828 41540
rect 17828 41520 17830 41540
rect 18758 43546 18814 43548
rect 18838 43546 18894 43548
rect 18918 43546 18974 43548
rect 18998 43546 19054 43548
rect 18758 43494 18804 43546
rect 18804 43494 18814 43546
rect 18838 43494 18868 43546
rect 18868 43494 18880 43546
rect 18880 43494 18894 43546
rect 18918 43494 18932 43546
rect 18932 43494 18944 43546
rect 18944 43494 18974 43546
rect 18998 43494 19008 43546
rect 19008 43494 19054 43546
rect 18758 43492 18814 43494
rect 18838 43492 18894 43494
rect 18918 43492 18974 43494
rect 18998 43492 19054 43494
rect 18758 42458 18814 42460
rect 18838 42458 18894 42460
rect 18918 42458 18974 42460
rect 18998 42458 19054 42460
rect 18758 42406 18804 42458
rect 18804 42406 18814 42458
rect 18838 42406 18868 42458
rect 18868 42406 18880 42458
rect 18880 42406 18894 42458
rect 18918 42406 18932 42458
rect 18932 42406 18944 42458
rect 18944 42406 18974 42458
rect 18998 42406 19008 42458
rect 19008 42406 19054 42458
rect 18758 42404 18814 42406
rect 18838 42404 18894 42406
rect 18918 42404 18974 42406
rect 18998 42404 19054 42406
rect 18418 41656 18474 41712
rect 18050 41384 18106 41440
rect 18510 38664 18566 38720
rect 18758 41370 18814 41372
rect 18838 41370 18894 41372
rect 18918 41370 18974 41372
rect 18998 41370 19054 41372
rect 18758 41318 18804 41370
rect 18804 41318 18814 41370
rect 18838 41318 18868 41370
rect 18868 41318 18880 41370
rect 18880 41318 18894 41370
rect 18918 41318 18932 41370
rect 18932 41318 18944 41370
rect 18944 41318 18974 41370
rect 18998 41318 19008 41370
rect 19008 41318 19054 41370
rect 18758 41316 18814 41318
rect 18838 41316 18894 41318
rect 18918 41316 18974 41318
rect 18998 41316 19054 41318
rect 18758 40282 18814 40284
rect 18838 40282 18894 40284
rect 18918 40282 18974 40284
rect 18998 40282 19054 40284
rect 18758 40230 18804 40282
rect 18804 40230 18814 40282
rect 18838 40230 18868 40282
rect 18868 40230 18880 40282
rect 18880 40230 18894 40282
rect 18918 40230 18932 40282
rect 18932 40230 18944 40282
rect 18944 40230 18974 40282
rect 18998 40230 19008 40282
rect 19008 40230 19054 40282
rect 18758 40228 18814 40230
rect 18838 40228 18894 40230
rect 18918 40228 18974 40230
rect 18998 40228 19054 40230
rect 18758 39194 18814 39196
rect 18838 39194 18894 39196
rect 18918 39194 18974 39196
rect 18998 39194 19054 39196
rect 18758 39142 18804 39194
rect 18804 39142 18814 39194
rect 18838 39142 18868 39194
rect 18868 39142 18880 39194
rect 18880 39142 18894 39194
rect 18918 39142 18932 39194
rect 18932 39142 18944 39194
rect 18944 39142 18974 39194
rect 18998 39142 19008 39194
rect 19008 39142 19054 39194
rect 18758 39140 18814 39142
rect 18838 39140 18894 39142
rect 18918 39140 18974 39142
rect 18998 39140 19054 39142
rect 19430 41656 19486 41712
rect 18758 38106 18814 38108
rect 18838 38106 18894 38108
rect 18918 38106 18974 38108
rect 18998 38106 19054 38108
rect 18758 38054 18804 38106
rect 18804 38054 18814 38106
rect 18838 38054 18868 38106
rect 18868 38054 18880 38106
rect 18880 38054 18894 38106
rect 18918 38054 18932 38106
rect 18932 38054 18944 38106
rect 18944 38054 18974 38106
rect 18998 38054 19008 38106
rect 19008 38054 19054 38106
rect 18758 38052 18814 38054
rect 18838 38052 18894 38054
rect 18918 38052 18974 38054
rect 18998 38052 19054 38054
rect 16854 31340 16910 31376
rect 16854 31320 16856 31340
rect 16856 31320 16908 31340
rect 16908 31320 16910 31340
rect 16946 29164 17002 29200
rect 16946 29144 16948 29164
rect 16948 29144 17000 29164
rect 17000 29144 17002 29164
rect 17038 28736 17094 28792
rect 17038 28600 17094 28656
rect 17130 27784 17186 27840
rect 16762 24792 16818 24848
rect 16578 23740 16580 23760
rect 16580 23740 16632 23760
rect 16632 23740 16634 23760
rect 16578 23704 16634 23740
rect 18142 32272 18198 32328
rect 17866 28328 17922 28384
rect 16578 21528 16634 21584
rect 16762 21664 16818 21720
rect 16946 21664 17002 21720
rect 17498 24812 17554 24848
rect 17498 24792 17500 24812
rect 17500 24792 17552 24812
rect 17552 24792 17554 24812
rect 17222 21528 17278 21584
rect 15474 16496 15530 16552
rect 15198 15544 15254 15600
rect 14922 11076 14978 11112
rect 14922 11056 14924 11076
rect 14924 11056 14976 11076
rect 14976 11056 14978 11076
rect 15106 10920 15162 10976
rect 15474 10784 15530 10840
rect 15791 17978 15847 17980
rect 15871 17978 15927 17980
rect 15951 17978 16007 17980
rect 16031 17978 16087 17980
rect 15791 17926 15837 17978
rect 15837 17926 15847 17978
rect 15871 17926 15901 17978
rect 15901 17926 15913 17978
rect 15913 17926 15927 17978
rect 15951 17926 15965 17978
rect 15965 17926 15977 17978
rect 15977 17926 16007 17978
rect 16031 17926 16041 17978
rect 16041 17926 16087 17978
rect 15791 17924 15847 17926
rect 15871 17924 15927 17926
rect 15951 17924 16007 17926
rect 16031 17924 16087 17926
rect 15791 16890 15847 16892
rect 15871 16890 15927 16892
rect 15951 16890 16007 16892
rect 16031 16890 16087 16892
rect 15791 16838 15837 16890
rect 15837 16838 15847 16890
rect 15871 16838 15901 16890
rect 15901 16838 15913 16890
rect 15913 16838 15927 16890
rect 15951 16838 15965 16890
rect 15965 16838 15977 16890
rect 15977 16838 16007 16890
rect 16031 16838 16041 16890
rect 16041 16838 16087 16890
rect 15791 16836 15847 16838
rect 15871 16836 15927 16838
rect 15951 16836 16007 16838
rect 16031 16836 16087 16838
rect 15842 15952 15898 16008
rect 15791 15802 15847 15804
rect 15871 15802 15927 15804
rect 15951 15802 16007 15804
rect 16031 15802 16087 15804
rect 15791 15750 15837 15802
rect 15837 15750 15847 15802
rect 15871 15750 15901 15802
rect 15901 15750 15913 15802
rect 15913 15750 15927 15802
rect 15951 15750 15965 15802
rect 15965 15750 15977 15802
rect 15977 15750 16007 15802
rect 16031 15750 16041 15802
rect 16041 15750 16087 15802
rect 15791 15748 15847 15750
rect 15871 15748 15927 15750
rect 15951 15748 16007 15750
rect 16031 15748 16087 15750
rect 16210 15136 16266 15192
rect 15791 14714 15847 14716
rect 15871 14714 15927 14716
rect 15951 14714 16007 14716
rect 16031 14714 16087 14716
rect 15791 14662 15837 14714
rect 15837 14662 15847 14714
rect 15871 14662 15901 14714
rect 15901 14662 15913 14714
rect 15913 14662 15927 14714
rect 15951 14662 15965 14714
rect 15965 14662 15977 14714
rect 15977 14662 16007 14714
rect 16031 14662 16041 14714
rect 16041 14662 16087 14714
rect 15791 14660 15847 14662
rect 15871 14660 15927 14662
rect 15951 14660 16007 14662
rect 16031 14660 16087 14662
rect 16118 14340 16174 14376
rect 16118 14320 16120 14340
rect 16120 14320 16172 14340
rect 16172 14320 16174 14340
rect 15791 13626 15847 13628
rect 15871 13626 15927 13628
rect 15951 13626 16007 13628
rect 16031 13626 16087 13628
rect 15791 13574 15837 13626
rect 15837 13574 15847 13626
rect 15871 13574 15901 13626
rect 15901 13574 15913 13626
rect 15913 13574 15927 13626
rect 15951 13574 15965 13626
rect 15965 13574 15977 13626
rect 15977 13574 16007 13626
rect 16031 13574 16041 13626
rect 16041 13574 16087 13626
rect 15791 13572 15847 13574
rect 15871 13572 15927 13574
rect 15951 13572 16007 13574
rect 16031 13572 16087 13574
rect 15791 12538 15847 12540
rect 15871 12538 15927 12540
rect 15951 12538 16007 12540
rect 16031 12538 16087 12540
rect 15791 12486 15837 12538
rect 15837 12486 15847 12538
rect 15871 12486 15901 12538
rect 15901 12486 15913 12538
rect 15913 12486 15927 12538
rect 15951 12486 15965 12538
rect 15965 12486 15977 12538
rect 15977 12486 16007 12538
rect 16031 12486 16041 12538
rect 16041 12486 16087 12538
rect 15791 12484 15847 12486
rect 15871 12484 15927 12486
rect 15951 12484 16007 12486
rect 16031 12484 16087 12486
rect 15791 11450 15847 11452
rect 15871 11450 15927 11452
rect 15951 11450 16007 11452
rect 16031 11450 16087 11452
rect 15791 11398 15837 11450
rect 15837 11398 15847 11450
rect 15871 11398 15901 11450
rect 15901 11398 15913 11450
rect 15913 11398 15927 11450
rect 15951 11398 15965 11450
rect 15965 11398 15977 11450
rect 15977 11398 16007 11450
rect 16031 11398 16041 11450
rect 16041 11398 16087 11450
rect 15791 11396 15847 11398
rect 15871 11396 15927 11398
rect 15951 11396 16007 11398
rect 16031 11396 16087 11398
rect 16854 17856 16910 17912
rect 17130 18944 17186 19000
rect 17038 18808 17094 18864
rect 16946 13776 17002 13832
rect 15791 10362 15847 10364
rect 15871 10362 15927 10364
rect 15951 10362 16007 10364
rect 16031 10362 16087 10364
rect 15791 10310 15837 10362
rect 15837 10310 15847 10362
rect 15871 10310 15901 10362
rect 15901 10310 15913 10362
rect 15913 10310 15927 10362
rect 15951 10310 15965 10362
rect 15965 10310 15977 10362
rect 15977 10310 16007 10362
rect 16031 10310 16041 10362
rect 16041 10310 16087 10362
rect 15791 10308 15847 10310
rect 15871 10308 15927 10310
rect 15951 10308 16007 10310
rect 16031 10308 16087 10310
rect 16578 11600 16634 11656
rect 16486 10648 16542 10704
rect 16210 9696 16266 9752
rect 15791 9274 15847 9276
rect 15871 9274 15927 9276
rect 15951 9274 16007 9276
rect 16031 9274 16087 9276
rect 15791 9222 15837 9274
rect 15837 9222 15847 9274
rect 15871 9222 15901 9274
rect 15901 9222 15913 9274
rect 15913 9222 15927 9274
rect 15951 9222 15965 9274
rect 15965 9222 15977 9274
rect 15977 9222 16007 9274
rect 16031 9222 16041 9274
rect 16041 9222 16087 9274
rect 15791 9220 15847 9222
rect 15871 9220 15927 9222
rect 15951 9220 16007 9222
rect 16031 9220 16087 9222
rect 15791 8186 15847 8188
rect 15871 8186 15927 8188
rect 15951 8186 16007 8188
rect 16031 8186 16087 8188
rect 15791 8134 15837 8186
rect 15837 8134 15847 8186
rect 15871 8134 15901 8186
rect 15901 8134 15913 8186
rect 15913 8134 15927 8186
rect 15951 8134 15965 8186
rect 15965 8134 15977 8186
rect 15977 8134 16007 8186
rect 16031 8134 16041 8186
rect 16041 8134 16087 8186
rect 15791 8132 15847 8134
rect 15871 8132 15927 8134
rect 15951 8132 16007 8134
rect 16031 8132 16087 8134
rect 15791 7098 15847 7100
rect 15871 7098 15927 7100
rect 15951 7098 16007 7100
rect 16031 7098 16087 7100
rect 15791 7046 15837 7098
rect 15837 7046 15847 7098
rect 15871 7046 15901 7098
rect 15901 7046 15913 7098
rect 15913 7046 15927 7098
rect 15951 7046 15965 7098
rect 15965 7046 15977 7098
rect 15977 7046 16007 7098
rect 16031 7046 16041 7098
rect 16041 7046 16087 7098
rect 15791 7044 15847 7046
rect 15871 7044 15927 7046
rect 15951 7044 16007 7046
rect 16031 7044 16087 7046
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 15566 4936 15622 4992
rect 15566 4564 15568 4584
rect 15568 4564 15620 4584
rect 15620 4564 15622 4584
rect 15566 4528 15622 4564
rect 15566 2488 15622 2544
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 16210 7928 16266 7984
rect 16210 5072 16266 5128
rect 17498 21664 17554 21720
rect 17866 20440 17922 20496
rect 17866 17040 17922 17096
rect 18234 30096 18290 30152
rect 18234 25744 18290 25800
rect 18418 30368 18474 30424
rect 18758 37018 18814 37020
rect 18838 37018 18894 37020
rect 18918 37018 18974 37020
rect 18998 37018 19054 37020
rect 18758 36966 18804 37018
rect 18804 36966 18814 37018
rect 18838 36966 18868 37018
rect 18868 36966 18880 37018
rect 18880 36966 18894 37018
rect 18918 36966 18932 37018
rect 18932 36966 18944 37018
rect 18944 36966 18974 37018
rect 18998 36966 19008 37018
rect 19008 36966 19054 37018
rect 18758 36964 18814 36966
rect 18838 36964 18894 36966
rect 18918 36964 18974 36966
rect 18998 36964 19054 36966
rect 19706 40160 19762 40216
rect 18758 35930 18814 35932
rect 18838 35930 18894 35932
rect 18918 35930 18974 35932
rect 18998 35930 19054 35932
rect 18758 35878 18804 35930
rect 18804 35878 18814 35930
rect 18838 35878 18868 35930
rect 18868 35878 18880 35930
rect 18880 35878 18894 35930
rect 18918 35878 18932 35930
rect 18932 35878 18944 35930
rect 18944 35878 18974 35930
rect 18998 35878 19008 35930
rect 19008 35878 19054 35930
rect 18758 35876 18814 35878
rect 18838 35876 18894 35878
rect 18918 35876 18974 35878
rect 18998 35876 19054 35878
rect 18878 35556 18934 35592
rect 18878 35536 18880 35556
rect 18880 35536 18932 35556
rect 18932 35536 18934 35556
rect 18758 34842 18814 34844
rect 18838 34842 18894 34844
rect 18918 34842 18974 34844
rect 18998 34842 19054 34844
rect 18758 34790 18804 34842
rect 18804 34790 18814 34842
rect 18838 34790 18868 34842
rect 18868 34790 18880 34842
rect 18880 34790 18894 34842
rect 18918 34790 18932 34842
rect 18932 34790 18944 34842
rect 18944 34790 18974 34842
rect 18998 34790 19008 34842
rect 19008 34790 19054 34842
rect 18758 34788 18814 34790
rect 18838 34788 18894 34790
rect 18918 34788 18974 34790
rect 18998 34788 19054 34790
rect 18758 33754 18814 33756
rect 18838 33754 18894 33756
rect 18918 33754 18974 33756
rect 18998 33754 19054 33756
rect 18758 33702 18804 33754
rect 18804 33702 18814 33754
rect 18838 33702 18868 33754
rect 18868 33702 18880 33754
rect 18880 33702 18894 33754
rect 18918 33702 18932 33754
rect 18932 33702 18944 33754
rect 18944 33702 18974 33754
rect 18998 33702 19008 33754
rect 19008 33702 19054 33754
rect 18758 33700 18814 33702
rect 18838 33700 18894 33702
rect 18918 33700 18974 33702
rect 18998 33700 19054 33702
rect 18878 33496 18934 33552
rect 18758 32666 18814 32668
rect 18838 32666 18894 32668
rect 18918 32666 18974 32668
rect 18998 32666 19054 32668
rect 18758 32614 18804 32666
rect 18804 32614 18814 32666
rect 18838 32614 18868 32666
rect 18868 32614 18880 32666
rect 18880 32614 18894 32666
rect 18918 32614 18932 32666
rect 18932 32614 18944 32666
rect 18944 32614 18974 32666
rect 18998 32614 19008 32666
rect 19008 32614 19054 32666
rect 18758 32612 18814 32614
rect 18838 32612 18894 32614
rect 18918 32612 18974 32614
rect 18998 32612 19054 32614
rect 18758 31578 18814 31580
rect 18838 31578 18894 31580
rect 18918 31578 18974 31580
rect 18998 31578 19054 31580
rect 18758 31526 18804 31578
rect 18804 31526 18814 31578
rect 18838 31526 18868 31578
rect 18868 31526 18880 31578
rect 18880 31526 18894 31578
rect 18918 31526 18932 31578
rect 18932 31526 18944 31578
rect 18944 31526 18974 31578
rect 18998 31526 19008 31578
rect 19008 31526 19054 31578
rect 18758 31524 18814 31526
rect 18838 31524 18894 31526
rect 18918 31524 18974 31526
rect 18998 31524 19054 31526
rect 18758 30490 18814 30492
rect 18838 30490 18894 30492
rect 18918 30490 18974 30492
rect 18998 30490 19054 30492
rect 18758 30438 18804 30490
rect 18804 30438 18814 30490
rect 18838 30438 18868 30490
rect 18868 30438 18880 30490
rect 18880 30438 18894 30490
rect 18918 30438 18932 30490
rect 18932 30438 18944 30490
rect 18944 30438 18974 30490
rect 18998 30438 19008 30490
rect 19008 30438 19054 30490
rect 18758 30436 18814 30438
rect 18838 30436 18894 30438
rect 18918 30436 18974 30438
rect 18998 30436 19054 30438
rect 18758 29402 18814 29404
rect 18838 29402 18894 29404
rect 18918 29402 18974 29404
rect 18998 29402 19054 29404
rect 18758 29350 18804 29402
rect 18804 29350 18814 29402
rect 18838 29350 18868 29402
rect 18868 29350 18880 29402
rect 18880 29350 18894 29402
rect 18918 29350 18932 29402
rect 18932 29350 18944 29402
rect 18944 29350 18974 29402
rect 18998 29350 19008 29402
rect 19008 29350 19054 29402
rect 18758 29348 18814 29350
rect 18838 29348 18894 29350
rect 18918 29348 18974 29350
rect 18998 29348 19054 29350
rect 19522 32444 19524 32464
rect 19524 32444 19576 32464
rect 19576 32444 19578 32464
rect 19522 32408 19578 32444
rect 18758 28314 18814 28316
rect 18838 28314 18894 28316
rect 18918 28314 18974 28316
rect 18998 28314 19054 28316
rect 18758 28262 18804 28314
rect 18804 28262 18814 28314
rect 18838 28262 18868 28314
rect 18868 28262 18880 28314
rect 18880 28262 18894 28314
rect 18918 28262 18932 28314
rect 18932 28262 18944 28314
rect 18944 28262 18974 28314
rect 18998 28262 19008 28314
rect 19008 28262 19054 28314
rect 18758 28260 18814 28262
rect 18838 28260 18894 28262
rect 18918 28260 18974 28262
rect 18998 28260 19054 28262
rect 19430 28736 19486 28792
rect 19430 28092 19432 28112
rect 19432 28092 19484 28112
rect 19484 28092 19486 28112
rect 18758 27226 18814 27228
rect 18838 27226 18894 27228
rect 18918 27226 18974 27228
rect 18998 27226 19054 27228
rect 18758 27174 18804 27226
rect 18804 27174 18814 27226
rect 18838 27174 18868 27226
rect 18868 27174 18880 27226
rect 18880 27174 18894 27226
rect 18918 27174 18932 27226
rect 18932 27174 18944 27226
rect 18944 27174 18974 27226
rect 18998 27174 19008 27226
rect 19008 27174 19054 27226
rect 18758 27172 18814 27174
rect 18838 27172 18894 27174
rect 18918 27172 18974 27174
rect 18998 27172 19054 27174
rect 18758 26138 18814 26140
rect 18838 26138 18894 26140
rect 18918 26138 18974 26140
rect 18998 26138 19054 26140
rect 18758 26086 18804 26138
rect 18804 26086 18814 26138
rect 18838 26086 18868 26138
rect 18868 26086 18880 26138
rect 18880 26086 18894 26138
rect 18918 26086 18932 26138
rect 18932 26086 18944 26138
rect 18944 26086 18974 26138
rect 18998 26086 19008 26138
rect 19008 26086 19054 26138
rect 18758 26084 18814 26086
rect 18838 26084 18894 26086
rect 18918 26084 18974 26086
rect 18998 26084 19054 26086
rect 19430 28056 19486 28092
rect 18758 25050 18814 25052
rect 18838 25050 18894 25052
rect 18918 25050 18974 25052
rect 18998 25050 19054 25052
rect 18758 24998 18804 25050
rect 18804 24998 18814 25050
rect 18838 24998 18868 25050
rect 18868 24998 18880 25050
rect 18880 24998 18894 25050
rect 18918 24998 18932 25050
rect 18932 24998 18944 25050
rect 18944 24998 18974 25050
rect 18998 24998 19008 25050
rect 19008 24998 19054 25050
rect 18758 24996 18814 24998
rect 18838 24996 18894 24998
rect 18918 24996 18974 24998
rect 18998 24996 19054 24998
rect 17498 15000 17554 15056
rect 17222 11328 17278 11384
rect 17038 11076 17094 11112
rect 17038 11056 17040 11076
rect 17040 11056 17092 11076
rect 17092 11056 17094 11076
rect 16394 5616 16450 5672
rect 16578 4664 16634 4720
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 16394 2388 16396 2408
rect 16396 2388 16448 2408
rect 16448 2388 16450 2408
rect 16394 2352 16450 2388
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 17774 14476 17830 14512
rect 17774 14456 17776 14476
rect 17776 14456 17828 14476
rect 17828 14456 17830 14476
rect 17958 11192 18014 11248
rect 17774 9424 17830 9480
rect 17498 5752 17554 5808
rect 17590 4664 17646 4720
rect 18142 8336 18198 8392
rect 17958 6704 18014 6760
rect 18142 6704 18198 6760
rect 18758 23962 18814 23964
rect 18838 23962 18894 23964
rect 18918 23962 18974 23964
rect 18998 23962 19054 23964
rect 18758 23910 18804 23962
rect 18804 23910 18814 23962
rect 18838 23910 18868 23962
rect 18868 23910 18880 23962
rect 18880 23910 18894 23962
rect 18918 23910 18932 23962
rect 18932 23910 18944 23962
rect 18944 23910 18974 23962
rect 18998 23910 19008 23962
rect 19008 23910 19054 23962
rect 18758 23908 18814 23910
rect 18838 23908 18894 23910
rect 18918 23908 18974 23910
rect 18998 23908 19054 23910
rect 20074 42064 20130 42120
rect 20718 42064 20774 42120
rect 20350 41692 20352 41712
rect 20352 41692 20404 41712
rect 20404 41692 20406 41712
rect 20350 41656 20406 41692
rect 20074 40024 20130 40080
rect 19982 39344 20038 39400
rect 20258 40296 20314 40352
rect 20442 38836 20444 38856
rect 20444 38836 20496 38856
rect 20496 38836 20498 38856
rect 20442 38800 20498 38836
rect 20626 40432 20682 40488
rect 20810 40160 20866 40216
rect 21362 41656 21418 41712
rect 20810 39480 20866 39536
rect 19706 24792 19762 24848
rect 18758 22874 18814 22876
rect 18838 22874 18894 22876
rect 18918 22874 18974 22876
rect 18998 22874 19054 22876
rect 18758 22822 18804 22874
rect 18804 22822 18814 22874
rect 18838 22822 18868 22874
rect 18868 22822 18880 22874
rect 18880 22822 18894 22874
rect 18918 22822 18932 22874
rect 18932 22822 18944 22874
rect 18944 22822 18974 22874
rect 18998 22822 19008 22874
rect 19008 22822 19054 22874
rect 18758 22820 18814 22822
rect 18838 22820 18894 22822
rect 18918 22820 18974 22822
rect 18998 22820 19054 22822
rect 18758 21786 18814 21788
rect 18838 21786 18894 21788
rect 18918 21786 18974 21788
rect 18998 21786 19054 21788
rect 18758 21734 18804 21786
rect 18804 21734 18814 21786
rect 18838 21734 18868 21786
rect 18868 21734 18880 21786
rect 18880 21734 18894 21786
rect 18918 21734 18932 21786
rect 18932 21734 18944 21786
rect 18944 21734 18974 21786
rect 18998 21734 19008 21786
rect 19008 21734 19054 21786
rect 18758 21732 18814 21734
rect 18838 21732 18894 21734
rect 18918 21732 18974 21734
rect 18998 21732 19054 21734
rect 18758 20698 18814 20700
rect 18838 20698 18894 20700
rect 18918 20698 18974 20700
rect 18998 20698 19054 20700
rect 18758 20646 18804 20698
rect 18804 20646 18814 20698
rect 18838 20646 18868 20698
rect 18868 20646 18880 20698
rect 18880 20646 18894 20698
rect 18918 20646 18932 20698
rect 18932 20646 18944 20698
rect 18944 20646 18974 20698
rect 18998 20646 19008 20698
rect 19008 20646 19054 20698
rect 18758 20644 18814 20646
rect 18838 20644 18894 20646
rect 18918 20644 18974 20646
rect 18998 20644 19054 20646
rect 18758 19610 18814 19612
rect 18838 19610 18894 19612
rect 18918 19610 18974 19612
rect 18998 19610 19054 19612
rect 18758 19558 18804 19610
rect 18804 19558 18814 19610
rect 18838 19558 18868 19610
rect 18868 19558 18880 19610
rect 18880 19558 18894 19610
rect 18918 19558 18932 19610
rect 18932 19558 18944 19610
rect 18944 19558 18974 19610
rect 18998 19558 19008 19610
rect 19008 19558 19054 19610
rect 18758 19556 18814 19558
rect 18838 19556 18894 19558
rect 18918 19556 18974 19558
rect 18998 19556 19054 19558
rect 18758 18522 18814 18524
rect 18838 18522 18894 18524
rect 18918 18522 18974 18524
rect 18998 18522 19054 18524
rect 18758 18470 18804 18522
rect 18804 18470 18814 18522
rect 18838 18470 18868 18522
rect 18868 18470 18880 18522
rect 18880 18470 18894 18522
rect 18918 18470 18932 18522
rect 18932 18470 18944 18522
rect 18944 18470 18974 18522
rect 18998 18470 19008 18522
rect 19008 18470 19054 18522
rect 18758 18468 18814 18470
rect 18838 18468 18894 18470
rect 18918 18468 18974 18470
rect 18998 18468 19054 18470
rect 18758 17434 18814 17436
rect 18838 17434 18894 17436
rect 18918 17434 18974 17436
rect 18998 17434 19054 17436
rect 18758 17382 18804 17434
rect 18804 17382 18814 17434
rect 18838 17382 18868 17434
rect 18868 17382 18880 17434
rect 18880 17382 18894 17434
rect 18918 17382 18932 17434
rect 18932 17382 18944 17434
rect 18944 17382 18974 17434
rect 18998 17382 19008 17434
rect 19008 17382 19054 17434
rect 18758 17380 18814 17382
rect 18838 17380 18894 17382
rect 18918 17380 18974 17382
rect 18998 17380 19054 17382
rect 20258 28736 20314 28792
rect 20074 25236 20076 25256
rect 20076 25236 20128 25256
rect 20128 25236 20130 25256
rect 20074 25200 20130 25236
rect 18758 16346 18814 16348
rect 18838 16346 18894 16348
rect 18918 16346 18974 16348
rect 18998 16346 19054 16348
rect 18758 16294 18804 16346
rect 18804 16294 18814 16346
rect 18838 16294 18868 16346
rect 18868 16294 18880 16346
rect 18880 16294 18894 16346
rect 18918 16294 18932 16346
rect 18932 16294 18944 16346
rect 18944 16294 18974 16346
rect 18998 16294 19008 16346
rect 19008 16294 19054 16346
rect 18758 16292 18814 16294
rect 18838 16292 18894 16294
rect 18918 16292 18974 16294
rect 18998 16292 19054 16294
rect 18758 15258 18814 15260
rect 18838 15258 18894 15260
rect 18918 15258 18974 15260
rect 18998 15258 19054 15260
rect 18758 15206 18804 15258
rect 18804 15206 18814 15258
rect 18838 15206 18868 15258
rect 18868 15206 18880 15258
rect 18880 15206 18894 15258
rect 18918 15206 18932 15258
rect 18932 15206 18944 15258
rect 18944 15206 18974 15258
rect 18998 15206 19008 15258
rect 19008 15206 19054 15258
rect 18758 15204 18814 15206
rect 18838 15204 18894 15206
rect 18918 15204 18974 15206
rect 18998 15204 19054 15206
rect 18758 14170 18814 14172
rect 18838 14170 18894 14172
rect 18918 14170 18974 14172
rect 18998 14170 19054 14172
rect 18758 14118 18804 14170
rect 18804 14118 18814 14170
rect 18838 14118 18868 14170
rect 18868 14118 18880 14170
rect 18880 14118 18894 14170
rect 18918 14118 18932 14170
rect 18932 14118 18944 14170
rect 18944 14118 18974 14170
rect 18998 14118 19008 14170
rect 19008 14118 19054 14170
rect 18758 14116 18814 14118
rect 18838 14116 18894 14118
rect 18918 14116 18974 14118
rect 18998 14116 19054 14118
rect 18758 13082 18814 13084
rect 18838 13082 18894 13084
rect 18918 13082 18974 13084
rect 18998 13082 19054 13084
rect 18758 13030 18804 13082
rect 18804 13030 18814 13082
rect 18838 13030 18868 13082
rect 18868 13030 18880 13082
rect 18880 13030 18894 13082
rect 18918 13030 18932 13082
rect 18932 13030 18944 13082
rect 18944 13030 18974 13082
rect 18998 13030 19008 13082
rect 19008 13030 19054 13082
rect 18758 13028 18814 13030
rect 18838 13028 18894 13030
rect 18918 13028 18974 13030
rect 18998 13028 19054 13030
rect 17958 6160 18014 6216
rect 17958 5616 18014 5672
rect 17038 2760 17094 2816
rect 17958 4120 18014 4176
rect 18758 11994 18814 11996
rect 18838 11994 18894 11996
rect 18918 11994 18974 11996
rect 18998 11994 19054 11996
rect 18758 11942 18804 11994
rect 18804 11942 18814 11994
rect 18838 11942 18868 11994
rect 18868 11942 18880 11994
rect 18880 11942 18894 11994
rect 18918 11942 18932 11994
rect 18932 11942 18944 11994
rect 18944 11942 18974 11994
rect 18998 11942 19008 11994
rect 19008 11942 19054 11994
rect 18758 11940 18814 11942
rect 18838 11940 18894 11942
rect 18918 11940 18974 11942
rect 18998 11940 19054 11942
rect 19522 13404 19524 13424
rect 19524 13404 19576 13424
rect 19576 13404 19578 13424
rect 19522 13368 19578 13404
rect 21725 43002 21781 43004
rect 21805 43002 21861 43004
rect 21885 43002 21941 43004
rect 21965 43002 22021 43004
rect 21725 42950 21771 43002
rect 21771 42950 21781 43002
rect 21805 42950 21835 43002
rect 21835 42950 21847 43002
rect 21847 42950 21861 43002
rect 21885 42950 21899 43002
rect 21899 42950 21911 43002
rect 21911 42950 21941 43002
rect 21965 42950 21975 43002
rect 21975 42950 22021 43002
rect 21725 42948 21781 42950
rect 21805 42948 21861 42950
rect 21885 42948 21941 42950
rect 21965 42948 22021 42950
rect 21914 42084 21970 42120
rect 21914 42064 21916 42084
rect 21916 42064 21968 42084
rect 21968 42064 21970 42084
rect 21725 41914 21781 41916
rect 21805 41914 21861 41916
rect 21885 41914 21941 41916
rect 21965 41914 22021 41916
rect 21725 41862 21771 41914
rect 21771 41862 21781 41914
rect 21805 41862 21835 41914
rect 21835 41862 21847 41914
rect 21847 41862 21861 41914
rect 21885 41862 21899 41914
rect 21899 41862 21911 41914
rect 21911 41862 21941 41914
rect 21965 41862 21975 41914
rect 21975 41862 22021 41914
rect 21725 41860 21781 41862
rect 21805 41860 21861 41862
rect 21885 41860 21941 41862
rect 21965 41860 22021 41862
rect 21638 41556 21640 41576
rect 21640 41556 21692 41576
rect 21692 41556 21694 41576
rect 21638 41520 21694 41556
rect 21546 40976 21602 41032
rect 21730 41112 21786 41168
rect 21725 40826 21781 40828
rect 21805 40826 21861 40828
rect 21885 40826 21941 40828
rect 21965 40826 22021 40828
rect 21725 40774 21771 40826
rect 21771 40774 21781 40826
rect 21805 40774 21835 40826
rect 21835 40774 21847 40826
rect 21847 40774 21861 40826
rect 21885 40774 21899 40826
rect 21899 40774 21911 40826
rect 21911 40774 21941 40826
rect 21965 40774 21975 40826
rect 21975 40774 22021 40826
rect 21725 40772 21781 40774
rect 21805 40772 21861 40774
rect 21885 40772 21941 40774
rect 21965 40772 22021 40774
rect 21725 39738 21781 39740
rect 21805 39738 21861 39740
rect 21885 39738 21941 39740
rect 21965 39738 22021 39740
rect 21725 39686 21771 39738
rect 21771 39686 21781 39738
rect 21805 39686 21835 39738
rect 21835 39686 21847 39738
rect 21847 39686 21861 39738
rect 21885 39686 21899 39738
rect 21899 39686 21911 39738
rect 21911 39686 21941 39738
rect 21965 39686 21975 39738
rect 21975 39686 22021 39738
rect 21725 39684 21781 39686
rect 21805 39684 21861 39686
rect 21885 39684 21941 39686
rect 21965 39684 22021 39686
rect 22282 39888 22338 39944
rect 23202 43288 23258 43344
rect 22650 40568 22706 40624
rect 21822 38836 21824 38856
rect 21824 38836 21876 38856
rect 21876 38836 21878 38856
rect 21822 38800 21878 38836
rect 21725 38650 21781 38652
rect 21805 38650 21861 38652
rect 21885 38650 21941 38652
rect 21965 38650 22021 38652
rect 21725 38598 21771 38650
rect 21771 38598 21781 38650
rect 21805 38598 21835 38650
rect 21835 38598 21847 38650
rect 21847 38598 21861 38650
rect 21885 38598 21899 38650
rect 21899 38598 21911 38650
rect 21911 38598 21941 38650
rect 21965 38598 21975 38650
rect 21975 38598 22021 38650
rect 21725 38596 21781 38598
rect 21805 38596 21861 38598
rect 21885 38596 21941 38598
rect 21965 38596 22021 38598
rect 21725 37562 21781 37564
rect 21805 37562 21861 37564
rect 21885 37562 21941 37564
rect 21965 37562 22021 37564
rect 21725 37510 21771 37562
rect 21771 37510 21781 37562
rect 21805 37510 21835 37562
rect 21835 37510 21847 37562
rect 21847 37510 21861 37562
rect 21885 37510 21899 37562
rect 21899 37510 21911 37562
rect 21911 37510 21941 37562
rect 21965 37510 21975 37562
rect 21975 37510 22021 37562
rect 21725 37508 21781 37510
rect 21805 37508 21861 37510
rect 21885 37508 21941 37510
rect 21965 37508 22021 37510
rect 21725 36474 21781 36476
rect 21805 36474 21861 36476
rect 21885 36474 21941 36476
rect 21965 36474 22021 36476
rect 21725 36422 21771 36474
rect 21771 36422 21781 36474
rect 21805 36422 21835 36474
rect 21835 36422 21847 36474
rect 21847 36422 21861 36474
rect 21885 36422 21899 36474
rect 21899 36422 21911 36474
rect 21911 36422 21941 36474
rect 21965 36422 21975 36474
rect 21975 36422 22021 36474
rect 21725 36420 21781 36422
rect 21805 36420 21861 36422
rect 21885 36420 21941 36422
rect 21965 36420 22021 36422
rect 21725 35386 21781 35388
rect 21805 35386 21861 35388
rect 21885 35386 21941 35388
rect 21965 35386 22021 35388
rect 21725 35334 21771 35386
rect 21771 35334 21781 35386
rect 21805 35334 21835 35386
rect 21835 35334 21847 35386
rect 21847 35334 21861 35386
rect 21885 35334 21899 35386
rect 21899 35334 21911 35386
rect 21911 35334 21941 35386
rect 21965 35334 21975 35386
rect 21975 35334 22021 35386
rect 21725 35332 21781 35334
rect 21805 35332 21861 35334
rect 21885 35332 21941 35334
rect 21965 35332 22021 35334
rect 23570 42064 23626 42120
rect 22926 40468 22928 40488
rect 22928 40468 22980 40488
rect 22980 40468 22982 40488
rect 22926 40432 22982 40468
rect 23018 40160 23074 40216
rect 23110 40024 23166 40080
rect 23754 40976 23810 41032
rect 23662 40876 23664 40896
rect 23664 40876 23716 40896
rect 23716 40876 23718 40896
rect 23662 40840 23718 40876
rect 23662 40296 23718 40352
rect 24692 43546 24748 43548
rect 24772 43546 24828 43548
rect 24852 43546 24908 43548
rect 24932 43546 24988 43548
rect 24692 43494 24738 43546
rect 24738 43494 24748 43546
rect 24772 43494 24802 43546
rect 24802 43494 24814 43546
rect 24814 43494 24828 43546
rect 24852 43494 24866 43546
rect 24866 43494 24878 43546
rect 24878 43494 24908 43546
rect 24932 43494 24942 43546
rect 24942 43494 24988 43546
rect 24692 43492 24748 43494
rect 24772 43492 24828 43494
rect 24852 43492 24908 43494
rect 24932 43492 24988 43494
rect 24692 42458 24748 42460
rect 24772 42458 24828 42460
rect 24852 42458 24908 42460
rect 24932 42458 24988 42460
rect 24692 42406 24738 42458
rect 24738 42406 24748 42458
rect 24772 42406 24802 42458
rect 24802 42406 24814 42458
rect 24814 42406 24828 42458
rect 24852 42406 24866 42458
rect 24866 42406 24878 42458
rect 24878 42406 24908 42458
rect 24932 42406 24942 42458
rect 24942 42406 24988 42458
rect 24692 42404 24748 42406
rect 24772 42404 24828 42406
rect 24852 42404 24908 42406
rect 24932 42404 24988 42406
rect 24122 41928 24178 41984
rect 23202 39888 23258 39944
rect 23018 39480 23074 39536
rect 22834 39344 22890 39400
rect 22742 35944 22798 36000
rect 21725 34298 21781 34300
rect 21805 34298 21861 34300
rect 21885 34298 21941 34300
rect 21965 34298 22021 34300
rect 21725 34246 21771 34298
rect 21771 34246 21781 34298
rect 21805 34246 21835 34298
rect 21835 34246 21847 34298
rect 21847 34246 21861 34298
rect 21885 34246 21899 34298
rect 21899 34246 21911 34298
rect 21911 34246 21941 34298
rect 21965 34246 21975 34298
rect 21975 34246 22021 34298
rect 21725 34244 21781 34246
rect 21805 34244 21861 34246
rect 21885 34244 21941 34246
rect 21965 34244 22021 34246
rect 21546 31864 21602 31920
rect 22374 33496 22430 33552
rect 21725 33210 21781 33212
rect 21805 33210 21861 33212
rect 21885 33210 21941 33212
rect 21965 33210 22021 33212
rect 21725 33158 21771 33210
rect 21771 33158 21781 33210
rect 21805 33158 21835 33210
rect 21835 33158 21847 33210
rect 21847 33158 21861 33210
rect 21885 33158 21899 33210
rect 21899 33158 21911 33210
rect 21911 33158 21941 33210
rect 21965 33158 21975 33210
rect 21975 33158 22021 33210
rect 21725 33156 21781 33158
rect 21805 33156 21861 33158
rect 21885 33156 21941 33158
rect 21965 33156 22021 33158
rect 21725 32122 21781 32124
rect 21805 32122 21861 32124
rect 21885 32122 21941 32124
rect 21965 32122 22021 32124
rect 21725 32070 21771 32122
rect 21771 32070 21781 32122
rect 21805 32070 21835 32122
rect 21835 32070 21847 32122
rect 21847 32070 21861 32122
rect 21885 32070 21899 32122
rect 21899 32070 21911 32122
rect 21911 32070 21941 32122
rect 21965 32070 21975 32122
rect 21975 32070 22021 32122
rect 21725 32068 21781 32070
rect 21805 32068 21861 32070
rect 21885 32068 21941 32070
rect 21965 32068 22021 32070
rect 20810 26832 20866 26888
rect 20718 26324 20720 26344
rect 20720 26324 20772 26344
rect 20772 26324 20774 26344
rect 20718 26288 20774 26324
rect 21362 30368 21418 30424
rect 21725 31034 21781 31036
rect 21805 31034 21861 31036
rect 21885 31034 21941 31036
rect 21965 31034 22021 31036
rect 21725 30982 21771 31034
rect 21771 30982 21781 31034
rect 21805 30982 21835 31034
rect 21835 30982 21847 31034
rect 21847 30982 21861 31034
rect 21885 30982 21899 31034
rect 21899 30982 21911 31034
rect 21911 30982 21941 31034
rect 21965 30982 21975 31034
rect 21975 30982 22021 31034
rect 21725 30980 21781 30982
rect 21805 30980 21861 30982
rect 21885 30980 21941 30982
rect 21965 30980 22021 30982
rect 21725 29946 21781 29948
rect 21805 29946 21861 29948
rect 21885 29946 21941 29948
rect 21965 29946 22021 29948
rect 21725 29894 21771 29946
rect 21771 29894 21781 29946
rect 21805 29894 21835 29946
rect 21835 29894 21847 29946
rect 21847 29894 21861 29946
rect 21885 29894 21899 29946
rect 21899 29894 21911 29946
rect 21911 29894 21941 29946
rect 21965 29894 21975 29946
rect 21975 29894 22021 29946
rect 21725 29892 21781 29894
rect 21805 29892 21861 29894
rect 21885 29892 21941 29894
rect 21965 29892 22021 29894
rect 21725 28858 21781 28860
rect 21805 28858 21861 28860
rect 21885 28858 21941 28860
rect 21965 28858 22021 28860
rect 21725 28806 21771 28858
rect 21771 28806 21781 28858
rect 21805 28806 21835 28858
rect 21835 28806 21847 28858
rect 21847 28806 21861 28858
rect 21885 28806 21899 28858
rect 21899 28806 21911 28858
rect 21911 28806 21941 28858
rect 21965 28806 21975 28858
rect 21975 28806 22021 28858
rect 21725 28804 21781 28806
rect 21805 28804 21861 28806
rect 21885 28804 21941 28806
rect 21965 28804 22021 28806
rect 22190 28092 22192 28112
rect 22192 28092 22244 28112
rect 22244 28092 22246 28112
rect 22190 28056 22246 28092
rect 21725 27770 21781 27772
rect 21805 27770 21861 27772
rect 21885 27770 21941 27772
rect 21965 27770 22021 27772
rect 21725 27718 21771 27770
rect 21771 27718 21781 27770
rect 21805 27718 21835 27770
rect 21835 27718 21847 27770
rect 21847 27718 21861 27770
rect 21885 27718 21899 27770
rect 21899 27718 21911 27770
rect 21911 27718 21941 27770
rect 21965 27718 21975 27770
rect 21975 27718 22021 27770
rect 21725 27716 21781 27718
rect 21805 27716 21861 27718
rect 21885 27716 21941 27718
rect 21965 27716 22021 27718
rect 19982 16360 20038 16416
rect 19430 11736 19486 11792
rect 18758 10906 18814 10908
rect 18838 10906 18894 10908
rect 18918 10906 18974 10908
rect 18998 10906 19054 10908
rect 18758 10854 18804 10906
rect 18804 10854 18814 10906
rect 18838 10854 18868 10906
rect 18868 10854 18880 10906
rect 18880 10854 18894 10906
rect 18918 10854 18932 10906
rect 18932 10854 18944 10906
rect 18944 10854 18974 10906
rect 18998 10854 19008 10906
rect 19008 10854 19054 10906
rect 18758 10852 18814 10854
rect 18838 10852 18894 10854
rect 18918 10852 18974 10854
rect 18998 10852 19054 10854
rect 19246 11056 19302 11112
rect 18758 9818 18814 9820
rect 18838 9818 18894 9820
rect 18918 9818 18974 9820
rect 18998 9818 19054 9820
rect 18758 9766 18804 9818
rect 18804 9766 18814 9818
rect 18838 9766 18868 9818
rect 18868 9766 18880 9818
rect 18880 9766 18894 9818
rect 18918 9766 18932 9818
rect 18932 9766 18944 9818
rect 18944 9766 18974 9818
rect 18998 9766 19008 9818
rect 19008 9766 19054 9818
rect 18758 9764 18814 9766
rect 18838 9764 18894 9766
rect 18918 9764 18974 9766
rect 18998 9764 19054 9766
rect 18758 8730 18814 8732
rect 18838 8730 18894 8732
rect 18918 8730 18974 8732
rect 18998 8730 19054 8732
rect 18758 8678 18804 8730
rect 18804 8678 18814 8730
rect 18838 8678 18868 8730
rect 18868 8678 18880 8730
rect 18880 8678 18894 8730
rect 18918 8678 18932 8730
rect 18932 8678 18944 8730
rect 18944 8678 18974 8730
rect 18998 8678 19008 8730
rect 19008 8678 19054 8730
rect 18758 8676 18814 8678
rect 18838 8676 18894 8678
rect 18918 8676 18974 8678
rect 18998 8676 19054 8678
rect 18694 8472 18750 8528
rect 18758 7642 18814 7644
rect 18838 7642 18894 7644
rect 18918 7642 18974 7644
rect 18998 7642 19054 7644
rect 18758 7590 18804 7642
rect 18804 7590 18814 7642
rect 18838 7590 18868 7642
rect 18868 7590 18880 7642
rect 18880 7590 18894 7642
rect 18918 7590 18932 7642
rect 18932 7590 18944 7642
rect 18944 7590 18974 7642
rect 18998 7590 19008 7642
rect 19008 7590 19054 7642
rect 18758 7588 18814 7590
rect 18838 7588 18894 7590
rect 18918 7588 18974 7590
rect 18998 7588 19054 7590
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 19062 5072 19118 5128
rect 19430 10804 19486 10840
rect 19430 10784 19432 10804
rect 19432 10784 19484 10804
rect 19484 10784 19486 10804
rect 19338 10698 19394 10704
rect 19338 10648 19340 10698
rect 19340 10648 19392 10698
rect 19392 10648 19394 10698
rect 19706 10784 19762 10840
rect 19430 6704 19486 6760
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18326 3984 18382 4040
rect 18234 3848 18290 3904
rect 18234 3440 18290 3496
rect 17222 2624 17278 2680
rect 16486 1300 16488 1320
rect 16488 1300 16540 1320
rect 16540 1300 16542 1320
rect 16486 1264 16542 1300
rect 17498 2624 17554 2680
rect 17958 2896 18014 2952
rect 17958 2624 18014 2680
rect 18142 3304 18198 3360
rect 18694 3712 18750 3768
rect 19154 3712 19210 3768
rect 18142 2352 18198 2408
rect 18602 3340 18604 3360
rect 18604 3340 18656 3360
rect 18656 3340 18658 3360
rect 18602 3304 18658 3340
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 19154 3168 19210 3224
rect 18694 2916 18750 2952
rect 18694 2896 18696 2916
rect 18696 2896 18748 2916
rect 18748 2896 18750 2916
rect 18510 2624 18566 2680
rect 18694 2624 18750 2680
rect 18602 2388 18604 2408
rect 18604 2388 18656 2408
rect 18656 2388 18658 2408
rect 18602 2352 18658 2388
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 20718 17992 20774 18048
rect 20626 15000 20682 15056
rect 19522 3984 19578 4040
rect 19430 2624 19486 2680
rect 20258 5344 20314 5400
rect 21725 26682 21781 26684
rect 21805 26682 21861 26684
rect 21885 26682 21941 26684
rect 21965 26682 22021 26684
rect 21725 26630 21771 26682
rect 21771 26630 21781 26682
rect 21805 26630 21835 26682
rect 21835 26630 21847 26682
rect 21847 26630 21861 26682
rect 21885 26630 21899 26682
rect 21899 26630 21911 26682
rect 21911 26630 21941 26682
rect 21965 26630 21975 26682
rect 21975 26630 22021 26682
rect 21725 26628 21781 26630
rect 21805 26628 21861 26630
rect 21885 26628 21941 26630
rect 21965 26628 22021 26630
rect 21725 25594 21781 25596
rect 21805 25594 21861 25596
rect 21885 25594 21941 25596
rect 21965 25594 22021 25596
rect 21725 25542 21771 25594
rect 21771 25542 21781 25594
rect 21805 25542 21835 25594
rect 21835 25542 21847 25594
rect 21847 25542 21861 25594
rect 21885 25542 21899 25594
rect 21899 25542 21911 25594
rect 21911 25542 21941 25594
rect 21965 25542 21975 25594
rect 21975 25542 22021 25594
rect 21725 25540 21781 25542
rect 21805 25540 21861 25542
rect 21885 25540 21941 25542
rect 21965 25540 22021 25542
rect 21730 24792 21786 24848
rect 21725 24506 21781 24508
rect 21805 24506 21861 24508
rect 21885 24506 21941 24508
rect 21965 24506 22021 24508
rect 21725 24454 21771 24506
rect 21771 24454 21781 24506
rect 21805 24454 21835 24506
rect 21835 24454 21847 24506
rect 21847 24454 21861 24506
rect 21885 24454 21899 24506
rect 21899 24454 21911 24506
rect 21911 24454 21941 24506
rect 21965 24454 21975 24506
rect 21975 24454 22021 24506
rect 21725 24452 21781 24454
rect 21805 24452 21861 24454
rect 21885 24452 21941 24454
rect 21965 24452 22021 24454
rect 21725 23418 21781 23420
rect 21805 23418 21861 23420
rect 21885 23418 21941 23420
rect 21965 23418 22021 23420
rect 21725 23366 21771 23418
rect 21771 23366 21781 23418
rect 21805 23366 21835 23418
rect 21835 23366 21847 23418
rect 21847 23366 21861 23418
rect 21885 23366 21899 23418
rect 21899 23366 21911 23418
rect 21911 23366 21941 23418
rect 21965 23366 21975 23418
rect 21975 23366 22021 23418
rect 21725 23364 21781 23366
rect 21805 23364 21861 23366
rect 21885 23364 21941 23366
rect 21965 23364 22021 23366
rect 21730 22480 21786 22536
rect 21725 22330 21781 22332
rect 21805 22330 21861 22332
rect 21885 22330 21941 22332
rect 21965 22330 22021 22332
rect 21725 22278 21771 22330
rect 21771 22278 21781 22330
rect 21805 22278 21835 22330
rect 21835 22278 21847 22330
rect 21847 22278 21861 22330
rect 21885 22278 21899 22330
rect 21899 22278 21911 22330
rect 21911 22278 21941 22330
rect 21965 22278 21975 22330
rect 21975 22278 22021 22330
rect 21725 22276 21781 22278
rect 21805 22276 21861 22278
rect 21885 22276 21941 22278
rect 21965 22276 22021 22278
rect 21546 19896 21602 19952
rect 22558 33360 22614 33416
rect 24122 37168 24178 37224
rect 22190 21392 22246 21448
rect 21725 21242 21781 21244
rect 21805 21242 21861 21244
rect 21885 21242 21941 21244
rect 21965 21242 22021 21244
rect 21725 21190 21771 21242
rect 21771 21190 21781 21242
rect 21805 21190 21835 21242
rect 21835 21190 21847 21242
rect 21847 21190 21861 21242
rect 21885 21190 21899 21242
rect 21899 21190 21911 21242
rect 21911 21190 21941 21242
rect 21965 21190 21975 21242
rect 21975 21190 22021 21242
rect 21725 21188 21781 21190
rect 21805 21188 21861 21190
rect 21885 21188 21941 21190
rect 21965 21188 22021 21190
rect 21725 20154 21781 20156
rect 21805 20154 21861 20156
rect 21885 20154 21941 20156
rect 21965 20154 22021 20156
rect 21725 20102 21771 20154
rect 21771 20102 21781 20154
rect 21805 20102 21835 20154
rect 21835 20102 21847 20154
rect 21847 20102 21861 20154
rect 21885 20102 21899 20154
rect 21899 20102 21911 20154
rect 21911 20102 21941 20154
rect 21965 20102 21975 20154
rect 21975 20102 22021 20154
rect 21725 20100 21781 20102
rect 21805 20100 21861 20102
rect 21885 20100 21941 20102
rect 21965 20100 22021 20102
rect 21725 19066 21781 19068
rect 21805 19066 21861 19068
rect 21885 19066 21941 19068
rect 21965 19066 22021 19068
rect 21725 19014 21771 19066
rect 21771 19014 21781 19066
rect 21805 19014 21835 19066
rect 21835 19014 21847 19066
rect 21847 19014 21861 19066
rect 21885 19014 21899 19066
rect 21899 19014 21911 19066
rect 21911 19014 21941 19066
rect 21965 19014 21975 19066
rect 21975 19014 22021 19066
rect 21725 19012 21781 19014
rect 21805 19012 21861 19014
rect 21885 19012 21941 19014
rect 21965 19012 22021 19014
rect 21638 18264 21694 18320
rect 21725 17978 21781 17980
rect 21805 17978 21861 17980
rect 21885 17978 21941 17980
rect 21965 17978 22021 17980
rect 21725 17926 21771 17978
rect 21771 17926 21781 17978
rect 21805 17926 21835 17978
rect 21835 17926 21847 17978
rect 21847 17926 21861 17978
rect 21885 17926 21899 17978
rect 21899 17926 21911 17978
rect 21911 17926 21941 17978
rect 21965 17926 21975 17978
rect 21975 17926 22021 17978
rect 21725 17924 21781 17926
rect 21805 17924 21861 17926
rect 21885 17924 21941 17926
rect 21965 17924 22021 17926
rect 22466 22480 22522 22536
rect 22282 19896 22338 19952
rect 22742 19760 22798 19816
rect 24398 39788 24400 39808
rect 24400 39788 24452 39808
rect 24452 39788 24454 39808
rect 24398 39752 24454 39788
rect 24398 38700 24400 38720
rect 24400 38700 24452 38720
rect 24452 38700 24454 38720
rect 24398 38664 24454 38700
rect 24398 37612 24400 37632
rect 24400 37612 24452 37632
rect 24452 37612 24454 37632
rect 24398 37576 24454 37612
rect 24398 36524 24400 36544
rect 24400 36524 24452 36544
rect 24452 36524 24454 36544
rect 24398 36488 24454 36524
rect 24398 35436 24400 35456
rect 24400 35436 24452 35456
rect 24452 35436 24454 35456
rect 24398 35400 24454 35436
rect 24398 34484 24400 34504
rect 24400 34484 24452 34504
rect 24452 34484 24454 34504
rect 24398 34448 24454 34484
rect 24398 33260 24400 33280
rect 24400 33260 24452 33280
rect 24452 33260 24454 33280
rect 24398 33224 24454 33260
rect 24398 32172 24400 32192
rect 24400 32172 24452 32192
rect 24452 32172 24454 32192
rect 24398 32136 24454 32172
rect 23570 23568 23626 23624
rect 21546 17448 21602 17504
rect 20902 14864 20958 14920
rect 20810 10648 20866 10704
rect 20810 9832 20866 9888
rect 21270 12688 21326 12744
rect 21178 12280 21234 12336
rect 22282 17720 22338 17776
rect 21725 16890 21781 16892
rect 21805 16890 21861 16892
rect 21885 16890 21941 16892
rect 21965 16890 22021 16892
rect 21725 16838 21771 16890
rect 21771 16838 21781 16890
rect 21805 16838 21835 16890
rect 21835 16838 21847 16890
rect 21847 16838 21861 16890
rect 21885 16838 21899 16890
rect 21899 16838 21911 16890
rect 21911 16838 21941 16890
rect 21965 16838 21975 16890
rect 21975 16838 22021 16890
rect 21725 16836 21781 16838
rect 21805 16836 21861 16838
rect 21885 16836 21941 16838
rect 21965 16836 22021 16838
rect 21725 15802 21781 15804
rect 21805 15802 21861 15804
rect 21885 15802 21941 15804
rect 21965 15802 22021 15804
rect 21725 15750 21771 15802
rect 21771 15750 21781 15802
rect 21805 15750 21835 15802
rect 21835 15750 21847 15802
rect 21847 15750 21861 15802
rect 21885 15750 21899 15802
rect 21899 15750 21911 15802
rect 21911 15750 21941 15802
rect 21965 15750 21975 15802
rect 21975 15750 22021 15802
rect 21725 15748 21781 15750
rect 21805 15748 21861 15750
rect 21885 15748 21941 15750
rect 21965 15748 22021 15750
rect 21725 14714 21781 14716
rect 21805 14714 21861 14716
rect 21885 14714 21941 14716
rect 21965 14714 22021 14716
rect 21725 14662 21771 14714
rect 21771 14662 21781 14714
rect 21805 14662 21835 14714
rect 21835 14662 21847 14714
rect 21847 14662 21861 14714
rect 21885 14662 21899 14714
rect 21899 14662 21911 14714
rect 21911 14662 21941 14714
rect 21965 14662 21975 14714
rect 21975 14662 22021 14714
rect 21725 14660 21781 14662
rect 21805 14660 21861 14662
rect 21885 14660 21941 14662
rect 21965 14660 22021 14662
rect 21725 13626 21781 13628
rect 21805 13626 21861 13628
rect 21885 13626 21941 13628
rect 21965 13626 22021 13628
rect 21725 13574 21771 13626
rect 21771 13574 21781 13626
rect 21805 13574 21835 13626
rect 21835 13574 21847 13626
rect 21847 13574 21861 13626
rect 21885 13574 21899 13626
rect 21899 13574 21911 13626
rect 21911 13574 21941 13626
rect 21965 13574 21975 13626
rect 21975 13574 22021 13626
rect 21725 13572 21781 13574
rect 21805 13572 21861 13574
rect 21885 13572 21941 13574
rect 21965 13572 22021 13574
rect 23846 21292 23848 21312
rect 23848 21292 23900 21312
rect 23900 21292 23902 21312
rect 23846 21256 23902 21292
rect 24030 20168 24086 20224
rect 24398 31084 24400 31104
rect 24400 31084 24452 31104
rect 24452 31084 24454 31104
rect 24398 31048 24454 31084
rect 24692 41370 24748 41372
rect 24772 41370 24828 41372
rect 24852 41370 24908 41372
rect 24932 41370 24988 41372
rect 24692 41318 24738 41370
rect 24738 41318 24748 41370
rect 24772 41318 24802 41370
rect 24802 41318 24814 41370
rect 24814 41318 24828 41370
rect 24852 41318 24866 41370
rect 24866 41318 24878 41370
rect 24878 41318 24908 41370
rect 24932 41318 24942 41370
rect 24942 41318 24988 41370
rect 24692 41316 24748 41318
rect 24772 41316 24828 41318
rect 24852 41316 24908 41318
rect 24932 41316 24988 41318
rect 25318 43016 25374 43072
rect 25134 42472 25190 42528
rect 25226 41384 25282 41440
rect 25134 40296 25190 40352
rect 24692 40282 24748 40284
rect 24772 40282 24828 40284
rect 24852 40282 24908 40284
rect 24932 40282 24988 40284
rect 24692 40230 24738 40282
rect 24738 40230 24748 40282
rect 24772 40230 24802 40282
rect 24802 40230 24814 40282
rect 24814 40230 24828 40282
rect 24852 40230 24866 40282
rect 24866 40230 24878 40282
rect 24878 40230 24908 40282
rect 24932 40230 24942 40282
rect 24942 40230 24988 40282
rect 24692 40228 24748 40230
rect 24772 40228 24828 40230
rect 24852 40228 24908 40230
rect 24932 40228 24988 40230
rect 25226 39244 25228 39264
rect 25228 39244 25280 39264
rect 25280 39244 25282 39264
rect 25226 39208 25282 39244
rect 24692 39194 24748 39196
rect 24772 39194 24828 39196
rect 24852 39194 24908 39196
rect 24932 39194 24988 39196
rect 24692 39142 24738 39194
rect 24738 39142 24748 39194
rect 24772 39142 24802 39194
rect 24802 39142 24814 39194
rect 24814 39142 24828 39194
rect 24852 39142 24866 39194
rect 24866 39142 24878 39194
rect 24878 39142 24908 39194
rect 24932 39142 24942 39194
rect 24942 39142 24988 39194
rect 24692 39140 24748 39142
rect 24772 39140 24828 39142
rect 24852 39140 24908 39142
rect 24932 39140 24988 39142
rect 25226 38156 25228 38176
rect 25228 38156 25280 38176
rect 25280 38156 25282 38176
rect 25226 38120 25282 38156
rect 24692 38106 24748 38108
rect 24772 38106 24828 38108
rect 24852 38106 24908 38108
rect 24932 38106 24988 38108
rect 24692 38054 24738 38106
rect 24738 38054 24748 38106
rect 24772 38054 24802 38106
rect 24802 38054 24814 38106
rect 24814 38054 24828 38106
rect 24852 38054 24866 38106
rect 24866 38054 24878 38106
rect 24878 38054 24908 38106
rect 24932 38054 24942 38106
rect 24942 38054 24988 38106
rect 24692 38052 24748 38054
rect 24772 38052 24828 38054
rect 24852 38052 24908 38054
rect 24932 38052 24988 38054
rect 24692 37018 24748 37020
rect 24772 37018 24828 37020
rect 24852 37018 24908 37020
rect 24932 37018 24988 37020
rect 24692 36966 24738 37018
rect 24738 36966 24748 37018
rect 24772 36966 24802 37018
rect 24802 36966 24814 37018
rect 24814 36966 24828 37018
rect 24852 36966 24866 37018
rect 24866 36966 24878 37018
rect 24878 36966 24908 37018
rect 24932 36966 24942 37018
rect 24942 36966 24988 37018
rect 24692 36964 24748 36966
rect 24772 36964 24828 36966
rect 24852 36964 24908 36966
rect 24932 36964 24988 36966
rect 25134 35944 25190 36000
rect 24692 35930 24748 35932
rect 24772 35930 24828 35932
rect 24852 35930 24908 35932
rect 24932 35930 24988 35932
rect 24692 35878 24738 35930
rect 24738 35878 24748 35930
rect 24772 35878 24802 35930
rect 24802 35878 24814 35930
rect 24814 35878 24828 35930
rect 24852 35878 24866 35930
rect 24866 35878 24878 35930
rect 24878 35878 24908 35930
rect 24932 35878 24942 35930
rect 24942 35878 24988 35930
rect 24692 35876 24748 35878
rect 24772 35876 24828 35878
rect 24852 35876 24908 35878
rect 24932 35876 24988 35878
rect 24692 34842 24748 34844
rect 24772 34842 24828 34844
rect 24852 34842 24908 34844
rect 24932 34842 24988 34844
rect 24692 34790 24738 34842
rect 24738 34790 24748 34842
rect 24772 34790 24802 34842
rect 24802 34790 24814 34842
rect 24814 34790 24828 34842
rect 24852 34790 24866 34842
rect 24866 34790 24878 34842
rect 24878 34790 24908 34842
rect 24932 34790 24942 34842
rect 24942 34790 24988 34842
rect 24692 34788 24748 34790
rect 24772 34788 24828 34790
rect 24852 34788 24908 34790
rect 24932 34788 24988 34790
rect 24692 33754 24748 33756
rect 24772 33754 24828 33756
rect 24852 33754 24908 33756
rect 24932 33754 24988 33756
rect 24692 33702 24738 33754
rect 24738 33702 24748 33754
rect 24772 33702 24802 33754
rect 24802 33702 24814 33754
rect 24814 33702 24828 33754
rect 24852 33702 24866 33754
rect 24866 33702 24878 33754
rect 24878 33702 24908 33754
rect 24932 33702 24942 33754
rect 24942 33702 24988 33754
rect 24692 33700 24748 33702
rect 24772 33700 24828 33702
rect 24852 33700 24908 33702
rect 24932 33700 24988 33702
rect 24692 32666 24748 32668
rect 24772 32666 24828 32668
rect 24852 32666 24908 32668
rect 24932 32666 24988 32668
rect 24692 32614 24738 32666
rect 24738 32614 24748 32666
rect 24772 32614 24802 32666
rect 24802 32614 24814 32666
rect 24814 32614 24828 32666
rect 24852 32614 24866 32666
rect 24866 32614 24878 32666
rect 24878 32614 24908 32666
rect 24932 32614 24942 32666
rect 24942 32614 24988 32666
rect 24692 32612 24748 32614
rect 24772 32612 24828 32614
rect 24852 32612 24908 32614
rect 24932 32612 24988 32614
rect 24692 31578 24748 31580
rect 24772 31578 24828 31580
rect 24852 31578 24908 31580
rect 24932 31578 24988 31580
rect 24692 31526 24738 31578
rect 24738 31526 24748 31578
rect 24772 31526 24802 31578
rect 24802 31526 24814 31578
rect 24814 31526 24828 31578
rect 24852 31526 24866 31578
rect 24866 31526 24878 31578
rect 24878 31526 24908 31578
rect 24932 31526 24942 31578
rect 24942 31526 24988 31578
rect 24692 31524 24748 31526
rect 24772 31524 24828 31526
rect 24852 31524 24908 31526
rect 24932 31524 24988 31526
rect 24398 29996 24400 30016
rect 24400 29996 24452 30016
rect 24452 29996 24454 30016
rect 24398 29960 24454 29996
rect 24398 28908 24400 28928
rect 24400 28908 24452 28928
rect 24452 28908 24454 28928
rect 24398 28872 24454 28908
rect 24398 27820 24400 27840
rect 24400 27820 24452 27840
rect 24452 27820 24454 27840
rect 24398 27784 24454 27820
rect 24398 26732 24400 26752
rect 24400 26732 24452 26752
rect 24452 26732 24454 26752
rect 24398 26696 24454 26732
rect 24398 25644 24400 25664
rect 24400 25644 24452 25664
rect 24452 25644 24454 25664
rect 24398 25608 24454 25644
rect 23846 19116 23848 19136
rect 23848 19116 23900 19136
rect 23900 19116 23902 19136
rect 23846 19080 23902 19116
rect 23018 17176 23074 17232
rect 22190 13640 22246 13696
rect 21725 12538 21781 12540
rect 21805 12538 21861 12540
rect 21885 12538 21941 12540
rect 21965 12538 22021 12540
rect 21725 12486 21771 12538
rect 21771 12486 21781 12538
rect 21805 12486 21835 12538
rect 21835 12486 21847 12538
rect 21847 12486 21861 12538
rect 21885 12486 21899 12538
rect 21899 12486 21911 12538
rect 21911 12486 21941 12538
rect 21965 12486 21975 12538
rect 21975 12486 22021 12538
rect 21725 12484 21781 12486
rect 21805 12484 21861 12486
rect 21885 12484 21941 12486
rect 21965 12484 22021 12486
rect 20718 6840 20774 6896
rect 20718 5208 20774 5264
rect 19798 2624 19854 2680
rect 20534 3848 20590 3904
rect 20902 6432 20958 6488
rect 20902 6060 20904 6080
rect 20904 6060 20956 6080
rect 20956 6060 20958 6080
rect 20902 6024 20958 6060
rect 21086 6432 21142 6488
rect 21454 6840 21510 6896
rect 21725 11450 21781 11452
rect 21805 11450 21861 11452
rect 21885 11450 21941 11452
rect 21965 11450 22021 11452
rect 21725 11398 21771 11450
rect 21771 11398 21781 11450
rect 21805 11398 21835 11450
rect 21835 11398 21847 11450
rect 21847 11398 21861 11450
rect 21885 11398 21899 11450
rect 21899 11398 21911 11450
rect 21911 11398 21941 11450
rect 21965 11398 21975 11450
rect 21975 11398 22021 11450
rect 21725 11396 21781 11398
rect 21805 11396 21861 11398
rect 21885 11396 21941 11398
rect 21965 11396 22021 11398
rect 22558 12552 22614 12608
rect 21725 10362 21781 10364
rect 21805 10362 21861 10364
rect 21885 10362 21941 10364
rect 21965 10362 22021 10364
rect 21725 10310 21771 10362
rect 21771 10310 21781 10362
rect 21805 10310 21835 10362
rect 21835 10310 21847 10362
rect 21847 10310 21861 10362
rect 21885 10310 21899 10362
rect 21899 10310 21911 10362
rect 21911 10310 21941 10362
rect 21965 10310 21975 10362
rect 21975 10310 22021 10362
rect 21725 10308 21781 10310
rect 21805 10308 21861 10310
rect 21885 10308 21941 10310
rect 21965 10308 22021 10310
rect 21725 9274 21781 9276
rect 21805 9274 21861 9276
rect 21885 9274 21941 9276
rect 21965 9274 22021 9276
rect 21725 9222 21771 9274
rect 21771 9222 21781 9274
rect 21805 9222 21835 9274
rect 21835 9222 21847 9274
rect 21847 9222 21861 9274
rect 21885 9222 21899 9274
rect 21899 9222 21911 9274
rect 21911 9222 21941 9274
rect 21965 9222 21975 9274
rect 21975 9222 22021 9274
rect 21725 9220 21781 9222
rect 21805 9220 21861 9222
rect 21885 9220 21941 9222
rect 21965 9220 22021 9222
rect 21725 8186 21781 8188
rect 21805 8186 21861 8188
rect 21885 8186 21941 8188
rect 21965 8186 22021 8188
rect 21725 8134 21771 8186
rect 21771 8134 21781 8186
rect 21805 8134 21835 8186
rect 21835 8134 21847 8186
rect 21847 8134 21861 8186
rect 21885 8134 21899 8186
rect 21899 8134 21911 8186
rect 21911 8134 21941 8186
rect 21965 8134 21975 8186
rect 21975 8134 22021 8186
rect 21725 8132 21781 8134
rect 21805 8132 21861 8134
rect 21885 8132 21941 8134
rect 21965 8132 22021 8134
rect 21725 7098 21781 7100
rect 21805 7098 21861 7100
rect 21885 7098 21941 7100
rect 21965 7098 22021 7100
rect 21725 7046 21771 7098
rect 21771 7046 21781 7098
rect 21805 7046 21835 7098
rect 21835 7046 21847 7098
rect 21847 7046 21861 7098
rect 21885 7046 21899 7098
rect 21899 7046 21911 7098
rect 21911 7046 21941 7098
rect 21965 7046 21975 7098
rect 21975 7046 22021 7098
rect 21725 7044 21781 7046
rect 21805 7044 21861 7046
rect 21885 7044 21941 7046
rect 21965 7044 22021 7046
rect 21822 6704 21878 6760
rect 21362 6160 21418 6216
rect 20902 3984 20958 4040
rect 20810 3576 20866 3632
rect 20718 2916 20774 2952
rect 20718 2896 20720 2916
rect 20720 2896 20772 2916
rect 20772 2896 20774 2916
rect 20718 2760 20774 2816
rect 20442 584 20498 640
rect 21914 6160 21970 6216
rect 21546 6024 21602 6080
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 22282 6160 22338 6216
rect 22098 5752 22154 5808
rect 21270 3440 21326 3496
rect 22006 5072 22062 5128
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 21546 4664 21602 4720
rect 21454 3984 21510 4040
rect 24398 24556 24400 24576
rect 24400 24556 24452 24576
rect 24452 24556 24454 24576
rect 24398 24520 24454 24556
rect 24398 23468 24400 23488
rect 24400 23468 24452 23488
rect 24452 23468 24454 23488
rect 24398 23432 24454 23468
rect 24490 22344 24546 22400
rect 24398 18028 24400 18048
rect 24400 18028 24452 18048
rect 24452 18028 24454 18048
rect 24398 17992 24454 18028
rect 24122 16940 24124 16960
rect 24124 16940 24176 16960
rect 24176 16940 24178 16960
rect 24122 16904 24178 16940
rect 23938 16496 23994 16552
rect 23018 12552 23074 12608
rect 23478 13368 23534 13424
rect 24122 15816 24178 15872
rect 24030 14764 24032 14784
rect 24032 14764 24084 14784
rect 24084 14764 24086 14784
rect 24030 14728 24086 14764
rect 24214 12588 24216 12608
rect 24216 12588 24268 12608
rect 24268 12588 24270 12608
rect 24214 12552 24270 12588
rect 23846 11500 23848 11520
rect 23848 11500 23900 11520
rect 23900 11500 23902 11520
rect 23846 11464 23902 11500
rect 22742 5480 22798 5536
rect 21362 1420 21418 1456
rect 21362 1400 21364 1420
rect 21364 1400 21416 1420
rect 21416 1400 21418 1420
rect 21086 1264 21142 1320
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 22650 4120 22706 4176
rect 22650 3032 22706 3088
rect 23386 10376 23442 10432
rect 23570 8916 23572 8936
rect 23572 8916 23624 8936
rect 23624 8916 23626 8936
rect 23570 8880 23626 8916
rect 24030 9288 24086 9344
rect 23202 6740 23204 6760
rect 23204 6740 23256 6760
rect 23256 6740 23258 6760
rect 23202 6704 23258 6740
rect 23754 7112 23810 7168
rect 23662 6840 23718 6896
rect 23386 6452 23442 6488
rect 23386 6432 23388 6452
rect 23388 6432 23440 6452
rect 23440 6432 23442 6452
rect 23386 6296 23442 6352
rect 23386 5480 23442 5536
rect 24692 30490 24748 30492
rect 24772 30490 24828 30492
rect 24852 30490 24908 30492
rect 24932 30490 24988 30492
rect 24692 30438 24738 30490
rect 24738 30438 24748 30490
rect 24772 30438 24802 30490
rect 24802 30438 24814 30490
rect 24814 30438 24828 30490
rect 24852 30438 24866 30490
rect 24866 30438 24878 30490
rect 24878 30438 24908 30490
rect 24932 30438 24942 30490
rect 24942 30438 24988 30490
rect 24692 30436 24748 30438
rect 24772 30436 24828 30438
rect 24852 30436 24908 30438
rect 24932 30436 24988 30438
rect 24692 29402 24748 29404
rect 24772 29402 24828 29404
rect 24852 29402 24908 29404
rect 24932 29402 24988 29404
rect 24692 29350 24738 29402
rect 24738 29350 24748 29402
rect 24772 29350 24802 29402
rect 24802 29350 24814 29402
rect 24814 29350 24828 29402
rect 24852 29350 24866 29402
rect 24866 29350 24878 29402
rect 24878 29350 24908 29402
rect 24932 29350 24942 29402
rect 24942 29350 24988 29402
rect 24692 29348 24748 29350
rect 24772 29348 24828 29350
rect 24852 29348 24908 29350
rect 24932 29348 24988 29350
rect 24692 28314 24748 28316
rect 24772 28314 24828 28316
rect 24852 28314 24908 28316
rect 24932 28314 24988 28316
rect 24692 28262 24738 28314
rect 24738 28262 24748 28314
rect 24772 28262 24802 28314
rect 24802 28262 24814 28314
rect 24814 28262 24828 28314
rect 24852 28262 24866 28314
rect 24866 28262 24878 28314
rect 24878 28262 24908 28314
rect 24932 28262 24942 28314
rect 24942 28262 24988 28314
rect 24692 28260 24748 28262
rect 24772 28260 24828 28262
rect 24852 28260 24908 28262
rect 24932 28260 24988 28262
rect 24692 27226 24748 27228
rect 24772 27226 24828 27228
rect 24852 27226 24908 27228
rect 24932 27226 24988 27228
rect 24692 27174 24738 27226
rect 24738 27174 24748 27226
rect 24772 27174 24802 27226
rect 24802 27174 24814 27226
rect 24814 27174 24828 27226
rect 24852 27174 24866 27226
rect 24866 27174 24878 27226
rect 24878 27174 24908 27226
rect 24932 27174 24942 27226
rect 24942 27174 24988 27226
rect 24692 27172 24748 27174
rect 24772 27172 24828 27174
rect 24852 27172 24908 27174
rect 24932 27172 24988 27174
rect 24692 26138 24748 26140
rect 24772 26138 24828 26140
rect 24852 26138 24908 26140
rect 24932 26138 24988 26140
rect 24692 26086 24738 26138
rect 24738 26086 24748 26138
rect 24772 26086 24802 26138
rect 24802 26086 24814 26138
rect 24814 26086 24828 26138
rect 24852 26086 24866 26138
rect 24866 26086 24878 26138
rect 24878 26086 24908 26138
rect 24932 26086 24942 26138
rect 24942 26086 24988 26138
rect 24692 26084 24748 26086
rect 24772 26084 24828 26086
rect 24852 26084 24908 26086
rect 24932 26084 24988 26086
rect 24692 25050 24748 25052
rect 24772 25050 24828 25052
rect 24852 25050 24908 25052
rect 24932 25050 24988 25052
rect 24692 24998 24738 25050
rect 24738 24998 24748 25050
rect 24772 24998 24802 25050
rect 24802 24998 24814 25050
rect 24814 24998 24828 25050
rect 24852 24998 24866 25050
rect 24866 24998 24878 25050
rect 24878 24998 24908 25050
rect 24932 24998 24942 25050
rect 24942 24998 24988 25050
rect 24692 24996 24748 24998
rect 24772 24996 24828 24998
rect 24852 24996 24908 24998
rect 24932 24996 24988 24998
rect 24692 23962 24748 23964
rect 24772 23962 24828 23964
rect 24852 23962 24908 23964
rect 24932 23962 24988 23964
rect 24692 23910 24738 23962
rect 24738 23910 24748 23962
rect 24772 23910 24802 23962
rect 24802 23910 24814 23962
rect 24814 23910 24828 23962
rect 24852 23910 24866 23962
rect 24866 23910 24878 23962
rect 24878 23910 24908 23962
rect 24932 23910 24942 23962
rect 24942 23910 24988 23962
rect 24692 23908 24748 23910
rect 24772 23908 24828 23910
rect 24852 23908 24908 23910
rect 24932 23908 24988 23910
rect 24692 22874 24748 22876
rect 24772 22874 24828 22876
rect 24852 22874 24908 22876
rect 24932 22874 24988 22876
rect 24692 22822 24738 22874
rect 24738 22822 24748 22874
rect 24772 22822 24802 22874
rect 24802 22822 24814 22874
rect 24814 22822 24828 22874
rect 24852 22822 24866 22874
rect 24866 22822 24878 22874
rect 24878 22822 24908 22874
rect 24932 22822 24942 22874
rect 24942 22822 24988 22874
rect 24692 22820 24748 22822
rect 24772 22820 24828 22822
rect 24852 22820 24908 22822
rect 24932 22820 24988 22822
rect 24692 21786 24748 21788
rect 24772 21786 24828 21788
rect 24852 21786 24908 21788
rect 24932 21786 24988 21788
rect 24692 21734 24738 21786
rect 24738 21734 24748 21786
rect 24772 21734 24802 21786
rect 24802 21734 24814 21786
rect 24814 21734 24828 21786
rect 24852 21734 24866 21786
rect 24866 21734 24878 21786
rect 24878 21734 24908 21786
rect 24932 21734 24942 21786
rect 24942 21734 24988 21786
rect 24692 21732 24748 21734
rect 24772 21732 24828 21734
rect 24852 21732 24908 21734
rect 24932 21732 24988 21734
rect 24692 20698 24748 20700
rect 24772 20698 24828 20700
rect 24852 20698 24908 20700
rect 24932 20698 24988 20700
rect 24692 20646 24738 20698
rect 24738 20646 24748 20698
rect 24772 20646 24802 20698
rect 24802 20646 24814 20698
rect 24814 20646 24828 20698
rect 24852 20646 24866 20698
rect 24866 20646 24878 20698
rect 24878 20646 24908 20698
rect 24932 20646 24942 20698
rect 24942 20646 24988 20698
rect 24692 20644 24748 20646
rect 24772 20644 24828 20646
rect 24852 20644 24908 20646
rect 24932 20644 24988 20646
rect 24692 19610 24748 19612
rect 24772 19610 24828 19612
rect 24852 19610 24908 19612
rect 24932 19610 24988 19612
rect 24692 19558 24738 19610
rect 24738 19558 24748 19610
rect 24772 19558 24802 19610
rect 24802 19558 24814 19610
rect 24814 19558 24828 19610
rect 24852 19558 24866 19610
rect 24866 19558 24878 19610
rect 24878 19558 24908 19610
rect 24932 19558 24942 19610
rect 24942 19558 24988 19610
rect 24692 19556 24748 19558
rect 24772 19556 24828 19558
rect 24852 19556 24908 19558
rect 24932 19556 24988 19558
rect 24692 18522 24748 18524
rect 24772 18522 24828 18524
rect 24852 18522 24908 18524
rect 24932 18522 24988 18524
rect 24692 18470 24738 18522
rect 24738 18470 24748 18522
rect 24772 18470 24802 18522
rect 24802 18470 24814 18522
rect 24814 18470 24828 18522
rect 24852 18470 24866 18522
rect 24866 18470 24878 18522
rect 24878 18470 24908 18522
rect 24932 18470 24942 18522
rect 24942 18470 24988 18522
rect 24692 18468 24748 18470
rect 24772 18468 24828 18470
rect 24852 18468 24908 18470
rect 24932 18468 24988 18470
rect 25226 34892 25228 34912
rect 25228 34892 25280 34912
rect 25280 34892 25282 34912
rect 25226 34856 25282 34892
rect 25226 33804 25228 33824
rect 25228 33804 25280 33824
rect 25280 33804 25282 33824
rect 25226 33768 25282 33804
rect 25226 32716 25228 32736
rect 25228 32716 25280 32736
rect 25280 32716 25282 32736
rect 25226 32680 25282 32716
rect 25134 31592 25190 31648
rect 25134 30504 25190 30560
rect 25134 29452 25136 29472
rect 25136 29452 25188 29472
rect 25188 29452 25190 29472
rect 25134 29416 25190 29452
rect 25134 28364 25136 28384
rect 25136 28364 25188 28384
rect 25188 28364 25190 28384
rect 25134 28328 25190 28364
rect 25134 27276 25136 27296
rect 25136 27276 25188 27296
rect 25188 27276 25190 27296
rect 25134 27240 25190 27276
rect 25134 26152 25190 26208
rect 25134 25064 25190 25120
rect 25134 24012 25136 24032
rect 25136 24012 25188 24032
rect 25188 24012 25190 24032
rect 25134 23976 25190 24012
rect 25134 22924 25136 22944
rect 25136 22924 25188 22944
rect 25188 22924 25190 22944
rect 25134 22888 25190 22924
rect 25134 21800 25190 21856
rect 25134 20712 25190 20768
rect 25134 18536 25190 18592
rect 24398 13676 24400 13696
rect 24400 13676 24452 13696
rect 24452 13676 24454 13696
rect 24398 13640 24454 13676
rect 24490 12688 24546 12744
rect 24306 9152 24362 9208
rect 25134 17448 25190 17504
rect 24692 17434 24748 17436
rect 24772 17434 24828 17436
rect 24852 17434 24908 17436
rect 24932 17434 24988 17436
rect 24692 17382 24738 17434
rect 24738 17382 24748 17434
rect 24772 17382 24802 17434
rect 24802 17382 24814 17434
rect 24814 17382 24828 17434
rect 24852 17382 24866 17434
rect 24866 17382 24878 17434
rect 24878 17382 24908 17434
rect 24932 17382 24942 17434
rect 24942 17382 24988 17434
rect 24692 17380 24748 17382
rect 24772 17380 24828 17382
rect 24852 17380 24908 17382
rect 24932 17380 24988 17382
rect 24692 16346 24748 16348
rect 24772 16346 24828 16348
rect 24852 16346 24908 16348
rect 24932 16346 24988 16348
rect 24692 16294 24738 16346
rect 24738 16294 24748 16346
rect 24772 16294 24802 16346
rect 24802 16294 24814 16346
rect 24814 16294 24828 16346
rect 24852 16294 24866 16346
rect 24866 16294 24878 16346
rect 24878 16294 24908 16346
rect 24932 16294 24942 16346
rect 24942 16294 24988 16346
rect 24692 16292 24748 16294
rect 24772 16292 24828 16294
rect 24852 16292 24908 16294
rect 24932 16292 24988 16294
rect 24692 15258 24748 15260
rect 24772 15258 24828 15260
rect 24852 15258 24908 15260
rect 24932 15258 24988 15260
rect 24692 15206 24738 15258
rect 24738 15206 24748 15258
rect 24772 15206 24802 15258
rect 24802 15206 24814 15258
rect 24814 15206 24828 15258
rect 24852 15206 24866 15258
rect 24866 15206 24878 15258
rect 24878 15206 24908 15258
rect 24932 15206 24942 15258
rect 24942 15206 24988 15258
rect 24692 15204 24748 15206
rect 24772 15204 24828 15206
rect 24852 15204 24908 15206
rect 24932 15204 24988 15206
rect 24692 14170 24748 14172
rect 24772 14170 24828 14172
rect 24852 14170 24908 14172
rect 24932 14170 24988 14172
rect 24692 14118 24738 14170
rect 24738 14118 24748 14170
rect 24772 14118 24802 14170
rect 24802 14118 24814 14170
rect 24814 14118 24828 14170
rect 24852 14118 24866 14170
rect 24866 14118 24878 14170
rect 24878 14118 24908 14170
rect 24932 14118 24942 14170
rect 24942 14118 24988 14170
rect 24692 14116 24748 14118
rect 24772 14116 24828 14118
rect 24852 14116 24908 14118
rect 24932 14116 24988 14118
rect 24692 13082 24748 13084
rect 24772 13082 24828 13084
rect 24852 13082 24908 13084
rect 24932 13082 24988 13084
rect 24692 13030 24738 13082
rect 24738 13030 24748 13082
rect 24772 13030 24802 13082
rect 24802 13030 24814 13082
rect 24814 13030 24828 13082
rect 24852 13030 24866 13082
rect 24866 13030 24878 13082
rect 24878 13030 24908 13082
rect 24932 13030 24942 13082
rect 24942 13030 24988 13082
rect 24692 13028 24748 13030
rect 24772 13028 24828 13030
rect 24852 13028 24908 13030
rect 24932 13028 24988 13030
rect 24692 11994 24748 11996
rect 24772 11994 24828 11996
rect 24852 11994 24908 11996
rect 24932 11994 24988 11996
rect 24692 11942 24738 11994
rect 24738 11942 24748 11994
rect 24772 11942 24802 11994
rect 24802 11942 24814 11994
rect 24814 11942 24828 11994
rect 24852 11942 24866 11994
rect 24866 11942 24878 11994
rect 24878 11942 24908 11994
rect 24932 11942 24942 11994
rect 24942 11942 24988 11994
rect 24692 11940 24748 11942
rect 24772 11940 24828 11942
rect 24852 11940 24908 11942
rect 24932 11940 24988 11942
rect 24692 10906 24748 10908
rect 24772 10906 24828 10908
rect 24852 10906 24908 10908
rect 24932 10906 24988 10908
rect 24692 10854 24738 10906
rect 24738 10854 24748 10906
rect 24772 10854 24802 10906
rect 24802 10854 24814 10906
rect 24814 10854 24828 10906
rect 24852 10854 24866 10906
rect 24866 10854 24878 10906
rect 24878 10854 24908 10906
rect 24932 10854 24942 10906
rect 24942 10854 24988 10906
rect 24692 10852 24748 10854
rect 24772 10852 24828 10854
rect 24852 10852 24908 10854
rect 24932 10852 24988 10854
rect 24692 9818 24748 9820
rect 24772 9818 24828 9820
rect 24852 9818 24908 9820
rect 24932 9818 24988 9820
rect 24692 9766 24738 9818
rect 24738 9766 24748 9818
rect 24772 9766 24802 9818
rect 24802 9766 24814 9818
rect 24814 9766 24828 9818
rect 24852 9766 24866 9818
rect 24866 9766 24878 9818
rect 24878 9766 24908 9818
rect 24932 9766 24942 9818
rect 24942 9766 24988 9818
rect 24692 9764 24748 9766
rect 24772 9764 24828 9766
rect 24852 9764 24908 9766
rect 24932 9764 24988 9766
rect 25134 14184 25190 14240
rect 25134 12688 25190 12744
rect 25226 12008 25282 12064
rect 25226 10920 25282 10976
rect 25502 19624 25558 19680
rect 25502 15272 25558 15328
rect 25318 9832 25374 9888
rect 24692 8730 24748 8732
rect 24772 8730 24828 8732
rect 24852 8730 24908 8732
rect 24932 8730 24988 8732
rect 24692 8678 24738 8730
rect 24738 8678 24748 8730
rect 24772 8678 24802 8730
rect 24802 8678 24814 8730
rect 24814 8678 24828 8730
rect 24852 8678 24866 8730
rect 24866 8678 24878 8730
rect 24878 8678 24908 8730
rect 24932 8678 24942 8730
rect 24942 8678 24988 8730
rect 24692 8676 24748 8678
rect 24772 8676 24828 8678
rect 24852 8676 24908 8678
rect 24932 8676 24988 8678
rect 24490 8200 24546 8256
rect 23662 6024 23718 6080
rect 23662 5344 23718 5400
rect 24692 7642 24748 7644
rect 24772 7642 24828 7644
rect 24852 7642 24908 7644
rect 24932 7642 24988 7644
rect 24692 7590 24738 7642
rect 24738 7590 24748 7642
rect 24772 7590 24802 7642
rect 24802 7590 24814 7642
rect 24814 7590 24828 7642
rect 24852 7590 24866 7642
rect 24866 7590 24878 7642
rect 24878 7590 24908 7642
rect 24932 7590 24942 7642
rect 24942 7590 24988 7642
rect 24692 7588 24748 7590
rect 24772 7588 24828 7590
rect 24852 7588 24908 7590
rect 24932 7588 24988 7590
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 25226 7656 25282 7712
rect 25226 4392 25282 4448
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
rect 25686 25200 25742 25256
rect 25686 5752 25742 5808
rect 25686 5480 25742 5536
rect 25686 3168 25742 3224
rect 25870 17176 25926 17232
rect 25594 2352 25650 2408
rect 25686 2216 25742 2272
<< metal3 >>
rect 25840 43618 26000 43648
rect 25086 43558 26000 43618
rect 6880 43552 7196 43553
rect 6880 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7196 43552
rect 6880 43487 7196 43488
rect 12814 43552 13130 43553
rect 12814 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13130 43552
rect 12814 43487 13130 43488
rect 18748 43552 19064 43553
rect 18748 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19064 43552
rect 18748 43487 19064 43488
rect 24682 43552 24998 43553
rect 24682 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 24998 43552
rect 24682 43487 24998 43488
rect 23197 43346 23263 43349
rect 25086 43346 25146 43558
rect 25840 43528 26000 43558
rect 23197 43344 25146 43346
rect 23197 43288 23202 43344
rect 23258 43288 25146 43344
rect 23197 43286 25146 43288
rect 23197 43283 23263 43286
rect 25313 43074 25379 43077
rect 25840 43074 26000 43104
rect 25313 43072 26000 43074
rect 25313 43016 25318 43072
rect 25374 43016 26000 43072
rect 25313 43014 26000 43016
rect 25313 43011 25379 43014
rect 3913 43008 4229 43009
rect 3913 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4229 43008
rect 3913 42943 4229 42944
rect 9847 43008 10163 43009
rect 9847 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10163 43008
rect 9847 42943 10163 42944
rect 15781 43008 16097 43009
rect 15781 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16097 43008
rect 15781 42943 16097 42944
rect 21715 43008 22031 43009
rect 21715 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22031 43008
rect 25840 42984 26000 43014
rect 21715 42943 22031 42944
rect 11697 42938 11763 42941
rect 12249 42940 12315 42941
rect 11830 42938 11836 42940
rect 11697 42936 11836 42938
rect 11697 42880 11702 42936
rect 11758 42880 11836 42936
rect 11697 42878 11836 42880
rect 11697 42875 11763 42878
rect 11830 42876 11836 42878
rect 11900 42876 11906 42940
rect 12198 42938 12204 42940
rect 12158 42878 12204 42938
rect 12268 42936 12315 42940
rect 12310 42880 12315 42936
rect 12198 42876 12204 42878
rect 12268 42876 12315 42880
rect 12249 42875 12315 42876
rect 12525 42940 12591 42941
rect 13813 42940 13879 42941
rect 12525 42936 12572 42940
rect 12636 42938 12642 42940
rect 12525 42880 12530 42936
rect 12525 42876 12572 42880
rect 12636 42878 12682 42938
rect 13813 42936 13860 42940
rect 13924 42938 13930 42940
rect 14273 42938 14339 42941
rect 14917 42940 14983 42941
rect 14406 42938 14412 42940
rect 13813 42880 13818 42936
rect 12636 42876 12642 42878
rect 13813 42876 13860 42880
rect 13924 42878 13970 42938
rect 14273 42936 14412 42938
rect 14273 42880 14278 42936
rect 14334 42880 14412 42936
rect 14273 42878 14412 42880
rect 13924 42876 13930 42878
rect 12525 42875 12591 42876
rect 13813 42875 13879 42876
rect 14273 42875 14339 42878
rect 14406 42876 14412 42878
rect 14476 42876 14482 42940
rect 14917 42936 14964 42940
rect 15028 42938 15034 42940
rect 14917 42880 14922 42936
rect 14917 42876 14964 42880
rect 15028 42878 15074 42938
rect 15028 42876 15034 42878
rect 15510 42876 15516 42940
rect 15580 42938 15586 42940
rect 15653 42938 15719 42941
rect 15580 42936 15719 42938
rect 15580 42880 15658 42936
rect 15714 42880 15719 42936
rect 15580 42878 15719 42880
rect 15580 42876 15586 42878
rect 14917 42875 14983 42876
rect 15653 42875 15719 42878
rect 8385 42802 8451 42805
rect 9397 42802 9463 42805
rect 8385 42800 9463 42802
rect 8385 42744 8390 42800
rect 8446 42744 9402 42800
rect 9458 42744 9463 42800
rect 8385 42742 9463 42744
rect 8385 42739 8451 42742
rect 9397 42739 9463 42742
rect 3049 42666 3115 42669
rect 9121 42666 9187 42669
rect 3049 42664 9187 42666
rect 3049 42608 3054 42664
rect 3110 42608 9126 42664
rect 9182 42608 9187 42664
rect 3049 42606 9187 42608
rect 3049 42603 3115 42606
rect 9121 42603 9187 42606
rect 25129 42530 25195 42533
rect 25840 42530 26000 42560
rect 25129 42528 26000 42530
rect 25129 42472 25134 42528
rect 25190 42472 26000 42528
rect 25129 42470 26000 42472
rect 25129 42467 25195 42470
rect 6880 42464 7196 42465
rect 6880 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7196 42464
rect 6880 42399 7196 42400
rect 12814 42464 13130 42465
rect 12814 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13130 42464
rect 12814 42399 13130 42400
rect 18748 42464 19064 42465
rect 18748 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19064 42464
rect 18748 42399 19064 42400
rect 24682 42464 24998 42465
rect 24682 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 24998 42464
rect 25840 42440 26000 42470
rect 24682 42399 24998 42400
rect 7598 42196 7604 42260
rect 7668 42258 7674 42260
rect 11789 42258 11855 42261
rect 7668 42256 11855 42258
rect 7668 42200 11794 42256
rect 11850 42200 11855 42256
rect 7668 42198 11855 42200
rect 7668 42196 7674 42198
rect 11789 42195 11855 42198
rect 1485 42122 1551 42125
rect 7373 42122 7439 42125
rect 7782 42122 7788 42124
rect 1485 42120 7298 42122
rect 1485 42064 1490 42120
rect 1546 42064 7298 42120
rect 1485 42062 7298 42064
rect 1485 42059 1551 42062
rect 7238 41986 7298 42062
rect 7373 42120 7788 42122
rect 7373 42064 7378 42120
rect 7434 42064 7788 42120
rect 7373 42062 7788 42064
rect 7373 42059 7439 42062
rect 7782 42060 7788 42062
rect 7852 42060 7858 42124
rect 8702 42060 8708 42124
rect 8772 42122 8778 42124
rect 9857 42122 9923 42125
rect 8772 42120 9923 42122
rect 8772 42064 9862 42120
rect 9918 42064 9923 42120
rect 8772 42062 9923 42064
rect 8772 42060 8778 42062
rect 9857 42059 9923 42062
rect 20069 42122 20135 42125
rect 20713 42122 20779 42125
rect 20069 42120 20779 42122
rect 20069 42064 20074 42120
rect 20130 42064 20718 42120
rect 20774 42064 20779 42120
rect 20069 42062 20779 42064
rect 20069 42059 20135 42062
rect 20713 42059 20779 42062
rect 21909 42122 21975 42125
rect 23565 42122 23631 42125
rect 21909 42120 23631 42122
rect 21909 42064 21914 42120
rect 21970 42064 23570 42120
rect 23626 42064 23631 42120
rect 21909 42062 23631 42064
rect 21909 42059 21975 42062
rect 23565 42059 23631 42062
rect 8293 41986 8359 41989
rect 7238 41984 8359 41986
rect 7238 41928 8298 41984
rect 8354 41928 8359 41984
rect 7238 41926 8359 41928
rect 8293 41923 8359 41926
rect 24117 41986 24183 41989
rect 25840 41986 26000 42016
rect 24117 41984 26000 41986
rect 24117 41928 24122 41984
rect 24178 41928 26000 41984
rect 24117 41926 26000 41928
rect 24117 41923 24183 41926
rect 3913 41920 4229 41921
rect 3913 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4229 41920
rect 3913 41855 4229 41856
rect 9847 41920 10163 41921
rect 9847 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10163 41920
rect 9847 41855 10163 41856
rect 15781 41920 16097 41921
rect 15781 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16097 41920
rect 15781 41855 16097 41856
rect 21715 41920 22031 41921
rect 21715 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22031 41920
rect 25840 41896 26000 41926
rect 21715 41855 22031 41856
rect 6177 41850 6243 41853
rect 6310 41850 6316 41852
rect 6177 41848 6316 41850
rect 6177 41792 6182 41848
rect 6238 41792 6316 41848
rect 6177 41790 6316 41792
rect 6177 41787 6243 41790
rect 6310 41788 6316 41790
rect 6380 41788 6386 41852
rect 7649 41850 7715 41853
rect 9397 41852 9463 41853
rect 8150 41850 8156 41852
rect 7649 41848 8156 41850
rect 7649 41792 7654 41848
rect 7710 41792 8156 41848
rect 7649 41790 8156 41792
rect 7649 41787 7715 41790
rect 8150 41788 8156 41790
rect 8220 41788 8226 41852
rect 9397 41848 9444 41852
rect 9508 41850 9514 41852
rect 17309 41850 17375 41853
rect 17534 41850 17540 41852
rect 9397 41792 9402 41848
rect 9397 41788 9444 41792
rect 9508 41790 9554 41850
rect 17309 41848 17540 41850
rect 17309 41792 17314 41848
rect 17370 41792 17540 41848
rect 17309 41790 17540 41792
rect 9508 41788 9514 41790
rect 9397 41787 9463 41788
rect 17309 41787 17375 41790
rect 17534 41788 17540 41790
rect 17604 41788 17610 41852
rect 1158 41652 1164 41716
rect 1228 41714 1234 41716
rect 6545 41714 6611 41717
rect 1228 41712 6611 41714
rect 1228 41656 6550 41712
rect 6606 41656 6611 41712
rect 1228 41654 6611 41656
rect 1228 41652 1234 41654
rect 6545 41651 6611 41654
rect 7925 41714 7991 41717
rect 16389 41716 16455 41717
rect 8518 41714 8524 41716
rect 7925 41712 8524 41714
rect 7925 41656 7930 41712
rect 7986 41656 8524 41712
rect 7925 41654 8524 41656
rect 7925 41651 7991 41654
rect 8518 41652 8524 41654
rect 8588 41652 8594 41716
rect 16389 41712 16436 41716
rect 16500 41714 16506 41716
rect 16389 41656 16394 41712
rect 16389 41652 16436 41656
rect 16500 41654 16546 41714
rect 16500 41652 16506 41654
rect 17350 41652 17356 41716
rect 17420 41714 17426 41716
rect 17585 41714 17651 41717
rect 17420 41712 17651 41714
rect 17420 41656 17590 41712
rect 17646 41656 17651 41712
rect 17420 41654 17651 41656
rect 17420 41652 17426 41654
rect 16389 41651 16455 41652
rect 17585 41651 17651 41654
rect 18413 41716 18479 41717
rect 19425 41716 19491 41717
rect 18413 41712 18460 41716
rect 18524 41714 18530 41716
rect 19374 41714 19380 41716
rect 18413 41656 18418 41712
rect 18413 41652 18460 41656
rect 18524 41654 18570 41714
rect 19334 41654 19380 41714
rect 19444 41712 19491 41716
rect 19486 41656 19491 41712
rect 18524 41652 18530 41654
rect 19374 41652 19380 41654
rect 19444 41652 19491 41656
rect 18413 41651 18479 41652
rect 19425 41651 19491 41652
rect 20345 41714 20411 41717
rect 21357 41714 21423 41717
rect 20345 41712 21423 41714
rect 20345 41656 20350 41712
rect 20406 41656 21362 41712
rect 21418 41656 21423 41712
rect 20345 41654 21423 41656
rect 20345 41651 20411 41654
rect 21357 41651 21423 41654
rect 790 41516 796 41580
rect 860 41578 866 41580
rect 4153 41578 4219 41581
rect 860 41576 4219 41578
rect 860 41520 4158 41576
rect 4214 41520 4219 41576
rect 860 41518 4219 41520
rect 860 41516 866 41518
rect 4153 41515 4219 41518
rect 4613 41580 4679 41581
rect 4613 41576 4660 41580
rect 4724 41578 4730 41580
rect 4613 41520 4618 41576
rect 4613 41516 4660 41520
rect 4724 41518 4770 41578
rect 4724 41516 4730 41518
rect 6126 41516 6132 41580
rect 6196 41578 6202 41580
rect 6729 41578 6795 41581
rect 6196 41576 6795 41578
rect 6196 41520 6734 41576
rect 6790 41520 6795 41576
rect 6196 41518 6795 41520
rect 6196 41516 6202 41518
rect 4613 41515 4679 41516
rect 6729 41515 6795 41518
rect 17769 41578 17835 41581
rect 21633 41578 21699 41581
rect 17769 41576 21699 41578
rect 17769 41520 17774 41576
rect 17830 41520 21638 41576
rect 21694 41520 21699 41576
rect 17769 41518 21699 41520
rect 17769 41515 17835 41518
rect 21633 41515 21699 41518
rect 974 41380 980 41444
rect 1044 41442 1050 41444
rect 3417 41442 3483 41445
rect 1044 41440 3483 41442
rect 1044 41384 3422 41440
rect 3478 41384 3483 41440
rect 1044 41382 3483 41384
rect 1044 41380 1050 41382
rect 3417 41379 3483 41382
rect 18045 41442 18111 41445
rect 18270 41442 18276 41444
rect 18045 41440 18276 41442
rect 18045 41384 18050 41440
rect 18106 41384 18276 41440
rect 18045 41382 18276 41384
rect 18045 41379 18111 41382
rect 18270 41380 18276 41382
rect 18340 41380 18346 41444
rect 25221 41442 25287 41445
rect 25840 41442 26000 41472
rect 25221 41440 26000 41442
rect 25221 41384 25226 41440
rect 25282 41384 26000 41440
rect 25221 41382 26000 41384
rect 25221 41379 25287 41382
rect 6880 41376 7196 41377
rect 6880 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7196 41376
rect 6880 41311 7196 41312
rect 12814 41376 13130 41377
rect 12814 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13130 41376
rect 12814 41311 13130 41312
rect 18748 41376 19064 41377
rect 18748 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19064 41376
rect 18748 41311 19064 41312
rect 24682 41376 24998 41377
rect 24682 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 24998 41376
rect 25840 41352 26000 41382
rect 24682 41311 24998 41312
rect 15101 41170 15167 41173
rect 21725 41170 21791 41173
rect 15101 41168 21791 41170
rect 15101 41112 15106 41168
rect 15162 41112 21730 41168
rect 21786 41112 21791 41168
rect 15101 41110 21791 41112
rect 15101 41107 15167 41110
rect 21725 41107 21791 41110
rect 21541 41034 21607 41037
rect 23749 41034 23815 41037
rect 21541 41032 23815 41034
rect 21541 40976 21546 41032
rect 21602 40976 23754 41032
rect 23810 40976 23815 41032
rect 21541 40974 23815 40976
rect 21541 40971 21607 40974
rect 23749 40971 23815 40974
rect 23657 40898 23723 40901
rect 25840 40898 26000 40928
rect 23657 40896 26000 40898
rect 23657 40840 23662 40896
rect 23718 40840 26000 40896
rect 23657 40838 26000 40840
rect 23657 40835 23723 40838
rect 3913 40832 4229 40833
rect 3913 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4229 40832
rect 3913 40767 4229 40768
rect 9847 40832 10163 40833
rect 9847 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10163 40832
rect 9847 40767 10163 40768
rect 15781 40832 16097 40833
rect 15781 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16097 40832
rect 15781 40767 16097 40768
rect 21715 40832 22031 40833
rect 21715 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22031 40832
rect 25840 40808 26000 40838
rect 21715 40767 22031 40768
rect 5809 40626 5875 40629
rect 14089 40626 14155 40629
rect 22645 40626 22711 40629
rect 5809 40624 22711 40626
rect 5809 40568 5814 40624
rect 5870 40568 14094 40624
rect 14150 40568 22650 40624
rect 22706 40568 22711 40624
rect 5809 40566 22711 40568
rect 5809 40563 5875 40566
rect 14089 40563 14155 40566
rect 22645 40563 22711 40566
rect 3785 40490 3851 40493
rect 6821 40490 6887 40493
rect 3785 40488 6887 40490
rect 3785 40432 3790 40488
rect 3846 40432 6826 40488
rect 6882 40432 6887 40488
rect 3785 40430 6887 40432
rect 3785 40427 3851 40430
rect 6821 40427 6887 40430
rect 20621 40490 20687 40493
rect 22921 40490 22987 40493
rect 20621 40488 22987 40490
rect 20621 40432 20626 40488
rect 20682 40432 22926 40488
rect 22982 40432 22987 40488
rect 20621 40430 22987 40432
rect 20621 40427 20687 40430
rect 22921 40427 22987 40430
rect 20253 40354 20319 40357
rect 23657 40354 23723 40357
rect 20253 40352 23723 40354
rect 20253 40296 20258 40352
rect 20314 40296 23662 40352
rect 23718 40296 23723 40352
rect 20253 40294 23723 40296
rect 20253 40291 20319 40294
rect 23657 40291 23723 40294
rect 25129 40354 25195 40357
rect 25840 40354 26000 40384
rect 25129 40352 26000 40354
rect 25129 40296 25134 40352
rect 25190 40296 26000 40352
rect 25129 40294 26000 40296
rect 25129 40291 25195 40294
rect 6880 40288 7196 40289
rect 6880 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7196 40288
rect 6880 40223 7196 40224
rect 12814 40288 13130 40289
rect 12814 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13130 40288
rect 12814 40223 13130 40224
rect 18748 40288 19064 40289
rect 18748 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19064 40288
rect 18748 40223 19064 40224
rect 24682 40288 24998 40289
rect 24682 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 24998 40288
rect 25840 40264 26000 40294
rect 24682 40223 24998 40224
rect 933 40218 999 40221
rect 4245 40218 4311 40221
rect 933 40216 4311 40218
rect 933 40160 938 40216
rect 994 40160 4250 40216
rect 4306 40160 4311 40216
rect 933 40158 4311 40160
rect 933 40155 999 40158
rect 4245 40155 4311 40158
rect 7465 40218 7531 40221
rect 8937 40218 9003 40221
rect 9121 40218 9187 40221
rect 7465 40216 9187 40218
rect 7465 40160 7470 40216
rect 7526 40160 8942 40216
rect 8998 40160 9126 40216
rect 9182 40160 9187 40216
rect 7465 40158 9187 40160
rect 7465 40155 7531 40158
rect 8937 40155 9003 40158
rect 9121 40155 9187 40158
rect 19701 40218 19767 40221
rect 20805 40218 20871 40221
rect 19701 40216 20871 40218
rect 19701 40160 19706 40216
rect 19762 40160 20810 40216
rect 20866 40160 20871 40216
rect 19701 40158 20871 40160
rect 19701 40155 19767 40158
rect 20805 40155 20871 40158
rect 22870 40156 22876 40220
rect 22940 40218 22946 40220
rect 23013 40218 23079 40221
rect 22940 40216 23079 40218
rect 22940 40160 23018 40216
rect 23074 40160 23079 40216
rect 22940 40158 23079 40160
rect 22940 40156 22946 40158
rect 23013 40155 23079 40158
rect 657 40082 723 40085
rect 3233 40082 3299 40085
rect 657 40080 3299 40082
rect 657 40024 662 40080
rect 718 40024 3238 40080
rect 3294 40024 3299 40080
rect 657 40022 3299 40024
rect 657 40019 723 40022
rect 3233 40019 3299 40022
rect 20069 40082 20135 40085
rect 23105 40082 23171 40085
rect 20069 40080 20362 40082
rect 20069 40024 20074 40080
rect 20130 40024 20362 40080
rect 20069 40022 20362 40024
rect 20069 40019 20135 40022
rect 20302 39946 20362 40022
rect 22050 40080 23171 40082
rect 22050 40024 23110 40080
rect 23166 40024 23171 40080
rect 22050 40022 23171 40024
rect 22050 39946 22110 40022
rect 23105 40019 23171 40022
rect 20302 39886 22110 39946
rect 22277 39946 22343 39949
rect 23197 39946 23263 39949
rect 22277 39944 23263 39946
rect 22277 39888 22282 39944
rect 22338 39888 23202 39944
rect 23258 39888 23263 39944
rect 22277 39886 23263 39888
rect 22277 39883 22343 39886
rect 23197 39883 23263 39886
rect 24393 39810 24459 39813
rect 25840 39810 26000 39840
rect 24393 39808 26000 39810
rect 24393 39752 24398 39808
rect 24454 39752 26000 39808
rect 24393 39750 26000 39752
rect 24393 39747 24459 39750
rect 3913 39744 4229 39745
rect 3913 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4229 39744
rect 3913 39679 4229 39680
rect 9847 39744 10163 39745
rect 9847 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10163 39744
rect 9847 39679 10163 39680
rect 15781 39744 16097 39745
rect 15781 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16097 39744
rect 15781 39679 16097 39680
rect 21715 39744 22031 39745
rect 21715 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22031 39744
rect 25840 39720 26000 39750
rect 21715 39679 22031 39680
rect 0 39538 160 39568
rect 1485 39538 1551 39541
rect 0 39536 1551 39538
rect 0 39480 1490 39536
rect 1546 39480 1551 39536
rect 0 39478 1551 39480
rect 0 39448 160 39478
rect 1485 39475 1551 39478
rect 20805 39538 20871 39541
rect 23013 39538 23079 39541
rect 20805 39536 23079 39538
rect 20805 39480 20810 39536
rect 20866 39480 23018 39536
rect 23074 39480 23079 39536
rect 20805 39478 23079 39480
rect 20805 39475 20871 39478
rect 23013 39475 23079 39478
rect 1393 39400 1459 39405
rect 1393 39344 1398 39400
rect 1454 39344 1459 39400
rect 1393 39339 1459 39344
rect 2221 39402 2287 39405
rect 8661 39402 8727 39405
rect 2221 39400 8727 39402
rect 2221 39344 2226 39400
rect 2282 39344 8666 39400
rect 8722 39344 8727 39400
rect 2221 39342 8727 39344
rect 2221 39339 2287 39342
rect 8661 39339 8727 39342
rect 19977 39402 20043 39405
rect 22829 39402 22895 39405
rect 19977 39400 22895 39402
rect 19977 39344 19982 39400
rect 20038 39344 22834 39400
rect 22890 39344 22895 39400
rect 19977 39342 22895 39344
rect 19977 39339 20043 39342
rect 22829 39339 22895 39342
rect 0 39266 160 39296
rect 1396 39266 1456 39339
rect 0 39206 1456 39266
rect 25221 39266 25287 39269
rect 25840 39266 26000 39296
rect 25221 39264 26000 39266
rect 25221 39208 25226 39264
rect 25282 39208 26000 39264
rect 25221 39206 26000 39208
rect 0 39176 160 39206
rect 25221 39203 25287 39206
rect 6880 39200 7196 39201
rect 6880 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7196 39200
rect 6880 39135 7196 39136
rect 12814 39200 13130 39201
rect 12814 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13130 39200
rect 12814 39135 13130 39136
rect 18748 39200 19064 39201
rect 18748 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19064 39200
rect 18748 39135 19064 39136
rect 24682 39200 24998 39201
rect 24682 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 24998 39200
rect 25840 39176 26000 39206
rect 24682 39135 24998 39136
rect 2630 39068 2636 39132
rect 2700 39130 2706 39132
rect 5257 39130 5323 39133
rect 2700 39128 5323 39130
rect 2700 39072 5262 39128
rect 5318 39072 5323 39128
rect 2700 39070 5323 39072
rect 2700 39068 2706 39070
rect 5257 39067 5323 39070
rect 0 38994 160 39024
rect 2773 38994 2839 38997
rect 0 38992 2839 38994
rect 0 38936 2778 38992
rect 2834 38936 2839 38992
rect 0 38934 2839 38936
rect 0 38904 160 38934
rect 2773 38931 2839 38934
rect 16849 38994 16915 38997
rect 22502 38994 22508 38996
rect 16849 38992 22508 38994
rect 16849 38936 16854 38992
rect 16910 38936 22508 38992
rect 16849 38934 22508 38936
rect 16849 38931 16915 38934
rect 22502 38932 22508 38934
rect 22572 38932 22578 38996
rect 3877 38858 3943 38861
rect 2730 38856 3943 38858
rect 2730 38800 3882 38856
rect 3938 38800 3943 38856
rect 2730 38798 3943 38800
rect 0 38722 160 38752
rect 2730 38722 2790 38798
rect 3877 38795 3943 38798
rect 20437 38858 20503 38861
rect 21817 38858 21883 38861
rect 20437 38856 21883 38858
rect 20437 38800 20442 38856
rect 20498 38800 21822 38856
rect 21878 38800 21883 38856
rect 20437 38798 21883 38800
rect 20437 38795 20503 38798
rect 21817 38795 21883 38798
rect 0 38662 2790 38722
rect 4705 38722 4771 38725
rect 9622 38722 9628 38724
rect 4705 38720 9628 38722
rect 4705 38664 4710 38720
rect 4766 38664 9628 38720
rect 4705 38662 9628 38664
rect 0 38632 160 38662
rect 4705 38659 4771 38662
rect 9622 38660 9628 38662
rect 9692 38660 9698 38724
rect 18505 38722 18571 38725
rect 19558 38722 19564 38724
rect 18505 38720 19564 38722
rect 18505 38664 18510 38720
rect 18566 38664 19564 38720
rect 18505 38662 19564 38664
rect 18505 38659 18571 38662
rect 19558 38660 19564 38662
rect 19628 38660 19634 38724
rect 24393 38722 24459 38725
rect 25840 38722 26000 38752
rect 24393 38720 26000 38722
rect 24393 38664 24398 38720
rect 24454 38664 26000 38720
rect 24393 38662 26000 38664
rect 24393 38659 24459 38662
rect 3913 38656 4229 38657
rect 3913 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4229 38656
rect 3913 38591 4229 38592
rect 9847 38656 10163 38657
rect 9847 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10163 38656
rect 9847 38591 10163 38592
rect 15781 38656 16097 38657
rect 15781 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16097 38656
rect 15781 38591 16097 38592
rect 21715 38656 22031 38657
rect 21715 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22031 38656
rect 25840 38632 26000 38662
rect 21715 38591 22031 38592
rect 0 38450 160 38480
rect 3049 38450 3115 38453
rect 0 38448 3115 38450
rect 0 38392 3054 38448
rect 3110 38392 3115 38448
rect 0 38390 3115 38392
rect 0 38360 160 38390
rect 3049 38387 3115 38390
rect 2221 38314 2287 38317
rect 5625 38314 5691 38317
rect 2221 38312 5691 38314
rect 2221 38256 2226 38312
rect 2282 38256 5630 38312
rect 5686 38256 5691 38312
rect 2221 38254 5691 38256
rect 2221 38251 2287 38254
rect 5625 38251 5691 38254
rect 0 38178 160 38208
rect 1209 38178 1275 38181
rect 0 38176 1275 38178
rect 0 38120 1214 38176
rect 1270 38120 1275 38176
rect 0 38118 1275 38120
rect 0 38088 160 38118
rect 1209 38115 1275 38118
rect 2814 38116 2820 38180
rect 2884 38178 2890 38180
rect 3049 38178 3115 38181
rect 2884 38176 3115 38178
rect 2884 38120 3054 38176
rect 3110 38120 3115 38176
rect 2884 38118 3115 38120
rect 2884 38116 2890 38118
rect 3049 38115 3115 38118
rect 25221 38178 25287 38181
rect 25840 38178 26000 38208
rect 25221 38176 26000 38178
rect 25221 38120 25226 38176
rect 25282 38120 26000 38176
rect 25221 38118 26000 38120
rect 25221 38115 25287 38118
rect 6880 38112 7196 38113
rect 6880 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7196 38112
rect 6880 38047 7196 38048
rect 12814 38112 13130 38113
rect 12814 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13130 38112
rect 12814 38047 13130 38048
rect 18748 38112 19064 38113
rect 18748 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19064 38112
rect 18748 38047 19064 38048
rect 24682 38112 24998 38113
rect 24682 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 24998 38112
rect 25840 38088 26000 38118
rect 24682 38047 24998 38048
rect 3417 38042 3483 38045
rect 1396 38040 3483 38042
rect 1396 37984 3422 38040
rect 3478 37984 3483 38040
rect 1396 37982 3483 37984
rect 0 37906 160 37936
rect 749 37906 815 37909
rect 0 37904 815 37906
rect 0 37848 754 37904
rect 810 37848 815 37904
rect 0 37846 815 37848
rect 0 37816 160 37846
rect 749 37843 815 37846
rect 0 37634 160 37664
rect 1396 37634 1456 37982
rect 3417 37979 3483 37982
rect 1669 37906 1735 37909
rect 5809 37906 5875 37909
rect 17902 37906 17908 37908
rect 1669 37904 5642 37906
rect 1669 37848 1674 37904
rect 1730 37848 5642 37904
rect 1669 37846 5642 37848
rect 1669 37843 1735 37846
rect 5582 37770 5642 37846
rect 5809 37904 17908 37906
rect 5809 37848 5814 37904
rect 5870 37848 17908 37904
rect 5809 37846 17908 37848
rect 5809 37843 5875 37846
rect 17902 37844 17908 37846
rect 17972 37844 17978 37908
rect 11094 37770 11100 37772
rect 5582 37710 11100 37770
rect 11094 37708 11100 37710
rect 11164 37708 11170 37772
rect 0 37574 1456 37634
rect 24393 37634 24459 37637
rect 25840 37634 26000 37664
rect 24393 37632 26000 37634
rect 24393 37576 24398 37632
rect 24454 37576 26000 37632
rect 24393 37574 26000 37576
rect 0 37544 160 37574
rect 24393 37571 24459 37574
rect 3913 37568 4229 37569
rect 3913 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4229 37568
rect 3913 37503 4229 37504
rect 9847 37568 10163 37569
rect 9847 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10163 37568
rect 9847 37503 10163 37504
rect 15781 37568 16097 37569
rect 15781 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16097 37568
rect 15781 37503 16097 37504
rect 21715 37568 22031 37569
rect 21715 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22031 37568
rect 25840 37544 26000 37574
rect 21715 37503 22031 37504
rect 2957 37500 3023 37501
rect 2957 37496 3004 37500
rect 3068 37498 3074 37500
rect 2957 37440 2962 37496
rect 2957 37436 3004 37440
rect 3068 37438 3114 37498
rect 3068 37436 3074 37438
rect 2957 37435 3023 37436
rect 0 37362 160 37392
rect 4889 37362 4955 37365
rect 0 37360 4955 37362
rect 0 37304 4894 37360
rect 4950 37304 4955 37360
rect 0 37302 4955 37304
rect 0 37272 160 37302
rect 4889 37299 4955 37302
rect 5533 37362 5599 37365
rect 6678 37362 6684 37364
rect 5533 37360 6684 37362
rect 5533 37304 5538 37360
rect 5594 37304 6684 37360
rect 5533 37302 6684 37304
rect 5533 37299 5599 37302
rect 6678 37300 6684 37302
rect 6748 37300 6754 37364
rect 8201 37362 8267 37365
rect 8886 37362 8892 37364
rect 8201 37360 8892 37362
rect 8201 37304 8206 37360
rect 8262 37304 8892 37360
rect 8201 37302 8892 37304
rect 8201 37299 8267 37302
rect 8886 37300 8892 37302
rect 8956 37300 8962 37364
rect 2773 37226 2839 37229
rect 12341 37226 12407 37229
rect 2773 37224 12407 37226
rect 2773 37168 2778 37224
rect 2834 37168 12346 37224
rect 12402 37168 12407 37224
rect 2773 37166 12407 37168
rect 2773 37163 2839 37166
rect 12341 37163 12407 37166
rect 24117 37226 24183 37229
rect 24117 37224 25146 37226
rect 24117 37168 24122 37224
rect 24178 37168 25146 37224
rect 24117 37166 25146 37168
rect 24117 37163 24183 37166
rect 0 37090 160 37120
rect 3877 37090 3943 37093
rect 0 37088 3943 37090
rect 0 37032 3882 37088
rect 3938 37032 3943 37088
rect 0 37030 3943 37032
rect 25086 37090 25146 37166
rect 25840 37090 26000 37120
rect 25086 37030 26000 37090
rect 0 37000 160 37030
rect 3877 37027 3943 37030
rect 6880 37024 7196 37025
rect 6880 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7196 37024
rect 6880 36959 7196 36960
rect 12814 37024 13130 37025
rect 12814 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13130 37024
rect 12814 36959 13130 36960
rect 18748 37024 19064 37025
rect 18748 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19064 37024
rect 18748 36959 19064 36960
rect 24682 37024 24998 37025
rect 24682 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 24998 37024
rect 25840 37000 26000 37030
rect 24682 36959 24998 36960
rect 289 36954 355 36957
rect 4337 36954 4403 36957
rect 289 36952 4403 36954
rect 289 36896 294 36952
rect 350 36896 4342 36952
rect 4398 36896 4403 36952
rect 289 36894 4403 36896
rect 289 36891 355 36894
rect 4337 36891 4403 36894
rect 0 36818 160 36848
rect 3141 36818 3207 36821
rect 0 36816 3207 36818
rect 0 36760 3146 36816
rect 3202 36760 3207 36816
rect 0 36758 3207 36760
rect 0 36728 160 36758
rect 3141 36755 3207 36758
rect 4061 36818 4127 36821
rect 7741 36818 7807 36821
rect 4061 36816 7807 36818
rect 4061 36760 4066 36816
rect 4122 36760 7746 36816
rect 7802 36760 7807 36816
rect 4061 36758 7807 36760
rect 4061 36755 4127 36758
rect 7741 36755 7807 36758
rect 1761 36682 1827 36685
rect 15561 36682 15627 36685
rect 1761 36680 15627 36682
rect 1761 36624 1766 36680
rect 1822 36624 15566 36680
rect 15622 36624 15627 36680
rect 1761 36622 15627 36624
rect 1761 36619 1827 36622
rect 15561 36619 15627 36622
rect 0 36546 160 36576
rect 1945 36546 2011 36549
rect 0 36544 2011 36546
rect 0 36488 1950 36544
rect 2006 36488 2011 36544
rect 0 36486 2011 36488
rect 0 36456 160 36486
rect 1945 36483 2011 36486
rect 2313 36546 2379 36549
rect 3785 36546 3851 36549
rect 2313 36544 3851 36546
rect 2313 36488 2318 36544
rect 2374 36488 3790 36544
rect 3846 36488 3851 36544
rect 2313 36486 3851 36488
rect 2313 36483 2379 36486
rect 3785 36483 3851 36486
rect 24393 36546 24459 36549
rect 25840 36546 26000 36576
rect 24393 36544 26000 36546
rect 24393 36488 24398 36544
rect 24454 36488 26000 36544
rect 24393 36486 26000 36488
rect 24393 36483 24459 36486
rect 3913 36480 4229 36481
rect 3913 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4229 36480
rect 3913 36415 4229 36416
rect 9847 36480 10163 36481
rect 9847 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10163 36480
rect 9847 36415 10163 36416
rect 15781 36480 16097 36481
rect 15781 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16097 36480
rect 15781 36415 16097 36416
rect 21715 36480 22031 36481
rect 21715 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22031 36480
rect 25840 36456 26000 36486
rect 21715 36415 22031 36416
rect 0 36274 160 36304
rect 1669 36274 1735 36277
rect 0 36272 1735 36274
rect 0 36216 1674 36272
rect 1730 36216 1735 36272
rect 0 36214 1735 36216
rect 0 36184 160 36214
rect 1669 36211 1735 36214
rect 2221 36138 2287 36141
rect 2446 36138 2452 36140
rect 2221 36136 2452 36138
rect 2221 36080 2226 36136
rect 2282 36080 2452 36136
rect 2221 36078 2452 36080
rect 2221 36075 2287 36078
rect 2446 36076 2452 36078
rect 2516 36076 2522 36140
rect 2998 36076 3004 36140
rect 3068 36138 3074 36140
rect 7373 36138 7439 36141
rect 3068 36136 7439 36138
rect 3068 36080 7378 36136
rect 7434 36080 7439 36136
rect 3068 36078 7439 36080
rect 3068 36076 3074 36078
rect 7373 36075 7439 36078
rect 8937 36138 9003 36141
rect 9397 36138 9463 36141
rect 8937 36136 9463 36138
rect 8937 36080 8942 36136
rect 8998 36080 9402 36136
rect 9458 36080 9463 36136
rect 8937 36078 9463 36080
rect 8937 36075 9003 36078
rect 9397 36075 9463 36078
rect 0 36002 160 36032
rect 3601 36002 3667 36005
rect 0 36000 3667 36002
rect 0 35944 3606 36000
rect 3662 35944 3667 36000
rect 0 35942 3667 35944
rect 0 35912 160 35942
rect 3601 35939 3667 35942
rect 3734 35940 3740 36004
rect 3804 36002 3810 36004
rect 4061 36002 4127 36005
rect 3804 36000 4127 36002
rect 3804 35944 4066 36000
rect 4122 35944 4127 36000
rect 3804 35942 4127 35944
rect 3804 35940 3810 35942
rect 4061 35939 4127 35942
rect 22737 36002 22803 36005
rect 22870 36002 22876 36004
rect 22737 36000 22876 36002
rect 22737 35944 22742 36000
rect 22798 35944 22876 36000
rect 22737 35942 22876 35944
rect 22737 35939 22803 35942
rect 22870 35940 22876 35942
rect 22940 35940 22946 36004
rect 25129 36002 25195 36005
rect 25840 36002 26000 36032
rect 25129 36000 26000 36002
rect 25129 35944 25134 36000
rect 25190 35944 26000 36000
rect 25129 35942 26000 35944
rect 25129 35939 25195 35942
rect 6880 35936 7196 35937
rect 6880 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7196 35936
rect 6880 35871 7196 35872
rect 12814 35936 13130 35937
rect 12814 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13130 35936
rect 12814 35871 13130 35872
rect 18748 35936 19064 35937
rect 18748 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19064 35936
rect 18748 35871 19064 35872
rect 24682 35936 24998 35937
rect 24682 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 24998 35936
rect 25840 35912 26000 35942
rect 24682 35871 24998 35872
rect 10409 35866 10475 35869
rect 10542 35866 10548 35868
rect 10409 35864 10548 35866
rect 10409 35808 10414 35864
rect 10470 35808 10548 35864
rect 10409 35806 10548 35808
rect 10409 35803 10475 35806
rect 10542 35804 10548 35806
rect 10612 35804 10618 35868
rect 0 35730 160 35760
rect 2773 35730 2839 35733
rect 0 35728 2839 35730
rect 0 35672 2778 35728
rect 2834 35672 2839 35728
rect 0 35670 2839 35672
rect 0 35640 160 35670
rect 2773 35667 2839 35670
rect 5625 35594 5691 35597
rect 11789 35594 11855 35597
rect 18873 35594 18939 35597
rect 5625 35592 10472 35594
rect 5625 35536 5630 35592
rect 5686 35536 10472 35592
rect 5625 35534 10472 35536
rect 5625 35531 5691 35534
rect 0 35458 160 35488
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35368 160 35398
rect 1577 35395 1643 35398
rect 6678 35396 6684 35460
rect 6748 35458 6754 35460
rect 8753 35458 8819 35461
rect 6748 35456 8819 35458
rect 6748 35400 8758 35456
rect 8814 35400 8819 35456
rect 6748 35398 8819 35400
rect 6748 35396 6754 35398
rect 8753 35395 8819 35398
rect 3913 35392 4229 35393
rect 3913 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4229 35392
rect 3913 35327 4229 35328
rect 9847 35392 10163 35393
rect 9847 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10163 35392
rect 9847 35327 10163 35328
rect 10412 35325 10472 35534
rect 11789 35592 18939 35594
rect 11789 35536 11794 35592
rect 11850 35536 18878 35592
rect 18934 35536 18939 35592
rect 11789 35534 18939 35536
rect 11789 35531 11855 35534
rect 18873 35531 18939 35534
rect 13537 35458 13603 35461
rect 11470 35456 13603 35458
rect 11470 35400 13542 35456
rect 13598 35400 13603 35456
rect 11470 35398 13603 35400
rect 10409 35322 10475 35325
rect 11470 35324 11530 35398
rect 13537 35395 13603 35398
rect 24393 35458 24459 35461
rect 25840 35458 26000 35488
rect 24393 35456 26000 35458
rect 24393 35400 24398 35456
rect 24454 35400 26000 35456
rect 24393 35398 26000 35400
rect 24393 35395 24459 35398
rect 15781 35392 16097 35393
rect 15781 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16097 35392
rect 15781 35327 16097 35328
rect 21715 35392 22031 35393
rect 21715 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22031 35392
rect 25840 35368 26000 35398
rect 21715 35327 22031 35328
rect 11462 35322 11468 35324
rect 10409 35320 11468 35322
rect 10409 35264 10414 35320
rect 10470 35264 11468 35320
rect 10409 35262 11468 35264
rect 10409 35259 10475 35262
rect 11462 35260 11468 35262
rect 11532 35260 11538 35324
rect 11605 35322 11671 35325
rect 14365 35322 14431 35325
rect 11605 35320 14431 35322
rect 11605 35264 11610 35320
rect 11666 35264 14370 35320
rect 14426 35264 14431 35320
rect 11605 35262 14431 35264
rect 11605 35259 11671 35262
rect 14365 35259 14431 35262
rect 0 35186 160 35216
rect 3785 35186 3851 35189
rect 0 35184 3851 35186
rect 0 35128 3790 35184
rect 3846 35128 3851 35184
rect 0 35126 3851 35128
rect 0 35096 160 35126
rect 3785 35123 3851 35126
rect 5441 35186 5507 35189
rect 5574 35186 5580 35188
rect 5441 35184 5580 35186
rect 5441 35128 5446 35184
rect 5502 35128 5580 35184
rect 5441 35126 5580 35128
rect 5441 35123 5507 35126
rect 5574 35124 5580 35126
rect 5644 35124 5650 35188
rect 10041 35186 10107 35189
rect 13169 35186 13235 35189
rect 9630 35184 13235 35186
rect 9630 35128 10046 35184
rect 10102 35128 13174 35184
rect 13230 35128 13235 35184
rect 9630 35126 13235 35128
rect 5901 35050 5967 35053
rect 9630 35050 9690 35126
rect 10041 35123 10107 35126
rect 13169 35123 13235 35126
rect 5901 35048 9690 35050
rect 5901 34992 5906 35048
rect 5962 34992 9690 35048
rect 5901 34990 9690 34992
rect 12985 35050 13051 35053
rect 13302 35050 13308 35052
rect 12985 35048 13308 35050
rect 12985 34992 12990 35048
rect 13046 34992 13308 35048
rect 12985 34990 13308 34992
rect 5901 34987 5967 34990
rect 12985 34987 13051 34990
rect 13302 34988 13308 34990
rect 13372 34988 13378 35052
rect 0 34914 160 34944
rect 1393 34914 1459 34917
rect 0 34912 1459 34914
rect 0 34856 1398 34912
rect 1454 34856 1459 34912
rect 0 34854 1459 34856
rect 0 34824 160 34854
rect 1393 34851 1459 34854
rect 4245 34914 4311 34917
rect 4981 34914 5047 34917
rect 4245 34912 5047 34914
rect 4245 34856 4250 34912
rect 4306 34856 4986 34912
rect 5042 34856 5047 34912
rect 4245 34854 5047 34856
rect 4245 34851 4311 34854
rect 4981 34851 5047 34854
rect 7833 34914 7899 34917
rect 9213 34914 9279 34917
rect 7833 34912 9279 34914
rect 7833 34856 7838 34912
rect 7894 34856 9218 34912
rect 9274 34856 9279 34912
rect 7833 34854 9279 34856
rect 7833 34851 7899 34854
rect 9213 34851 9279 34854
rect 9581 34914 9647 34917
rect 11789 34914 11855 34917
rect 12341 34914 12407 34917
rect 9581 34912 9690 34914
rect 9581 34856 9586 34912
rect 9642 34856 9690 34912
rect 9581 34851 9690 34856
rect 11789 34912 12407 34914
rect 11789 34856 11794 34912
rect 11850 34856 12346 34912
rect 12402 34856 12407 34912
rect 11789 34854 12407 34856
rect 11789 34851 11855 34854
rect 12341 34851 12407 34854
rect 25221 34914 25287 34917
rect 25840 34914 26000 34944
rect 25221 34912 26000 34914
rect 25221 34856 25226 34912
rect 25282 34856 26000 34912
rect 25221 34854 26000 34856
rect 25221 34851 25287 34854
rect 6880 34848 7196 34849
rect 6880 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7196 34848
rect 6880 34783 7196 34784
rect 9630 34778 9690 34851
rect 12814 34848 13130 34849
rect 12814 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13130 34848
rect 12814 34783 13130 34784
rect 18748 34848 19064 34849
rect 18748 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19064 34848
rect 18748 34783 19064 34784
rect 24682 34848 24998 34849
rect 24682 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 24998 34848
rect 25840 34824 26000 34854
rect 24682 34783 24998 34784
rect 9630 34718 12450 34778
rect 0 34642 160 34672
rect 749 34642 815 34645
rect 2037 34644 2103 34645
rect 2037 34642 2084 34644
rect 0 34640 815 34642
rect 0 34584 754 34640
rect 810 34584 815 34640
rect 0 34582 815 34584
rect 1992 34640 2084 34642
rect 1992 34584 2042 34640
rect 1992 34582 2084 34584
rect 0 34552 160 34582
rect 749 34579 815 34582
rect 2037 34580 2084 34582
rect 2148 34580 2154 34644
rect 4470 34580 4476 34644
rect 4540 34642 4546 34644
rect 5073 34642 5139 34645
rect 8293 34642 8359 34645
rect 9029 34642 9095 34645
rect 10685 34642 10751 34645
rect 4540 34640 8954 34642
rect 4540 34584 5078 34640
rect 5134 34584 8298 34640
rect 8354 34584 8954 34640
rect 4540 34582 8954 34584
rect 4540 34580 4546 34582
rect 2037 34579 2103 34580
rect 5073 34579 5139 34582
rect 8293 34579 8359 34582
rect 4061 34506 4127 34509
rect 2730 34504 4127 34506
rect 2730 34448 4066 34504
rect 4122 34448 4127 34504
rect 2730 34446 4127 34448
rect 0 34370 160 34400
rect 2730 34370 2790 34446
rect 4061 34443 4127 34446
rect 5390 34444 5396 34508
rect 5460 34506 5466 34508
rect 5533 34506 5599 34509
rect 5460 34504 5599 34506
rect 5460 34448 5538 34504
rect 5594 34448 5599 34504
rect 5460 34446 5599 34448
rect 8894 34506 8954 34582
rect 9029 34640 10751 34642
rect 9029 34584 9034 34640
rect 9090 34584 10690 34640
rect 10746 34584 10751 34640
rect 9029 34582 10751 34584
rect 12390 34642 12450 34718
rect 13261 34642 13327 34645
rect 12390 34640 13327 34642
rect 12390 34584 13266 34640
rect 13322 34584 13327 34640
rect 12390 34582 13327 34584
rect 9029 34579 9095 34582
rect 10685 34579 10751 34582
rect 13261 34579 13327 34582
rect 11605 34506 11671 34509
rect 8894 34504 11671 34506
rect 8894 34448 11610 34504
rect 11666 34448 11671 34504
rect 8894 34446 11671 34448
rect 5460 34444 5466 34446
rect 5533 34443 5599 34446
rect 11605 34443 11671 34446
rect 24393 34506 24459 34509
rect 24393 34504 25146 34506
rect 24393 34448 24398 34504
rect 24454 34448 25146 34504
rect 24393 34446 25146 34448
rect 24393 34443 24459 34446
rect 0 34310 2790 34370
rect 9121 34370 9187 34373
rect 9489 34370 9555 34373
rect 9121 34368 9555 34370
rect 9121 34312 9126 34368
rect 9182 34312 9494 34368
rect 9550 34312 9555 34368
rect 9121 34310 9555 34312
rect 25086 34370 25146 34446
rect 25840 34370 26000 34400
rect 25086 34310 26000 34370
rect 0 34280 160 34310
rect 9121 34307 9187 34310
rect 9489 34307 9555 34310
rect 3913 34304 4229 34305
rect 3913 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4229 34304
rect 3913 34239 4229 34240
rect 9847 34304 10163 34305
rect 9847 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10163 34304
rect 9847 34239 10163 34240
rect 15781 34304 16097 34305
rect 15781 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16097 34304
rect 15781 34239 16097 34240
rect 21715 34304 22031 34305
rect 21715 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22031 34304
rect 25840 34280 26000 34310
rect 21715 34239 22031 34240
rect 0 34098 160 34128
rect 3417 34098 3483 34101
rect 0 34096 3483 34098
rect 0 34040 3422 34096
rect 3478 34040 3483 34096
rect 0 34038 3483 34040
rect 0 34008 160 34038
rect 3417 34035 3483 34038
rect 3601 34098 3667 34101
rect 4654 34098 4660 34100
rect 3601 34096 4660 34098
rect 3601 34040 3606 34096
rect 3662 34040 4660 34096
rect 3601 34038 4660 34040
rect 3601 34035 3667 34038
rect 4654 34036 4660 34038
rect 4724 34036 4730 34100
rect 8753 34098 8819 34101
rect 11697 34098 11763 34101
rect 8753 34096 11763 34098
rect 8753 34040 8758 34096
rect 8814 34040 11702 34096
rect 11758 34040 11763 34096
rect 8753 34038 11763 34040
rect 8753 34035 8819 34038
rect 11697 34035 11763 34038
rect 2681 33962 2747 33965
rect 1396 33960 2747 33962
rect 1396 33904 2686 33960
rect 2742 33904 2747 33960
rect 1396 33902 2747 33904
rect 0 33826 160 33856
rect 1396 33826 1456 33902
rect 2681 33899 2747 33902
rect 6177 33962 6243 33965
rect 8937 33962 9003 33965
rect 11237 33962 11303 33965
rect 6177 33960 11303 33962
rect 6177 33904 6182 33960
rect 6238 33904 8942 33960
rect 8998 33904 11242 33960
rect 11298 33904 11303 33960
rect 6177 33902 11303 33904
rect 6177 33899 6243 33902
rect 8937 33899 9003 33902
rect 11237 33899 11303 33902
rect 0 33766 1456 33826
rect 2681 33826 2747 33829
rect 2998 33826 3004 33828
rect 2681 33824 3004 33826
rect 2681 33768 2686 33824
rect 2742 33768 3004 33824
rect 2681 33766 3004 33768
rect 0 33736 160 33766
rect 2681 33763 2747 33766
rect 2998 33764 3004 33766
rect 3068 33764 3074 33828
rect 25221 33826 25287 33829
rect 25840 33826 26000 33856
rect 25221 33824 26000 33826
rect 25221 33768 25226 33824
rect 25282 33768 26000 33824
rect 25221 33766 26000 33768
rect 25221 33763 25287 33766
rect 6880 33760 7196 33761
rect 6880 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7196 33760
rect 6880 33695 7196 33696
rect 12814 33760 13130 33761
rect 12814 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13130 33760
rect 12814 33695 13130 33696
rect 18748 33760 19064 33761
rect 18748 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19064 33760
rect 18748 33695 19064 33696
rect 24682 33760 24998 33761
rect 24682 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 24998 33760
rect 25840 33736 26000 33766
rect 24682 33695 24998 33696
rect 3734 33628 3740 33692
rect 3804 33690 3810 33692
rect 4337 33690 4403 33693
rect 7833 33690 7899 33693
rect 8109 33690 8175 33693
rect 3804 33688 6792 33690
rect 3804 33632 4342 33688
rect 4398 33632 6792 33688
rect 3804 33630 6792 33632
rect 3804 33628 3810 33630
rect 4337 33627 4403 33630
rect 0 33554 160 33584
rect 1209 33554 1275 33557
rect 0 33552 1275 33554
rect 0 33496 1214 33552
rect 1270 33496 1275 33552
rect 0 33494 1275 33496
rect 6732 33554 6792 33630
rect 7833 33688 8175 33690
rect 7833 33632 7838 33688
rect 7894 33632 8114 33688
rect 8170 33632 8175 33688
rect 7833 33630 8175 33632
rect 7833 33627 7899 33630
rect 8109 33627 8175 33630
rect 10910 33554 10916 33556
rect 6732 33494 10916 33554
rect 0 33464 160 33494
rect 1209 33491 1275 33494
rect 10910 33492 10916 33494
rect 10980 33554 10986 33556
rect 13721 33554 13787 33557
rect 10980 33552 13787 33554
rect 10980 33496 13726 33552
rect 13782 33496 13787 33552
rect 10980 33494 13787 33496
rect 10980 33492 10986 33494
rect 13721 33491 13787 33494
rect 18873 33554 18939 33557
rect 22369 33554 22435 33557
rect 18873 33552 22435 33554
rect 18873 33496 18878 33552
rect 18934 33496 22374 33552
rect 22430 33496 22435 33552
rect 18873 33494 22435 33496
rect 18873 33491 18939 33494
rect 22369 33491 22435 33494
rect 2446 33356 2452 33420
rect 2516 33418 2522 33420
rect 6913 33418 6979 33421
rect 2516 33416 6979 33418
rect 2516 33360 6918 33416
rect 6974 33360 6979 33416
rect 2516 33358 6979 33360
rect 2516 33356 2522 33358
rect 6913 33355 6979 33358
rect 7189 33418 7255 33421
rect 9857 33418 9923 33421
rect 7189 33416 9923 33418
rect 7189 33360 7194 33416
rect 7250 33360 9862 33416
rect 9918 33360 9923 33416
rect 7189 33358 9923 33360
rect 7189 33355 7255 33358
rect 9857 33355 9923 33358
rect 12617 33418 12683 33421
rect 12617 33416 19810 33418
rect 12617 33360 12622 33416
rect 12678 33360 19810 33416
rect 12617 33358 19810 33360
rect 12617 33355 12683 33358
rect 0 33282 160 33312
rect 2865 33282 2931 33285
rect 0 33280 2931 33282
rect 0 33224 2870 33280
rect 2926 33224 2931 33280
rect 0 33222 2931 33224
rect 0 33192 160 33222
rect 2865 33219 2931 33222
rect 6269 33282 6335 33285
rect 9397 33282 9463 33285
rect 6269 33280 9463 33282
rect 6269 33224 6274 33280
rect 6330 33224 9402 33280
rect 9458 33224 9463 33280
rect 6269 33222 9463 33224
rect 6269 33219 6335 33222
rect 9397 33219 9463 33222
rect 12525 33282 12591 33285
rect 15469 33282 15535 33285
rect 19750 33284 19810 33358
rect 19926 33356 19932 33420
rect 19996 33418 20002 33420
rect 22553 33418 22619 33421
rect 19996 33416 22619 33418
rect 19996 33360 22558 33416
rect 22614 33360 22619 33416
rect 19996 33358 22619 33360
rect 19996 33356 20002 33358
rect 22553 33355 22619 33358
rect 12525 33280 15535 33282
rect 12525 33224 12530 33280
rect 12586 33224 15474 33280
rect 15530 33224 15535 33280
rect 12525 33222 15535 33224
rect 12525 33219 12591 33222
rect 15469 33219 15535 33222
rect 19742 33220 19748 33284
rect 19812 33220 19818 33284
rect 24393 33282 24459 33285
rect 25840 33282 26000 33312
rect 24393 33280 26000 33282
rect 24393 33224 24398 33280
rect 24454 33224 26000 33280
rect 24393 33222 26000 33224
rect 24393 33219 24459 33222
rect 3913 33216 4229 33217
rect 3913 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4229 33216
rect 3913 33151 4229 33152
rect 9847 33216 10163 33217
rect 9847 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10163 33216
rect 9847 33151 10163 33152
rect 15781 33216 16097 33217
rect 15781 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16097 33216
rect 15781 33151 16097 33152
rect 21715 33216 22031 33217
rect 21715 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22031 33216
rect 25840 33192 26000 33222
rect 21715 33151 22031 33152
rect 0 33010 160 33040
rect 1485 33010 1551 33013
rect 0 33008 1551 33010
rect 0 32952 1490 33008
rect 1546 32952 1551 33008
rect 0 32950 1551 32952
rect 0 32920 160 32950
rect 1485 32947 1551 32950
rect 9622 32948 9628 33012
rect 9692 33010 9698 33012
rect 11237 33010 11303 33013
rect 9692 33008 11303 33010
rect 9692 32952 11242 33008
rect 11298 32952 11303 33008
rect 9692 32950 11303 32952
rect 9692 32948 9698 32950
rect 11237 32947 11303 32950
rect 1669 32874 1735 32877
rect 10358 32874 10364 32876
rect 1669 32872 10364 32874
rect 1669 32816 1674 32872
rect 1730 32816 10364 32872
rect 1669 32814 10364 32816
rect 1669 32811 1735 32814
rect 10358 32812 10364 32814
rect 10428 32812 10434 32876
rect 12157 32874 12223 32877
rect 16021 32874 16087 32877
rect 12157 32872 16087 32874
rect 12157 32816 12162 32872
rect 12218 32816 16026 32872
rect 16082 32816 16087 32872
rect 12157 32814 16087 32816
rect 12157 32811 12223 32814
rect 16021 32811 16087 32814
rect 0 32738 160 32768
rect 2773 32738 2839 32741
rect 11513 32738 11579 32741
rect 0 32736 2839 32738
rect 0 32680 2778 32736
rect 2834 32680 2839 32736
rect 0 32678 2839 32680
rect 0 32648 160 32678
rect 2773 32675 2839 32678
rect 9630 32736 11579 32738
rect 9630 32680 11518 32736
rect 11574 32680 11579 32736
rect 9630 32678 11579 32680
rect 6880 32672 7196 32673
rect 6880 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7196 32672
rect 6880 32607 7196 32608
rect 2497 32602 2563 32605
rect 6637 32602 6703 32605
rect 9630 32602 9690 32678
rect 11513 32675 11579 32678
rect 25221 32738 25287 32741
rect 25840 32738 26000 32768
rect 25221 32736 26000 32738
rect 25221 32680 25226 32736
rect 25282 32680 26000 32736
rect 25221 32678 26000 32680
rect 25221 32675 25287 32678
rect 12814 32672 13130 32673
rect 12814 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13130 32672
rect 12814 32607 13130 32608
rect 18748 32672 19064 32673
rect 18748 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19064 32672
rect 18748 32607 19064 32608
rect 24682 32672 24998 32673
rect 24682 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 24998 32672
rect 25840 32648 26000 32678
rect 24682 32607 24998 32608
rect 2497 32600 6703 32602
rect 2497 32544 2502 32600
rect 2558 32544 6642 32600
rect 6698 32544 6703 32600
rect 2497 32542 6703 32544
rect 2497 32539 2563 32542
rect 6637 32539 6703 32542
rect 7422 32542 9690 32602
rect 14181 32602 14247 32605
rect 15009 32602 15075 32605
rect 14181 32600 15075 32602
rect 14181 32544 14186 32600
rect 14242 32544 15014 32600
rect 15070 32544 15075 32600
rect 14181 32542 15075 32544
rect 0 32466 160 32496
rect 1209 32466 1275 32469
rect 0 32464 1275 32466
rect 0 32408 1214 32464
rect 1270 32408 1275 32464
rect 0 32406 1275 32408
rect 0 32376 160 32406
rect 1209 32403 1275 32406
rect 1853 32466 1919 32469
rect 7422 32466 7482 32542
rect 14181 32539 14247 32542
rect 15009 32539 15075 32542
rect 1853 32464 7482 32466
rect 1853 32408 1858 32464
rect 1914 32408 7482 32464
rect 1853 32406 7482 32408
rect 8201 32466 8267 32469
rect 19517 32466 19583 32469
rect 8201 32464 19583 32466
rect 8201 32408 8206 32464
rect 8262 32408 19522 32464
rect 19578 32408 19583 32464
rect 8201 32406 19583 32408
rect 1853 32403 1919 32406
rect 8201 32403 8267 32406
rect 19517 32403 19583 32406
rect 3550 32268 3556 32332
rect 3620 32330 3626 32332
rect 4613 32330 4679 32333
rect 3620 32328 4679 32330
rect 3620 32272 4618 32328
rect 4674 32272 4679 32328
rect 3620 32270 4679 32272
rect 3620 32268 3626 32270
rect 4613 32267 4679 32270
rect 10133 32330 10199 32333
rect 18137 32330 18203 32333
rect 10133 32328 18203 32330
rect 10133 32272 10138 32328
rect 10194 32272 18142 32328
rect 18198 32272 18203 32328
rect 10133 32270 18203 32272
rect 10133 32267 10199 32270
rect 18137 32267 18203 32270
rect 0 32194 160 32224
rect 1117 32194 1183 32197
rect 0 32192 1183 32194
rect 0 32136 1122 32192
rect 1178 32136 1183 32192
rect 0 32134 1183 32136
rect 0 32104 160 32134
rect 1117 32131 1183 32134
rect 24393 32194 24459 32197
rect 25840 32194 26000 32224
rect 24393 32192 26000 32194
rect 24393 32136 24398 32192
rect 24454 32136 26000 32192
rect 24393 32134 26000 32136
rect 24393 32131 24459 32134
rect 3913 32128 4229 32129
rect 3913 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4229 32128
rect 3913 32063 4229 32064
rect 9847 32128 10163 32129
rect 9847 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10163 32128
rect 9847 32063 10163 32064
rect 15781 32128 16097 32129
rect 15781 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16097 32128
rect 15781 32063 16097 32064
rect 21715 32128 22031 32129
rect 21715 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22031 32128
rect 25840 32104 26000 32134
rect 21715 32063 22031 32064
rect 0 31922 160 31952
rect 1209 31922 1275 31925
rect 0 31920 1275 31922
rect 0 31864 1214 31920
rect 1270 31864 1275 31920
rect 0 31862 1275 31864
rect 0 31832 160 31862
rect 1209 31859 1275 31862
rect 1485 31922 1551 31925
rect 6637 31922 6703 31925
rect 7097 31922 7163 31925
rect 1485 31920 7163 31922
rect 1485 31864 1490 31920
rect 1546 31864 6642 31920
rect 6698 31864 7102 31920
rect 7158 31864 7163 31920
rect 1485 31862 7163 31864
rect 1485 31859 1551 31862
rect 6637 31859 6703 31862
rect 7097 31859 7163 31862
rect 10869 31922 10935 31925
rect 13629 31922 13695 31925
rect 10869 31920 13695 31922
rect 10869 31864 10874 31920
rect 10930 31864 13634 31920
rect 13690 31864 13695 31920
rect 10869 31862 13695 31864
rect 10869 31859 10935 31862
rect 13629 31859 13695 31862
rect 15193 31922 15259 31925
rect 21541 31922 21607 31925
rect 15193 31920 21607 31922
rect 15193 31864 15198 31920
rect 15254 31864 21546 31920
rect 21602 31864 21607 31920
rect 15193 31862 21607 31864
rect 15193 31859 15259 31862
rect 21541 31859 21607 31862
rect 841 31786 907 31789
rect 5901 31786 5967 31789
rect 841 31784 5967 31786
rect 841 31728 846 31784
rect 902 31728 5906 31784
rect 5962 31728 5967 31784
rect 841 31726 5967 31728
rect 841 31723 907 31726
rect 5901 31723 5967 31726
rect 12014 31724 12020 31788
rect 12084 31786 12090 31788
rect 12617 31786 12683 31789
rect 12084 31784 12683 31786
rect 12084 31728 12622 31784
rect 12678 31728 12683 31784
rect 12084 31726 12683 31728
rect 12084 31724 12090 31726
rect 12617 31723 12683 31726
rect 0 31650 160 31680
rect 3785 31650 3851 31653
rect 0 31648 3851 31650
rect 0 31592 3790 31648
rect 3846 31592 3851 31648
rect 0 31590 3851 31592
rect 0 31560 160 31590
rect 3785 31587 3851 31590
rect 25129 31650 25195 31653
rect 25840 31650 26000 31680
rect 25129 31648 26000 31650
rect 25129 31592 25134 31648
rect 25190 31592 26000 31648
rect 25129 31590 26000 31592
rect 25129 31587 25195 31590
rect 6880 31584 7196 31585
rect 6880 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7196 31584
rect 6880 31519 7196 31520
rect 12814 31584 13130 31585
rect 12814 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13130 31584
rect 12814 31519 13130 31520
rect 18748 31584 19064 31585
rect 18748 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19064 31584
rect 18748 31519 19064 31520
rect 24682 31584 24998 31585
rect 24682 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 24998 31584
rect 25840 31560 26000 31590
rect 24682 31519 24998 31520
rect 4429 31514 4495 31517
rect 8569 31514 8635 31517
rect 12433 31514 12499 31517
rect 4429 31512 4722 31514
rect 4429 31456 4434 31512
rect 4490 31456 4722 31512
rect 4429 31454 4722 31456
rect 4429 31451 4495 31454
rect 0 31378 160 31408
rect 1393 31378 1459 31381
rect 4662 31380 4722 31454
rect 8569 31512 12499 31514
rect 8569 31456 8574 31512
rect 8630 31456 12438 31512
rect 12494 31456 12499 31512
rect 8569 31454 12499 31456
rect 8569 31451 8635 31454
rect 12433 31451 12499 31454
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 160 31318
rect 1393 31315 1459 31318
rect 4654 31316 4660 31380
rect 4724 31316 4730 31380
rect 5441 31378 5507 31381
rect 7414 31378 7420 31380
rect 5441 31376 7420 31378
rect 5441 31320 5446 31376
rect 5502 31320 7420 31376
rect 5441 31318 7420 31320
rect 5441 31315 5507 31318
rect 7414 31316 7420 31318
rect 7484 31316 7490 31380
rect 8017 31378 8083 31381
rect 16849 31378 16915 31381
rect 8017 31376 16915 31378
rect 8017 31320 8022 31376
rect 8078 31320 16854 31376
rect 16910 31320 16915 31376
rect 8017 31318 16915 31320
rect 8017 31315 8083 31318
rect 16849 31315 16915 31318
rect 4429 31242 4495 31245
rect 7598 31242 7604 31244
rect 4429 31240 7604 31242
rect 4429 31184 4434 31240
rect 4490 31184 7604 31240
rect 4429 31182 7604 31184
rect 4429 31179 4495 31182
rect 7598 31180 7604 31182
rect 7668 31180 7674 31244
rect 7833 31242 7899 31245
rect 21030 31242 21036 31244
rect 7833 31240 21036 31242
rect 7833 31184 7838 31240
rect 7894 31184 21036 31240
rect 7833 31182 21036 31184
rect 7833 31179 7899 31182
rect 21030 31180 21036 31182
rect 21100 31180 21106 31244
rect 0 31106 160 31136
rect 2773 31106 2839 31109
rect 0 31104 2839 31106
rect 0 31048 2778 31104
rect 2834 31048 2839 31104
rect 0 31046 2839 31048
rect 0 31016 160 31046
rect 2773 31043 2839 31046
rect 4889 31106 4955 31109
rect 9673 31106 9739 31109
rect 4889 31104 9739 31106
rect 4889 31048 4894 31104
rect 4950 31048 9678 31104
rect 9734 31048 9739 31104
rect 4889 31046 9739 31048
rect 4889 31043 4955 31046
rect 9673 31043 9739 31046
rect 11237 31106 11303 31109
rect 15101 31106 15167 31109
rect 11237 31104 15167 31106
rect 11237 31048 11242 31104
rect 11298 31048 15106 31104
rect 15162 31048 15167 31104
rect 11237 31046 15167 31048
rect 11237 31043 11303 31046
rect 15101 31043 15167 31046
rect 24393 31106 24459 31109
rect 25840 31106 26000 31136
rect 24393 31104 26000 31106
rect 24393 31048 24398 31104
rect 24454 31048 26000 31104
rect 24393 31046 26000 31048
rect 24393 31043 24459 31046
rect 3913 31040 4229 31041
rect 3913 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4229 31040
rect 3913 30975 4229 30976
rect 9847 31040 10163 31041
rect 9847 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10163 31040
rect 9847 30975 10163 30976
rect 15781 31040 16097 31041
rect 15781 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16097 31040
rect 15781 30975 16097 30976
rect 21715 31040 22031 31041
rect 21715 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22031 31040
rect 25840 31016 26000 31046
rect 21715 30975 22031 30976
rect 6177 30970 6243 30973
rect 8017 30970 8083 30973
rect 6177 30968 8083 30970
rect 6177 30912 6182 30968
rect 6238 30912 8022 30968
rect 8078 30912 8083 30968
rect 6177 30910 8083 30912
rect 6177 30907 6243 30910
rect 8017 30907 8083 30910
rect 0 30834 160 30864
rect 1301 30834 1367 30837
rect 0 30832 1367 30834
rect 0 30776 1306 30832
rect 1362 30776 1367 30832
rect 0 30774 1367 30776
rect 0 30744 160 30774
rect 1301 30771 1367 30774
rect 2405 30834 2471 30837
rect 5441 30834 5507 30837
rect 2405 30832 5507 30834
rect 2405 30776 2410 30832
rect 2466 30776 5446 30832
rect 5502 30776 5507 30832
rect 2405 30774 5507 30776
rect 2405 30771 2471 30774
rect 5441 30771 5507 30774
rect 2262 30636 2268 30700
rect 2332 30698 2338 30700
rect 2589 30698 2655 30701
rect 10133 30698 10199 30701
rect 2332 30696 10199 30698
rect 2332 30640 2594 30696
rect 2650 30640 10138 30696
rect 10194 30640 10199 30696
rect 2332 30638 10199 30640
rect 2332 30636 2338 30638
rect 2589 30635 2655 30638
rect 10133 30635 10199 30638
rect 11462 30636 11468 30700
rect 11532 30698 11538 30700
rect 12065 30698 12131 30701
rect 11532 30696 12131 30698
rect 11532 30640 12070 30696
rect 12126 30640 12131 30696
rect 11532 30638 12131 30640
rect 11532 30636 11538 30638
rect 12065 30635 12131 30638
rect 0 30562 160 30592
rect 3693 30562 3759 30565
rect 0 30560 3759 30562
rect 0 30504 3698 30560
rect 3754 30504 3759 30560
rect 0 30502 3759 30504
rect 0 30472 160 30502
rect 3693 30499 3759 30502
rect 25129 30562 25195 30565
rect 25840 30562 26000 30592
rect 25129 30560 26000 30562
rect 25129 30504 25134 30560
rect 25190 30504 26000 30560
rect 25129 30502 26000 30504
rect 25129 30499 25195 30502
rect 6880 30496 7196 30497
rect 6880 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7196 30496
rect 6880 30431 7196 30432
rect 12814 30496 13130 30497
rect 12814 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13130 30496
rect 12814 30431 13130 30432
rect 18748 30496 19064 30497
rect 18748 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19064 30496
rect 18748 30431 19064 30432
rect 24682 30496 24998 30497
rect 24682 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 24998 30496
rect 25840 30472 26000 30502
rect 24682 30431 24998 30432
rect 3141 30426 3207 30429
rect 3366 30426 3372 30428
rect 3141 30424 3372 30426
rect 3141 30368 3146 30424
rect 3202 30368 3372 30424
rect 3141 30366 3372 30368
rect 3141 30363 3207 30366
rect 3366 30364 3372 30366
rect 3436 30364 3442 30428
rect 3877 30426 3943 30429
rect 4889 30428 4955 30429
rect 3877 30424 4170 30426
rect 3877 30368 3882 30424
rect 3938 30368 4170 30424
rect 3877 30366 4170 30368
rect 3877 30363 3943 30366
rect 0 30290 160 30320
rect 3785 30290 3851 30293
rect 0 30288 3851 30290
rect 0 30232 3790 30288
rect 3846 30232 3851 30288
rect 0 30230 3851 30232
rect 4110 30290 4170 30366
rect 4838 30364 4844 30428
rect 4908 30426 4955 30428
rect 18413 30426 18479 30429
rect 4908 30424 5000 30426
rect 4950 30368 5000 30424
rect 4908 30366 5000 30368
rect 18278 30424 18479 30426
rect 18278 30368 18418 30424
rect 18474 30368 18479 30424
rect 18278 30366 18479 30368
rect 4908 30364 4955 30366
rect 4889 30363 4955 30364
rect 4470 30290 4476 30292
rect 4110 30230 4476 30290
rect 0 30200 160 30230
rect 3785 30227 3851 30230
rect 4470 30228 4476 30230
rect 4540 30228 4546 30292
rect 8753 30290 8819 30293
rect 4846 30288 8819 30290
rect 4846 30232 8758 30288
rect 8814 30232 8819 30288
rect 4846 30230 8819 30232
rect 1485 30154 1551 30157
rect 798 30152 1551 30154
rect 798 30096 1490 30152
rect 1546 30096 1551 30152
rect 798 30094 1551 30096
rect 0 30018 160 30048
rect 798 30018 858 30094
rect 1485 30091 1551 30094
rect 2129 30154 2195 30157
rect 4846 30154 4906 30230
rect 8753 30227 8819 30230
rect 18278 30157 18338 30366
rect 18413 30363 18479 30366
rect 21357 30426 21423 30429
rect 21582 30426 21588 30428
rect 21357 30424 21588 30426
rect 21357 30368 21362 30424
rect 21418 30368 21588 30424
rect 21357 30366 21588 30368
rect 21357 30363 21423 30366
rect 21582 30364 21588 30366
rect 21652 30364 21658 30428
rect 2129 30152 4906 30154
rect 2129 30096 2134 30152
rect 2190 30096 4906 30152
rect 2129 30094 4906 30096
rect 18229 30152 18338 30157
rect 18229 30096 18234 30152
rect 18290 30096 18338 30152
rect 18229 30094 18338 30096
rect 2129 30091 2195 30094
rect 18229 30091 18295 30094
rect 0 29958 858 30018
rect 24393 30018 24459 30021
rect 25840 30018 26000 30048
rect 24393 30016 26000 30018
rect 24393 29960 24398 30016
rect 24454 29960 26000 30016
rect 24393 29958 26000 29960
rect 0 29928 160 29958
rect 24393 29955 24459 29958
rect 3913 29952 4229 29953
rect 3913 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4229 29952
rect 3913 29887 4229 29888
rect 9847 29952 10163 29953
rect 9847 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10163 29952
rect 9847 29887 10163 29888
rect 15781 29952 16097 29953
rect 15781 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16097 29952
rect 15781 29887 16097 29888
rect 21715 29952 22031 29953
rect 21715 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22031 29952
rect 25840 29928 26000 29958
rect 21715 29887 22031 29888
rect 4294 29822 7850 29882
rect 0 29746 160 29776
rect 933 29746 999 29749
rect 0 29744 999 29746
rect 0 29688 938 29744
rect 994 29688 999 29744
rect 0 29686 999 29688
rect 0 29656 160 29686
rect 933 29683 999 29686
rect 2814 29684 2820 29748
rect 2884 29746 2890 29748
rect 4294 29746 4354 29822
rect 2884 29686 4354 29746
rect 4705 29746 4771 29749
rect 5390 29746 5396 29748
rect 4705 29744 5396 29746
rect 4705 29688 4710 29744
rect 4766 29688 5396 29744
rect 4705 29686 5396 29688
rect 2884 29684 2890 29686
rect 4705 29683 4771 29686
rect 5390 29684 5396 29686
rect 5460 29684 5466 29748
rect 7790 29746 7850 29822
rect 14089 29746 14155 29749
rect 6088 29686 7666 29746
rect 7790 29744 14155 29746
rect 7790 29688 14094 29744
rect 14150 29688 14155 29744
rect 7790 29686 14155 29688
rect 6088 29613 6148 29686
rect 6085 29608 6151 29613
rect 6085 29552 6090 29608
rect 6146 29552 6151 29608
rect 6085 29547 6151 29552
rect 7097 29610 7163 29613
rect 7606 29610 7666 29686
rect 14089 29683 14155 29686
rect 12709 29610 12775 29613
rect 13486 29610 13492 29612
rect 7097 29608 7482 29610
rect 7097 29552 7102 29608
rect 7158 29552 7482 29608
rect 7097 29550 7482 29552
rect 7606 29608 13492 29610
rect 7606 29552 12714 29608
rect 12770 29552 13492 29608
rect 7606 29550 13492 29552
rect 7097 29547 7163 29550
rect 0 29474 160 29504
rect 1301 29474 1367 29477
rect 0 29472 1367 29474
rect 0 29416 1306 29472
rect 1362 29416 1367 29472
rect 0 29414 1367 29416
rect 0 29384 160 29414
rect 1301 29411 1367 29414
rect 1577 29474 1643 29477
rect 6453 29474 6519 29477
rect 1577 29472 6519 29474
rect 1577 29416 1582 29472
rect 1638 29416 6458 29472
rect 6514 29416 6519 29472
rect 1577 29414 6519 29416
rect 7422 29474 7482 29550
rect 12709 29547 12775 29550
rect 13486 29548 13492 29550
rect 13556 29548 13562 29612
rect 7557 29474 7623 29477
rect 11053 29474 11119 29477
rect 7422 29472 11119 29474
rect 7422 29416 7562 29472
rect 7618 29416 11058 29472
rect 11114 29416 11119 29472
rect 7422 29414 11119 29416
rect 1577 29411 1643 29414
rect 6453 29411 6519 29414
rect 7557 29411 7623 29414
rect 11053 29411 11119 29414
rect 25129 29474 25195 29477
rect 25840 29474 26000 29504
rect 25129 29472 26000 29474
rect 25129 29416 25134 29472
rect 25190 29416 26000 29472
rect 25129 29414 26000 29416
rect 25129 29411 25195 29414
rect 6880 29408 7196 29409
rect 6880 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7196 29408
rect 6880 29343 7196 29344
rect 12814 29408 13130 29409
rect 12814 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13130 29408
rect 12814 29343 13130 29344
rect 18748 29408 19064 29409
rect 18748 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19064 29408
rect 18748 29343 19064 29344
rect 24682 29408 24998 29409
rect 24682 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 24998 29408
rect 25840 29384 26000 29414
rect 24682 29343 24998 29344
rect 565 29338 631 29341
rect 3233 29338 3299 29341
rect 6729 29338 6795 29341
rect 565 29336 3299 29338
rect 565 29280 570 29336
rect 626 29280 3238 29336
rect 3294 29280 3299 29336
rect 565 29278 3299 29280
rect 565 29275 631 29278
rect 3233 29275 3299 29278
rect 3558 29336 6795 29338
rect 3558 29280 6734 29336
rect 6790 29280 6795 29336
rect 3558 29278 6795 29280
rect 0 29202 160 29232
rect 3325 29202 3391 29205
rect 0 29200 3391 29202
rect 0 29144 3330 29200
rect 3386 29144 3391 29200
rect 0 29142 3391 29144
rect 0 29112 160 29142
rect 3325 29139 3391 29142
rect 2078 29004 2084 29068
rect 2148 29066 2154 29068
rect 3558 29066 3618 29278
rect 6729 29275 6795 29278
rect 10542 29276 10548 29340
rect 10612 29338 10618 29340
rect 10685 29338 10751 29341
rect 10612 29336 10751 29338
rect 10612 29280 10690 29336
rect 10746 29280 10751 29336
rect 10612 29278 10751 29280
rect 10612 29276 10618 29278
rect 10685 29275 10751 29278
rect 15377 29338 15443 29341
rect 16205 29338 16271 29341
rect 15377 29336 16271 29338
rect 15377 29280 15382 29336
rect 15438 29280 16210 29336
rect 16266 29280 16271 29336
rect 15377 29278 16271 29280
rect 15377 29275 15443 29278
rect 16205 29275 16271 29278
rect 7649 29202 7715 29205
rect 16614 29202 16620 29204
rect 7649 29200 16620 29202
rect 7649 29144 7654 29200
rect 7710 29144 16620 29200
rect 7649 29142 16620 29144
rect 7649 29139 7715 29142
rect 16614 29140 16620 29142
rect 16684 29202 16690 29204
rect 16941 29202 17007 29205
rect 16684 29200 17007 29202
rect 16684 29144 16946 29200
rect 17002 29144 17007 29200
rect 16684 29142 17007 29144
rect 16684 29140 16690 29142
rect 16941 29139 17007 29142
rect 2148 29006 3618 29066
rect 5165 29066 5231 29069
rect 5390 29066 5396 29068
rect 5165 29064 5396 29066
rect 5165 29008 5170 29064
rect 5226 29008 5396 29064
rect 5165 29006 5396 29008
rect 2148 29004 2154 29006
rect 5165 29003 5231 29006
rect 5390 29004 5396 29006
rect 5460 29004 5466 29068
rect 5625 29066 5691 29069
rect 6085 29066 6151 29069
rect 5625 29064 6151 29066
rect 5625 29008 5630 29064
rect 5686 29008 6090 29064
rect 6146 29008 6151 29064
rect 5625 29006 6151 29008
rect 5625 29003 5691 29006
rect 6085 29003 6151 29006
rect 7097 29066 7163 29069
rect 8293 29066 8359 29069
rect 7097 29064 8359 29066
rect 7097 29008 7102 29064
rect 7158 29008 8298 29064
rect 8354 29008 8359 29064
rect 7097 29006 8359 29008
rect 7097 29003 7163 29006
rect 8293 29003 8359 29006
rect 8937 29066 9003 29069
rect 10869 29066 10935 29069
rect 8937 29064 10935 29066
rect 8937 29008 8942 29064
rect 8998 29008 10874 29064
rect 10930 29008 10935 29064
rect 8937 29006 10935 29008
rect 8937 29003 9003 29006
rect 10869 29003 10935 29006
rect 11053 29066 11119 29069
rect 15561 29066 15627 29069
rect 11053 29064 15627 29066
rect 11053 29008 11058 29064
rect 11114 29008 15566 29064
rect 15622 29008 15627 29064
rect 11053 29006 15627 29008
rect 11053 29003 11119 29006
rect 15561 29003 15627 29006
rect 15745 29066 15811 29069
rect 16246 29066 16252 29068
rect 15745 29064 16252 29066
rect 15745 29008 15750 29064
rect 15806 29008 16252 29064
rect 15745 29006 16252 29008
rect 15745 29003 15811 29006
rect 16246 29004 16252 29006
rect 16316 29004 16322 29068
rect 0 28930 160 28960
rect 3601 28930 3667 28933
rect 0 28928 3667 28930
rect 0 28872 3606 28928
rect 3662 28872 3667 28928
rect 0 28870 3667 28872
rect 0 28840 160 28870
rect 3601 28867 3667 28870
rect 24393 28930 24459 28933
rect 25840 28930 26000 28960
rect 24393 28928 26000 28930
rect 24393 28872 24398 28928
rect 24454 28872 26000 28928
rect 24393 28870 26000 28872
rect 24393 28867 24459 28870
rect 3913 28864 4229 28865
rect 3913 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4229 28864
rect 3913 28799 4229 28800
rect 9847 28864 10163 28865
rect 9847 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10163 28864
rect 9847 28799 10163 28800
rect 15781 28864 16097 28865
rect 15781 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16097 28864
rect 15781 28799 16097 28800
rect 21715 28864 22031 28865
rect 21715 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22031 28864
rect 25840 28840 26000 28870
rect 21715 28799 22031 28800
rect 1485 28794 1551 28797
rect 798 28792 1551 28794
rect 798 28736 1490 28792
rect 1546 28736 1551 28792
rect 798 28734 1551 28736
rect 0 28658 160 28688
rect 798 28658 858 28734
rect 1485 28731 1551 28734
rect 4981 28794 5047 28797
rect 9397 28794 9463 28797
rect 4981 28792 9463 28794
rect 4981 28736 4986 28792
rect 5042 28736 9402 28792
rect 9458 28736 9463 28792
rect 4981 28734 9463 28736
rect 4981 28731 5047 28734
rect 9397 28731 9463 28734
rect 10358 28732 10364 28796
rect 10428 28794 10434 28796
rect 11881 28794 11947 28797
rect 10428 28792 11947 28794
rect 10428 28736 11886 28792
rect 11942 28736 11947 28792
rect 10428 28734 11947 28736
rect 10428 28732 10434 28734
rect 11881 28731 11947 28734
rect 16798 28732 16804 28796
rect 16868 28794 16874 28796
rect 17033 28794 17099 28797
rect 16868 28792 17099 28794
rect 16868 28736 17038 28792
rect 17094 28736 17099 28792
rect 16868 28734 17099 28736
rect 16868 28732 16874 28734
rect 17033 28731 17099 28734
rect 19425 28794 19491 28797
rect 20253 28794 20319 28797
rect 19425 28792 20319 28794
rect 19425 28736 19430 28792
rect 19486 28736 20258 28792
rect 20314 28736 20319 28792
rect 19425 28734 20319 28736
rect 19425 28731 19491 28734
rect 20253 28731 20319 28734
rect 1945 28660 2011 28661
rect 1894 28658 1900 28660
rect 0 28598 858 28658
rect 1854 28598 1900 28658
rect 1964 28658 2011 28660
rect 17033 28658 17099 28661
rect 17166 28658 17172 28660
rect 1964 28656 17172 28658
rect 2006 28600 17038 28656
rect 17094 28600 17172 28656
rect 0 28568 160 28598
rect 1894 28596 1900 28598
rect 1964 28598 17172 28600
rect 1964 28596 2011 28598
rect 1945 28595 2011 28596
rect 17033 28595 17099 28598
rect 17166 28596 17172 28598
rect 17236 28596 17242 28660
rect 2589 28524 2655 28525
rect 2589 28522 2636 28524
rect 2544 28520 2636 28522
rect 2544 28464 2594 28520
rect 2544 28462 2636 28464
rect 2589 28460 2636 28462
rect 2700 28460 2706 28524
rect 4153 28522 4219 28525
rect 4981 28524 5047 28525
rect 4981 28522 5028 28524
rect 4153 28520 5028 28522
rect 4153 28464 4158 28520
rect 4214 28464 4986 28520
rect 4153 28462 5028 28464
rect 2589 28459 2655 28460
rect 4153 28459 4219 28462
rect 4981 28460 5028 28462
rect 5092 28460 5098 28524
rect 7465 28522 7531 28525
rect 5168 28520 7531 28522
rect 5168 28464 7470 28520
rect 7526 28464 7531 28520
rect 5168 28462 7531 28464
rect 4981 28459 5047 28460
rect 0 28386 160 28416
rect 749 28386 815 28389
rect 0 28384 815 28386
rect 0 28328 754 28384
rect 810 28328 815 28384
rect 0 28326 815 28328
rect 0 28296 160 28326
rect 749 28323 815 28326
rect 1710 28324 1716 28388
rect 1780 28386 1786 28388
rect 2313 28386 2379 28389
rect 5168 28386 5228 28462
rect 7465 28459 7531 28462
rect 9397 28522 9463 28525
rect 13670 28522 13676 28524
rect 9397 28520 13676 28522
rect 9397 28464 9402 28520
rect 9458 28464 13676 28520
rect 9397 28462 13676 28464
rect 9397 28459 9463 28462
rect 13670 28460 13676 28462
rect 13740 28522 13746 28524
rect 14733 28522 14799 28525
rect 13740 28520 14799 28522
rect 13740 28464 14738 28520
rect 14794 28464 14799 28520
rect 13740 28462 14799 28464
rect 13740 28460 13746 28462
rect 14733 28459 14799 28462
rect 1780 28384 5228 28386
rect 1780 28328 2318 28384
rect 2374 28328 5228 28384
rect 1780 28326 5228 28328
rect 9581 28386 9647 28389
rect 11145 28386 11211 28389
rect 9581 28384 11211 28386
rect 9581 28328 9586 28384
rect 9642 28328 11150 28384
rect 11206 28328 11211 28384
rect 9581 28326 11211 28328
rect 1780 28324 1786 28326
rect 2313 28323 2379 28326
rect 9581 28323 9647 28326
rect 11145 28323 11211 28326
rect 13813 28386 13879 28389
rect 17861 28386 17927 28389
rect 13813 28384 17927 28386
rect 13813 28328 13818 28384
rect 13874 28328 17866 28384
rect 17922 28328 17927 28384
rect 13813 28326 17927 28328
rect 13813 28323 13879 28326
rect 17861 28323 17927 28326
rect 25129 28386 25195 28389
rect 25840 28386 26000 28416
rect 25129 28384 26000 28386
rect 25129 28328 25134 28384
rect 25190 28328 26000 28384
rect 25129 28326 26000 28328
rect 25129 28323 25195 28326
rect 6880 28320 7196 28321
rect 6880 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7196 28320
rect 6880 28255 7196 28256
rect 12814 28320 13130 28321
rect 12814 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13130 28320
rect 12814 28255 13130 28256
rect 18748 28320 19064 28321
rect 18748 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19064 28320
rect 18748 28255 19064 28256
rect 24682 28320 24998 28321
rect 24682 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 24998 28320
rect 25840 28296 26000 28326
rect 24682 28255 24998 28256
rect 606 28188 612 28252
rect 676 28250 682 28252
rect 5533 28250 5599 28253
rect 676 28248 5599 28250
rect 676 28192 5538 28248
rect 5594 28192 5599 28248
rect 676 28190 5599 28192
rect 676 28188 682 28190
rect 5533 28187 5599 28190
rect 7465 28250 7531 28253
rect 11513 28250 11579 28253
rect 7465 28248 11579 28250
rect 7465 28192 7470 28248
rect 7526 28192 11518 28248
rect 11574 28192 11579 28248
rect 7465 28190 11579 28192
rect 7465 28187 7531 28190
rect 11513 28187 11579 28190
rect 0 28114 160 28144
rect 3141 28114 3207 28117
rect 0 28112 3207 28114
rect 0 28056 3146 28112
rect 3202 28056 3207 28112
rect 0 28054 3207 28056
rect 0 28024 160 28054
rect 3141 28051 3207 28054
rect 4061 28114 4127 28117
rect 5257 28114 5323 28117
rect 4061 28112 5323 28114
rect 4061 28056 4066 28112
rect 4122 28056 5262 28112
rect 5318 28056 5323 28112
rect 4061 28054 5323 28056
rect 4061 28051 4127 28054
rect 5257 28051 5323 28054
rect 6821 28114 6887 28117
rect 13629 28114 13695 28117
rect 6821 28112 13695 28114
rect 6821 28056 6826 28112
rect 6882 28056 13634 28112
rect 13690 28056 13695 28112
rect 6821 28054 13695 28056
rect 6821 28051 6887 28054
rect 13629 28051 13695 28054
rect 19425 28114 19491 28117
rect 22185 28114 22251 28117
rect 19425 28112 22251 28114
rect 19425 28056 19430 28112
rect 19486 28056 22190 28112
rect 22246 28056 22251 28112
rect 19425 28054 22251 28056
rect 19425 28051 19491 28054
rect 22185 28051 22251 28054
rect 4245 27978 4311 27981
rect 5625 27978 5691 27981
rect 4245 27976 5691 27978
rect 4245 27920 4250 27976
rect 4306 27920 5630 27976
rect 5686 27920 5691 27976
rect 4245 27918 5691 27920
rect 4245 27915 4311 27918
rect 5625 27915 5691 27918
rect 6085 27978 6151 27981
rect 10501 27978 10567 27981
rect 6085 27976 10567 27978
rect 6085 27920 6090 27976
rect 6146 27920 10506 27976
rect 10562 27920 10567 27976
rect 6085 27918 10567 27920
rect 6085 27915 6151 27918
rect 10501 27915 10567 27918
rect 15009 27978 15075 27981
rect 20662 27978 20668 27980
rect 15009 27976 20668 27978
rect 15009 27920 15014 27976
rect 15070 27920 20668 27976
rect 15009 27918 20668 27920
rect 15009 27915 15075 27918
rect 20662 27916 20668 27918
rect 20732 27916 20738 27980
rect 0 27842 160 27872
rect 749 27842 815 27845
rect 0 27840 815 27842
rect 0 27784 754 27840
rect 810 27784 815 27840
rect 0 27782 815 27784
rect 0 27752 160 27782
rect 749 27779 815 27782
rect 4429 27842 4495 27845
rect 7189 27842 7255 27845
rect 4429 27840 7255 27842
rect 4429 27784 4434 27840
rect 4490 27784 7194 27840
rect 7250 27784 7255 27840
rect 4429 27782 7255 27784
rect 4429 27779 4495 27782
rect 7189 27779 7255 27782
rect 16246 27780 16252 27844
rect 16316 27842 16322 27844
rect 17125 27842 17191 27845
rect 16316 27840 17191 27842
rect 16316 27784 17130 27840
rect 17186 27784 17191 27840
rect 16316 27782 17191 27784
rect 16316 27780 16322 27782
rect 17125 27779 17191 27782
rect 24393 27842 24459 27845
rect 25840 27842 26000 27872
rect 24393 27840 26000 27842
rect 24393 27784 24398 27840
rect 24454 27784 26000 27840
rect 24393 27782 26000 27784
rect 24393 27779 24459 27782
rect 3913 27776 4229 27777
rect 3913 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4229 27776
rect 3913 27711 4229 27712
rect 9847 27776 10163 27777
rect 9847 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10163 27776
rect 9847 27711 10163 27712
rect 15781 27776 16097 27777
rect 15781 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16097 27776
rect 15781 27711 16097 27712
rect 21715 27776 22031 27777
rect 21715 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22031 27776
rect 25840 27752 26000 27782
rect 21715 27711 22031 27712
rect 2037 27706 2103 27709
rect 982 27704 2103 27706
rect 982 27648 2042 27704
rect 2098 27648 2103 27704
rect 982 27646 2103 27648
rect 0 27570 160 27600
rect 982 27570 1042 27646
rect 2037 27643 2103 27646
rect 11513 27706 11579 27709
rect 12341 27706 12407 27709
rect 11513 27704 12407 27706
rect 11513 27648 11518 27704
rect 11574 27648 12346 27704
rect 12402 27648 12407 27704
rect 11513 27646 12407 27648
rect 11513 27643 11579 27646
rect 12341 27643 12407 27646
rect 17534 27644 17540 27708
rect 17604 27706 17610 27708
rect 20846 27706 20852 27708
rect 17604 27646 20852 27706
rect 17604 27644 17610 27646
rect 20846 27644 20852 27646
rect 20916 27644 20922 27708
rect 2313 27570 2379 27573
rect 0 27510 1042 27570
rect 1166 27568 2379 27570
rect 1166 27512 2318 27568
rect 2374 27512 2379 27568
rect 1166 27510 2379 27512
rect 0 27480 160 27510
rect 0 27298 160 27328
rect 1166 27298 1226 27510
rect 2313 27507 2379 27510
rect 2681 27570 2747 27573
rect 7097 27570 7163 27573
rect 2681 27568 7163 27570
rect 2681 27512 2686 27568
rect 2742 27512 7102 27568
rect 7158 27512 7163 27568
rect 2681 27510 7163 27512
rect 2681 27507 2747 27510
rect 7097 27507 7163 27510
rect 10409 27570 10475 27573
rect 12249 27570 12315 27573
rect 10409 27568 12315 27570
rect 10409 27512 10414 27568
rect 10470 27512 12254 27568
rect 12310 27512 12315 27568
rect 10409 27510 12315 27512
rect 10409 27507 10475 27510
rect 12249 27507 12315 27510
rect 1761 27432 1827 27437
rect 2957 27436 3023 27437
rect 2957 27434 3004 27436
rect 1761 27376 1766 27432
rect 1822 27376 1827 27432
rect 1761 27371 1827 27376
rect 2912 27432 3004 27434
rect 2912 27376 2962 27432
rect 2912 27374 3004 27376
rect 2957 27372 3004 27374
rect 3068 27372 3074 27436
rect 5942 27372 5948 27436
rect 6012 27434 6018 27436
rect 7465 27434 7531 27437
rect 6012 27432 7531 27434
rect 6012 27376 7470 27432
rect 7526 27376 7531 27432
rect 6012 27374 7531 27376
rect 6012 27372 6018 27374
rect 2957 27371 3023 27372
rect 7465 27371 7531 27374
rect 0 27238 1226 27298
rect 0 27208 160 27238
rect 0 27026 160 27056
rect 1764 27026 1824 27371
rect 2957 27298 3023 27301
rect 6729 27298 6795 27301
rect 2957 27296 6795 27298
rect 2957 27240 2962 27296
rect 3018 27240 6734 27296
rect 6790 27240 6795 27296
rect 2957 27238 6795 27240
rect 2957 27235 3023 27238
rect 6729 27235 6795 27238
rect 25129 27298 25195 27301
rect 25840 27298 26000 27328
rect 25129 27296 26000 27298
rect 25129 27240 25134 27296
rect 25190 27240 26000 27296
rect 25129 27238 26000 27240
rect 25129 27235 25195 27238
rect 6880 27232 7196 27233
rect 6880 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7196 27232
rect 6880 27167 7196 27168
rect 12814 27232 13130 27233
rect 12814 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13130 27232
rect 12814 27167 13130 27168
rect 18748 27232 19064 27233
rect 18748 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19064 27232
rect 18748 27167 19064 27168
rect 24682 27232 24998 27233
rect 24682 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 24998 27232
rect 25840 27208 26000 27238
rect 24682 27167 24998 27168
rect 0 26966 1824 27026
rect 2221 27026 2287 27029
rect 7465 27026 7531 27029
rect 2221 27024 7531 27026
rect 2221 26968 2226 27024
rect 2282 26968 7470 27024
rect 7526 26968 7531 27024
rect 2221 26966 7531 26968
rect 0 26936 160 26966
rect 2221 26963 2287 26966
rect 7465 26963 7531 26966
rect 1342 26828 1348 26892
rect 1412 26890 1418 26892
rect 1577 26890 1643 26893
rect 1412 26888 1643 26890
rect 1412 26832 1582 26888
rect 1638 26832 1643 26888
rect 1412 26830 1643 26832
rect 1412 26828 1418 26830
rect 1534 26827 1643 26830
rect 1761 26890 1827 26893
rect 2078 26890 2084 26892
rect 1761 26888 2084 26890
rect 1761 26832 1766 26888
rect 1822 26832 2084 26888
rect 1761 26830 2084 26832
rect 1761 26827 1827 26830
rect 2078 26828 2084 26830
rect 2148 26828 2154 26892
rect 2773 26890 2839 26893
rect 7281 26890 7347 26893
rect 2773 26888 7347 26890
rect 2773 26832 2778 26888
rect 2834 26832 7286 26888
rect 7342 26832 7347 26888
rect 2773 26830 7347 26832
rect 2773 26827 2839 26830
rect 7281 26827 7347 26830
rect 20805 26892 20871 26893
rect 20805 26888 20852 26892
rect 20916 26890 20922 26892
rect 20805 26832 20810 26888
rect 20805 26828 20852 26832
rect 20916 26830 20962 26890
rect 20916 26828 20922 26830
rect 20805 26827 20871 26828
rect 0 26754 160 26784
rect 1534 26754 1594 26827
rect 2446 26754 2452 26756
rect 0 26694 1456 26754
rect 1534 26694 2452 26754
rect 0 26664 160 26694
rect 1396 26618 1456 26694
rect 2446 26692 2452 26694
rect 2516 26754 2522 26756
rect 2516 26694 2790 26754
rect 2516 26692 2522 26694
rect 2589 26618 2655 26621
rect 1396 26616 2655 26618
rect 1396 26560 2594 26616
rect 2650 26560 2655 26616
rect 1396 26558 2655 26560
rect 2589 26555 2655 26558
rect 0 26482 160 26512
rect 1209 26482 1275 26485
rect 0 26480 1275 26482
rect 0 26424 1214 26480
rect 1270 26424 1275 26480
rect 0 26422 1275 26424
rect 2730 26482 2790 26694
rect 11278 26692 11284 26756
rect 11348 26754 11354 26756
rect 13261 26754 13327 26757
rect 11348 26752 13327 26754
rect 11348 26696 13266 26752
rect 13322 26696 13327 26752
rect 11348 26694 13327 26696
rect 11348 26692 11354 26694
rect 13261 26691 13327 26694
rect 24393 26754 24459 26757
rect 25840 26754 26000 26784
rect 24393 26752 26000 26754
rect 24393 26696 24398 26752
rect 24454 26696 26000 26752
rect 24393 26694 26000 26696
rect 24393 26691 24459 26694
rect 3913 26688 4229 26689
rect 3913 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4229 26688
rect 3913 26623 4229 26624
rect 9847 26688 10163 26689
rect 9847 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10163 26688
rect 9847 26623 10163 26624
rect 15781 26688 16097 26689
rect 15781 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16097 26688
rect 15781 26623 16097 26624
rect 21715 26688 22031 26689
rect 21715 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22031 26688
rect 25840 26664 26000 26694
rect 21715 26623 22031 26624
rect 6729 26482 6795 26485
rect 2730 26480 6795 26482
rect 2730 26424 6734 26480
rect 6790 26424 6795 26480
rect 2730 26422 6795 26424
rect 0 26392 160 26422
rect 1209 26419 1275 26422
rect 6729 26419 6795 26422
rect 9254 26420 9260 26484
rect 9324 26482 9330 26484
rect 13537 26482 13603 26485
rect 9324 26480 13603 26482
rect 9324 26424 13542 26480
rect 13598 26424 13603 26480
rect 9324 26422 13603 26424
rect 9324 26420 9330 26422
rect 13537 26419 13603 26422
rect 1117 26346 1183 26349
rect 7649 26346 7715 26349
rect 10317 26346 10383 26349
rect 20713 26346 20779 26349
rect 1117 26344 7715 26346
rect 1117 26288 1122 26344
rect 1178 26288 7654 26344
rect 7710 26288 7715 26344
rect 1117 26286 7715 26288
rect 1117 26283 1183 26286
rect 7649 26283 7715 26286
rect 9630 26344 20779 26346
rect 9630 26288 10322 26344
rect 10378 26288 20718 26344
rect 20774 26288 20779 26344
rect 9630 26286 20779 26288
rect 0 26210 160 26240
rect 3785 26210 3851 26213
rect 0 26208 3851 26210
rect 0 26152 3790 26208
rect 3846 26152 3851 26208
rect 0 26150 3851 26152
rect 0 26120 160 26150
rect 3785 26147 3851 26150
rect 5533 26210 5599 26213
rect 6126 26210 6132 26212
rect 5533 26208 6132 26210
rect 5533 26152 5538 26208
rect 5594 26152 6132 26208
rect 5533 26150 6132 26152
rect 5533 26147 5599 26150
rect 6126 26148 6132 26150
rect 6196 26148 6202 26212
rect 8661 26210 8727 26213
rect 9630 26210 9690 26286
rect 10317 26283 10383 26286
rect 20713 26283 20779 26286
rect 8661 26208 9690 26210
rect 8661 26152 8666 26208
rect 8722 26152 9690 26208
rect 8661 26150 9690 26152
rect 25129 26210 25195 26213
rect 25840 26210 26000 26240
rect 25129 26208 26000 26210
rect 25129 26152 25134 26208
rect 25190 26152 26000 26208
rect 25129 26150 26000 26152
rect 8661 26147 8727 26150
rect 25129 26147 25195 26150
rect 6880 26144 7196 26145
rect 6880 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7196 26144
rect 6880 26079 7196 26080
rect 12814 26144 13130 26145
rect 12814 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13130 26144
rect 12814 26079 13130 26080
rect 18748 26144 19064 26145
rect 18748 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19064 26144
rect 18748 26079 19064 26080
rect 24682 26144 24998 26145
rect 24682 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 24998 26144
rect 25840 26120 26000 26150
rect 24682 26079 24998 26080
rect 2037 26074 2103 26077
rect 2262 26074 2268 26076
rect 2037 26072 2268 26074
rect 2037 26016 2042 26072
rect 2098 26016 2268 26072
rect 2037 26014 2268 26016
rect 2037 26011 2103 26014
rect 2262 26012 2268 26014
rect 2332 26012 2338 26076
rect 2446 26012 2452 26076
rect 2516 26074 2522 26076
rect 2773 26074 2839 26077
rect 2516 26072 2839 26074
rect 2516 26016 2778 26072
rect 2834 26016 2839 26072
rect 2516 26014 2839 26016
rect 2516 26012 2522 26014
rect 2773 26011 2839 26014
rect 10041 26074 10107 26077
rect 10041 26072 11162 26074
rect 10041 26016 10046 26072
rect 10102 26016 11162 26072
rect 10041 26014 11162 26016
rect 10041 26011 10107 26014
rect 0 25938 160 25968
rect 3417 25938 3483 25941
rect 0 25936 3483 25938
rect 0 25880 3422 25936
rect 3478 25880 3483 25936
rect 0 25878 3483 25880
rect 0 25848 160 25878
rect 3417 25875 3483 25878
rect 4654 25876 4660 25940
rect 4724 25938 4730 25940
rect 6494 25938 6500 25940
rect 4724 25878 6500 25938
rect 4724 25876 4730 25878
rect 6494 25876 6500 25878
rect 6564 25876 6570 25940
rect 7649 25938 7715 25941
rect 8937 25938 9003 25941
rect 10961 25938 11027 25941
rect 7649 25936 9003 25938
rect 7649 25880 7654 25936
rect 7710 25880 8942 25936
rect 8998 25880 9003 25936
rect 7649 25878 9003 25880
rect 7649 25875 7715 25878
rect 8937 25875 9003 25878
rect 10550 25936 11027 25938
rect 10550 25880 10966 25936
rect 11022 25880 11027 25936
rect 10550 25878 11027 25880
rect 11102 25938 11162 26014
rect 13445 25938 13511 25941
rect 11102 25936 13511 25938
rect 11102 25880 13450 25936
rect 13506 25880 13511 25936
rect 11102 25878 13511 25880
rect 1577 25802 1643 25805
rect 8753 25802 8819 25805
rect 9857 25802 9923 25805
rect 10550 25802 10610 25878
rect 10961 25875 11027 25878
rect 13445 25875 13511 25878
rect 1577 25800 8819 25802
rect 1577 25744 1582 25800
rect 1638 25744 8758 25800
rect 8814 25744 8819 25800
rect 1577 25742 8819 25744
rect 1577 25739 1643 25742
rect 8753 25739 8819 25742
rect 9630 25800 10610 25802
rect 9630 25744 9862 25800
rect 9918 25744 10610 25800
rect 9630 25742 10610 25744
rect 0 25666 160 25696
rect 2865 25666 2931 25669
rect 0 25664 2931 25666
rect 0 25608 2870 25664
rect 2926 25608 2931 25664
rect 0 25606 2931 25608
rect 0 25576 160 25606
rect 2865 25603 2931 25606
rect 4981 25666 5047 25669
rect 6126 25666 6132 25668
rect 4981 25664 6132 25666
rect 4981 25608 4986 25664
rect 5042 25608 6132 25664
rect 4981 25606 6132 25608
rect 4981 25603 5047 25606
rect 6126 25604 6132 25606
rect 6196 25604 6202 25668
rect 3913 25600 4229 25601
rect 3913 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4229 25600
rect 3913 25535 4229 25536
rect 6821 25530 6887 25533
rect 8753 25530 8819 25533
rect 6821 25528 8819 25530
rect 6821 25472 6826 25528
rect 6882 25472 8758 25528
rect 8814 25472 8819 25528
rect 6821 25470 8819 25472
rect 6821 25467 6887 25470
rect 8753 25467 8819 25470
rect 0 25394 160 25424
rect 1301 25394 1367 25397
rect 0 25392 1367 25394
rect 0 25336 1306 25392
rect 1362 25336 1367 25392
rect 0 25334 1367 25336
rect 0 25304 160 25334
rect 1301 25331 1367 25334
rect 1853 25394 1919 25397
rect 9630 25394 9690 25742
rect 9857 25739 9923 25742
rect 10726 25740 10732 25804
rect 10796 25802 10802 25804
rect 18229 25802 18295 25805
rect 10796 25800 18295 25802
rect 10796 25744 18234 25800
rect 18290 25744 18295 25800
rect 10796 25742 18295 25744
rect 10796 25740 10802 25742
rect 18229 25739 18295 25742
rect 24393 25666 24459 25669
rect 25840 25666 26000 25696
rect 24393 25664 26000 25666
rect 24393 25608 24398 25664
rect 24454 25608 26000 25664
rect 24393 25606 26000 25608
rect 24393 25603 24459 25606
rect 9847 25600 10163 25601
rect 9847 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10163 25600
rect 9847 25535 10163 25536
rect 15781 25600 16097 25601
rect 15781 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16097 25600
rect 15781 25535 16097 25536
rect 21715 25600 22031 25601
rect 21715 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22031 25600
rect 25840 25576 26000 25606
rect 21715 25535 22031 25536
rect 10317 25396 10383 25397
rect 10317 25394 10364 25396
rect 1853 25392 9690 25394
rect 1853 25336 1858 25392
rect 1914 25336 9690 25392
rect 1853 25334 9690 25336
rect 10272 25392 10364 25394
rect 10272 25336 10322 25392
rect 10272 25334 10364 25336
rect 1853 25331 1919 25334
rect 10317 25332 10364 25334
rect 10428 25332 10434 25396
rect 10317 25331 10383 25332
rect 1209 25256 1275 25261
rect 1209 25200 1214 25256
rect 1270 25200 1275 25256
rect 1209 25195 1275 25200
rect 1853 25258 1919 25261
rect 6821 25258 6887 25261
rect 1853 25256 6887 25258
rect 1853 25200 1858 25256
rect 1914 25200 6826 25256
rect 6882 25200 6887 25256
rect 1853 25198 6887 25200
rect 1853 25195 1919 25198
rect 6821 25195 6887 25198
rect 7005 25258 7071 25261
rect 8109 25258 8175 25261
rect 7005 25256 8175 25258
rect 7005 25200 7010 25256
rect 7066 25200 8114 25256
rect 8170 25200 8175 25256
rect 7005 25198 8175 25200
rect 7005 25195 7071 25198
rect 8109 25195 8175 25198
rect 16297 25258 16363 25261
rect 16614 25258 16620 25260
rect 16297 25256 16620 25258
rect 16297 25200 16302 25256
rect 16358 25200 16620 25256
rect 16297 25198 16620 25200
rect 16297 25195 16363 25198
rect 16614 25196 16620 25198
rect 16684 25258 16690 25260
rect 20069 25258 20135 25261
rect 16684 25256 20135 25258
rect 16684 25200 20074 25256
rect 20130 25200 20135 25256
rect 16684 25198 20135 25200
rect 16684 25196 16690 25198
rect 20069 25195 20135 25198
rect 21582 25196 21588 25260
rect 21652 25258 21658 25260
rect 25681 25258 25747 25261
rect 21652 25256 25747 25258
rect 21652 25200 25686 25256
rect 25742 25200 25747 25256
rect 21652 25198 25747 25200
rect 21652 25196 21658 25198
rect 25681 25195 25747 25198
rect 0 25122 160 25152
rect 1212 25122 1272 25195
rect 0 25062 1272 25122
rect 25129 25122 25195 25125
rect 25840 25122 26000 25152
rect 25129 25120 26000 25122
rect 25129 25064 25134 25120
rect 25190 25064 26000 25120
rect 25129 25062 26000 25064
rect 0 25032 160 25062
rect 25129 25059 25195 25062
rect 6880 25056 7196 25057
rect 6880 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7196 25056
rect 6880 24991 7196 24992
rect 12814 25056 13130 25057
rect 12814 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13130 25056
rect 12814 24991 13130 24992
rect 18748 25056 19064 25057
rect 18748 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19064 25056
rect 18748 24991 19064 24992
rect 24682 25056 24998 25057
rect 24682 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 24998 25056
rect 25840 25032 26000 25062
rect 24682 24991 24998 24992
rect 8201 24986 8267 24989
rect 11605 24986 11671 24989
rect 8201 24984 11671 24986
rect 8201 24928 8206 24984
rect 8262 24928 11610 24984
rect 11666 24928 11671 24984
rect 8201 24926 11671 24928
rect 8201 24923 8267 24926
rect 11605 24923 11671 24926
rect 0 24850 160 24880
rect 2129 24850 2195 24853
rect 0 24848 2195 24850
rect 0 24792 2134 24848
rect 2190 24792 2195 24848
rect 0 24790 2195 24792
rect 0 24760 160 24790
rect 2129 24787 2195 24790
rect 5574 24788 5580 24852
rect 5644 24850 5650 24852
rect 9489 24850 9555 24853
rect 5644 24848 9555 24850
rect 5644 24792 9494 24848
rect 9550 24792 9555 24848
rect 5644 24790 9555 24792
rect 5644 24788 5650 24790
rect 9489 24787 9555 24790
rect 16757 24850 16823 24853
rect 17493 24850 17559 24853
rect 16757 24848 17559 24850
rect 16757 24792 16762 24848
rect 16818 24792 17498 24848
rect 17554 24792 17559 24848
rect 16757 24790 17559 24792
rect 16757 24787 16823 24790
rect 17493 24787 17559 24790
rect 19701 24850 19767 24853
rect 21725 24850 21791 24853
rect 19701 24848 21791 24850
rect 19701 24792 19706 24848
rect 19762 24792 21730 24848
rect 21786 24792 21791 24848
rect 19701 24790 21791 24792
rect 19701 24787 19767 24790
rect 21725 24787 21791 24790
rect 381 24714 447 24717
rect 2865 24714 2931 24717
rect 5717 24714 5783 24717
rect 381 24712 2931 24714
rect 381 24656 386 24712
rect 442 24656 2870 24712
rect 2926 24656 2931 24712
rect 381 24654 2931 24656
rect 381 24651 447 24654
rect 2865 24651 2931 24654
rect 5582 24712 5783 24714
rect 5582 24656 5722 24712
rect 5778 24656 5783 24712
rect 5582 24654 5783 24656
rect 0 24578 160 24608
rect 1117 24578 1183 24581
rect 0 24576 1183 24578
rect 0 24520 1122 24576
rect 1178 24520 1183 24576
rect 0 24518 1183 24520
rect 0 24488 160 24518
rect 1117 24515 1183 24518
rect 3913 24512 4229 24513
rect 3913 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4229 24512
rect 3913 24447 4229 24448
rect 0 24306 160 24336
rect 5582 24309 5642 24654
rect 5717 24651 5783 24654
rect 10685 24714 10751 24717
rect 12198 24714 12204 24716
rect 10685 24712 12204 24714
rect 10685 24656 10690 24712
rect 10746 24656 12204 24712
rect 10685 24654 12204 24656
rect 10685 24651 10751 24654
rect 12198 24652 12204 24654
rect 12268 24652 12274 24716
rect 24393 24578 24459 24581
rect 25840 24578 26000 24608
rect 24393 24576 26000 24578
rect 24393 24520 24398 24576
rect 24454 24520 26000 24576
rect 24393 24518 26000 24520
rect 24393 24515 24459 24518
rect 9847 24512 10163 24513
rect 9847 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10163 24512
rect 9847 24447 10163 24448
rect 15781 24512 16097 24513
rect 15781 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16097 24512
rect 15781 24447 16097 24448
rect 21715 24512 22031 24513
rect 21715 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22031 24512
rect 25840 24488 26000 24518
rect 21715 24447 22031 24448
rect 1669 24306 1735 24309
rect 0 24304 1735 24306
rect 0 24248 1674 24304
rect 1730 24248 1735 24304
rect 0 24246 1735 24248
rect 0 24216 160 24246
rect 1669 24243 1735 24246
rect 2998 24244 3004 24308
rect 3068 24306 3074 24308
rect 5073 24306 5139 24309
rect 3068 24304 5139 24306
rect 3068 24248 5078 24304
rect 5134 24248 5139 24304
rect 3068 24246 5139 24248
rect 5582 24304 5691 24309
rect 10869 24308 10935 24309
rect 10869 24306 10916 24308
rect 5582 24248 5630 24304
rect 5686 24248 5691 24304
rect 5582 24246 5691 24248
rect 10824 24304 10916 24306
rect 10824 24248 10874 24304
rect 10824 24246 10916 24248
rect 3068 24244 3074 24246
rect 5073 24243 5139 24246
rect 5625 24243 5691 24246
rect 10869 24244 10916 24246
rect 10980 24244 10986 24308
rect 10869 24243 10935 24244
rect 933 24170 999 24173
rect 4061 24170 4127 24173
rect 933 24168 4127 24170
rect 933 24112 938 24168
rect 994 24112 4066 24168
rect 4122 24112 4127 24168
rect 933 24110 4127 24112
rect 933 24107 999 24110
rect 4061 24107 4127 24110
rect 0 24034 160 24064
rect 1393 24034 1459 24037
rect 0 24032 1459 24034
rect 0 23976 1398 24032
rect 1454 23976 1459 24032
rect 0 23974 1459 23976
rect 0 23944 160 23974
rect 1393 23971 1459 23974
rect 9581 24034 9647 24037
rect 12341 24034 12407 24037
rect 9581 24032 12407 24034
rect 9581 23976 9586 24032
rect 9642 23976 12346 24032
rect 12402 23976 12407 24032
rect 9581 23974 12407 23976
rect 9581 23971 9647 23974
rect 12341 23971 12407 23974
rect 25129 24034 25195 24037
rect 25840 24034 26000 24064
rect 25129 24032 26000 24034
rect 25129 23976 25134 24032
rect 25190 23976 26000 24032
rect 25129 23974 26000 23976
rect 25129 23971 25195 23974
rect 6880 23968 7196 23969
rect 6880 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7196 23968
rect 6880 23903 7196 23904
rect 12814 23968 13130 23969
rect 12814 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13130 23968
rect 12814 23903 13130 23904
rect 18748 23968 19064 23969
rect 18748 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19064 23968
rect 18748 23903 19064 23904
rect 24682 23968 24998 23969
rect 24682 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 24998 23968
rect 25840 23944 26000 23974
rect 24682 23903 24998 23904
rect 2773 23900 2839 23901
rect 2773 23898 2820 23900
rect 2728 23896 2820 23898
rect 2728 23840 2778 23896
rect 2728 23838 2820 23840
rect 2773 23836 2820 23838
rect 2884 23836 2890 23900
rect 9765 23898 9831 23901
rect 9765 23896 12082 23898
rect 9765 23840 9770 23896
rect 9826 23840 12082 23896
rect 9765 23838 12082 23840
rect 2773 23835 2839 23836
rect 9765 23835 9831 23838
rect 0 23762 160 23792
rect 1025 23762 1091 23765
rect 0 23760 1091 23762
rect 0 23704 1030 23760
rect 1086 23704 1091 23760
rect 0 23702 1091 23704
rect 0 23672 160 23702
rect 1025 23699 1091 23702
rect 1761 23762 1827 23765
rect 9581 23762 9647 23765
rect 1761 23760 9647 23762
rect 1761 23704 1766 23760
rect 1822 23704 9586 23760
rect 9642 23704 9647 23760
rect 1761 23702 9647 23704
rect 1761 23699 1827 23702
rect 9581 23699 9647 23702
rect 9765 23762 9831 23765
rect 11697 23762 11763 23765
rect 9765 23760 11763 23762
rect 9765 23704 9770 23760
rect 9826 23704 11702 23760
rect 11758 23704 11763 23760
rect 9765 23702 11763 23704
rect 12022 23762 12082 23838
rect 16573 23762 16639 23765
rect 12022 23760 16639 23762
rect 12022 23704 16578 23760
rect 16634 23704 16639 23760
rect 12022 23702 16639 23704
rect 9765 23699 9831 23702
rect 11697 23699 11763 23702
rect 16573 23699 16639 23702
rect 1301 23626 1367 23629
rect 10133 23626 10199 23629
rect 1301 23624 10199 23626
rect 1301 23568 1306 23624
rect 1362 23568 10138 23624
rect 10194 23568 10199 23624
rect 1301 23566 10199 23568
rect 1301 23563 1367 23566
rect 10133 23563 10199 23566
rect 21398 23564 21404 23628
rect 21468 23626 21474 23628
rect 23565 23626 23631 23629
rect 21468 23624 23631 23626
rect 21468 23568 23570 23624
rect 23626 23568 23631 23624
rect 21468 23566 23631 23568
rect 21468 23564 21474 23566
rect 23565 23563 23631 23566
rect 0 23490 160 23520
rect 749 23490 815 23493
rect 0 23488 815 23490
rect 0 23432 754 23488
rect 810 23432 815 23488
rect 0 23430 815 23432
rect 0 23400 160 23430
rect 749 23427 815 23430
rect 1710 23428 1716 23492
rect 1780 23490 1786 23492
rect 2129 23490 2195 23493
rect 1780 23488 2195 23490
rect 1780 23432 2134 23488
rect 2190 23432 2195 23488
rect 1780 23430 2195 23432
rect 1780 23428 1786 23430
rect 2129 23427 2195 23430
rect 4838 23428 4844 23492
rect 4908 23490 4914 23492
rect 4981 23490 5047 23493
rect 5942 23490 5948 23492
rect 4908 23488 5047 23490
rect 4908 23432 4986 23488
rect 5042 23432 5047 23488
rect 4908 23430 5047 23432
rect 4908 23428 4914 23430
rect 4981 23427 5047 23430
rect 5168 23430 5948 23490
rect 3913 23424 4229 23425
rect 3913 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4229 23424
rect 3913 23359 4229 23360
rect 0 23218 160 23248
rect 1577 23218 1643 23221
rect 0 23216 1643 23218
rect 0 23160 1582 23216
rect 1638 23160 1643 23216
rect 0 23158 1643 23160
rect 0 23128 160 23158
rect 1577 23155 1643 23158
rect 5168 23082 5228 23430
rect 5942 23428 5948 23430
rect 6012 23428 6018 23492
rect 6494 23428 6500 23492
rect 6564 23490 6570 23492
rect 9673 23490 9739 23493
rect 6564 23488 9739 23490
rect 6564 23432 9678 23488
rect 9734 23432 9739 23488
rect 6564 23430 9739 23432
rect 6564 23428 6570 23430
rect 9673 23427 9739 23430
rect 12249 23490 12315 23493
rect 13486 23490 13492 23492
rect 12249 23488 13492 23490
rect 12249 23432 12254 23488
rect 12310 23432 13492 23488
rect 12249 23430 13492 23432
rect 12249 23427 12315 23430
rect 13486 23428 13492 23430
rect 13556 23490 13562 23492
rect 14457 23490 14523 23493
rect 13556 23488 14523 23490
rect 13556 23432 14462 23488
rect 14518 23432 14523 23488
rect 13556 23430 14523 23432
rect 13556 23428 13562 23430
rect 14457 23427 14523 23430
rect 24393 23490 24459 23493
rect 25840 23490 26000 23520
rect 24393 23488 26000 23490
rect 24393 23432 24398 23488
rect 24454 23432 26000 23488
rect 24393 23430 26000 23432
rect 24393 23427 24459 23430
rect 9847 23424 10163 23425
rect 9847 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10163 23424
rect 9847 23359 10163 23360
rect 15781 23424 16097 23425
rect 15781 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16097 23424
rect 15781 23359 16097 23360
rect 21715 23424 22031 23425
rect 21715 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22031 23424
rect 25840 23400 26000 23430
rect 21715 23359 22031 23360
rect 13721 23356 13787 23357
rect 13670 23292 13676 23356
rect 13740 23354 13787 23356
rect 13740 23352 13832 23354
rect 13782 23296 13832 23352
rect 13740 23294 13832 23296
rect 13740 23292 13787 23294
rect 13721 23291 13787 23292
rect 5441 23218 5507 23221
rect 10133 23218 10199 23221
rect 5441 23216 10199 23218
rect 5441 23160 5446 23216
rect 5502 23160 10138 23216
rect 10194 23160 10199 23216
rect 5441 23158 10199 23160
rect 5441 23155 5507 23158
rect 10133 23155 10199 23158
rect 11646 23156 11652 23220
rect 11716 23218 11722 23220
rect 13537 23218 13603 23221
rect 11716 23216 13603 23218
rect 11716 23160 13542 23216
rect 13598 23160 13603 23216
rect 11716 23158 13603 23160
rect 11716 23156 11722 23158
rect 13537 23155 13603 23158
rect 2730 23022 5228 23082
rect 6453 23082 6519 23085
rect 8109 23082 8175 23085
rect 17534 23082 17540 23084
rect 6453 23080 7482 23082
rect 6453 23024 6458 23080
rect 6514 23024 7482 23080
rect 6453 23022 7482 23024
rect 0 22946 160 22976
rect 1301 22946 1367 22949
rect 0 22944 1367 22946
rect 0 22888 1306 22944
rect 1362 22888 1367 22944
rect 0 22886 1367 22888
rect 0 22856 160 22886
rect 1301 22883 1367 22886
rect 0 22674 160 22704
rect 0 22614 1594 22674
rect 0 22584 160 22614
rect 1534 22538 1594 22614
rect 2262 22612 2268 22676
rect 2332 22674 2338 22676
rect 2730 22674 2790 23022
rect 6453 23019 6519 23022
rect 3969 22946 4035 22949
rect 3006 22944 4035 22946
rect 3006 22888 3974 22944
rect 4030 22888 4035 22944
rect 3006 22886 4035 22888
rect 7422 22946 7482 23022
rect 8109 23080 17540 23082
rect 8109 23024 8114 23080
rect 8170 23024 17540 23080
rect 8109 23022 17540 23024
rect 8109 23019 8175 23022
rect 17534 23020 17540 23022
rect 17604 23020 17610 23084
rect 12014 22946 12020 22948
rect 7422 22886 12020 22946
rect 2332 22614 2790 22674
rect 2865 22672 2931 22677
rect 2865 22616 2870 22672
rect 2926 22616 2931 22672
rect 2332 22612 2338 22614
rect 2865 22611 2931 22616
rect 2868 22538 2928 22611
rect 1534 22478 2928 22538
rect 0 22402 160 22432
rect 1485 22402 1551 22405
rect 0 22400 1551 22402
rect 0 22344 1490 22400
rect 1546 22344 1551 22400
rect 0 22342 1551 22344
rect 0 22312 160 22342
rect 1485 22339 1551 22342
rect 381 22266 447 22269
rect 3006 22266 3066 22886
rect 3969 22883 4035 22886
rect 12014 22884 12020 22886
rect 12084 22884 12090 22948
rect 13537 22946 13603 22949
rect 13670 22946 13676 22948
rect 13537 22944 13676 22946
rect 13537 22888 13542 22944
rect 13598 22888 13676 22944
rect 13537 22886 13676 22888
rect 13537 22883 13603 22886
rect 13670 22884 13676 22886
rect 13740 22884 13746 22948
rect 25129 22946 25195 22949
rect 25840 22946 26000 22976
rect 25129 22944 26000 22946
rect 25129 22888 25134 22944
rect 25190 22888 26000 22944
rect 25129 22886 26000 22888
rect 25129 22883 25195 22886
rect 6880 22880 7196 22881
rect 6880 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7196 22880
rect 6880 22815 7196 22816
rect 12814 22880 13130 22881
rect 12814 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13130 22880
rect 12814 22815 13130 22816
rect 18748 22880 19064 22881
rect 18748 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19064 22880
rect 18748 22815 19064 22816
rect 24682 22880 24998 22881
rect 24682 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 24998 22880
rect 25840 22856 26000 22886
rect 24682 22815 24998 22816
rect 4613 22812 4679 22813
rect 4613 22808 4660 22812
rect 4724 22810 4730 22812
rect 4613 22752 4618 22808
rect 4613 22748 4660 22752
rect 4724 22750 4770 22810
rect 4724 22748 4730 22750
rect 4613 22747 4679 22748
rect 3141 22674 3207 22677
rect 3141 22672 12450 22674
rect 3141 22616 3146 22672
rect 3202 22616 12450 22672
rect 3141 22614 12450 22616
rect 3141 22611 3207 22614
rect 11094 22538 11100 22540
rect 381 22264 3066 22266
rect 381 22208 386 22264
rect 442 22208 3066 22264
rect 381 22206 3066 22208
rect 3374 22478 11100 22538
rect 381 22203 447 22206
rect 0 22130 160 22160
rect 3233 22130 3299 22133
rect 0 22128 3299 22130
rect 0 22072 3238 22128
rect 3294 22072 3299 22128
rect 0 22070 3299 22072
rect 0 22040 160 22070
rect 3233 22067 3299 22070
rect 1761 21994 1827 21997
rect 1894 21994 1900 21996
rect 1761 21992 1900 21994
rect 1761 21936 1766 21992
rect 1822 21936 1900 21992
rect 1761 21934 1900 21936
rect 1761 21931 1827 21934
rect 1894 21932 1900 21934
rect 1964 21932 1970 21996
rect 0 21858 160 21888
rect 1301 21858 1367 21861
rect 0 21856 1367 21858
rect 0 21800 1306 21856
rect 1362 21800 1367 21856
rect 0 21798 1367 21800
rect 0 21768 160 21798
rect 1301 21795 1367 21798
rect 3233 21858 3299 21861
rect 3374 21858 3434 22478
rect 11094 22476 11100 22478
rect 11164 22476 11170 22540
rect 11462 22476 11468 22540
rect 11532 22538 11538 22540
rect 11789 22538 11855 22541
rect 11532 22536 11855 22538
rect 11532 22480 11794 22536
rect 11850 22480 11855 22536
rect 11532 22478 11855 22480
rect 12390 22538 12450 22614
rect 16113 22538 16179 22541
rect 12390 22536 16179 22538
rect 12390 22480 16118 22536
rect 16174 22480 16179 22536
rect 12390 22478 16179 22480
rect 11532 22476 11538 22478
rect 11789 22475 11855 22478
rect 16113 22475 16179 22478
rect 21725 22538 21791 22541
rect 22461 22538 22527 22541
rect 21725 22536 22527 22538
rect 21725 22480 21730 22536
rect 21786 22480 22466 22536
rect 22522 22480 22527 22536
rect 21725 22478 22527 22480
rect 21725 22475 21791 22478
rect 22461 22475 22527 22478
rect 24485 22402 24551 22405
rect 25840 22402 26000 22432
rect 24485 22400 26000 22402
rect 24485 22344 24490 22400
rect 24546 22344 26000 22400
rect 24485 22342 26000 22344
rect 24485 22339 24551 22342
rect 3913 22336 4229 22337
rect 3913 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4229 22336
rect 3913 22271 4229 22272
rect 9847 22336 10163 22337
rect 9847 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10163 22336
rect 9847 22271 10163 22272
rect 15781 22336 16097 22337
rect 15781 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16097 22336
rect 15781 22271 16097 22272
rect 21715 22336 22031 22337
rect 21715 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22031 22336
rect 25840 22312 26000 22342
rect 21715 22271 22031 22272
rect 4613 22266 4679 22269
rect 8477 22266 8543 22269
rect 9581 22266 9647 22269
rect 4613 22264 9647 22266
rect 4613 22208 4618 22264
rect 4674 22208 8482 22264
rect 8538 22208 9586 22264
rect 9642 22208 9647 22264
rect 4613 22206 9647 22208
rect 4613 22203 4679 22206
rect 8477 22203 8543 22206
rect 9581 22203 9647 22206
rect 3969 22130 4035 22133
rect 5257 22130 5323 22133
rect 3969 22128 5323 22130
rect 3969 22072 3974 22128
rect 4030 22072 5262 22128
rect 5318 22072 5323 22128
rect 3969 22070 5323 22072
rect 3969 22067 4035 22070
rect 5257 22067 5323 22070
rect 6821 22130 6887 22133
rect 11697 22130 11763 22133
rect 6821 22128 11763 22130
rect 6821 22072 6826 22128
rect 6882 22072 11702 22128
rect 11758 22072 11763 22128
rect 6821 22070 11763 22072
rect 6821 22067 6887 22070
rect 11697 22067 11763 22070
rect 5390 21932 5396 21996
rect 5460 21994 5466 21996
rect 5460 21934 10058 21994
rect 5460 21932 5466 21934
rect 6177 21860 6243 21861
rect 6126 21858 6132 21860
rect 3233 21856 3434 21858
rect 3233 21800 3238 21856
rect 3294 21800 3434 21856
rect 3233 21798 3434 21800
rect 6086 21798 6132 21858
rect 6196 21856 6243 21860
rect 6238 21800 6243 21856
rect 3233 21795 3299 21798
rect 6126 21796 6132 21798
rect 6196 21796 6243 21800
rect 6177 21795 6243 21796
rect 7649 21858 7715 21861
rect 9254 21858 9260 21860
rect 7649 21856 9260 21858
rect 7649 21800 7654 21856
rect 7710 21800 9260 21856
rect 7649 21798 9260 21800
rect 7649 21795 7715 21798
rect 9254 21796 9260 21798
rect 9324 21796 9330 21860
rect 6880 21792 7196 21793
rect 6880 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7196 21792
rect 6880 21727 7196 21728
rect 1669 21722 1735 21725
rect 3417 21722 3483 21725
rect 1669 21720 3483 21722
rect 1669 21664 1674 21720
rect 1730 21664 3422 21720
rect 3478 21664 3483 21720
rect 1669 21662 3483 21664
rect 1669 21659 1735 21662
rect 3417 21659 3483 21662
rect 0 21586 160 21616
rect 1209 21586 1275 21589
rect 0 21584 1275 21586
rect 0 21528 1214 21584
rect 1270 21528 1275 21584
rect 0 21526 1275 21528
rect 0 21496 160 21526
rect 1209 21523 1275 21526
rect 4613 21586 4679 21589
rect 9857 21586 9923 21589
rect 4613 21584 9923 21586
rect 4613 21528 4618 21584
rect 4674 21528 9862 21584
rect 9918 21528 9923 21584
rect 4613 21526 9923 21528
rect 9998 21586 10058 21934
rect 25129 21858 25195 21861
rect 25840 21858 26000 21888
rect 25129 21856 26000 21858
rect 25129 21800 25134 21856
rect 25190 21800 26000 21856
rect 25129 21798 26000 21800
rect 25129 21795 25195 21798
rect 12814 21792 13130 21793
rect 12814 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13130 21792
rect 12814 21727 13130 21728
rect 18748 21792 19064 21793
rect 18748 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19064 21792
rect 18748 21727 19064 21728
rect 24682 21792 24998 21793
rect 24682 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 24998 21792
rect 25840 21768 26000 21798
rect 24682 21727 24998 21728
rect 16757 21724 16823 21725
rect 16757 21722 16804 21724
rect 16712 21720 16804 21722
rect 16712 21664 16762 21720
rect 16712 21662 16804 21664
rect 16757 21660 16804 21662
rect 16868 21660 16874 21724
rect 16941 21722 17007 21725
rect 17493 21722 17559 21725
rect 16941 21720 17559 21722
rect 16941 21664 16946 21720
rect 17002 21664 17498 21720
rect 17554 21664 17559 21720
rect 16941 21662 17559 21664
rect 16757 21659 16823 21660
rect 16941 21659 17007 21662
rect 17493 21659 17559 21662
rect 10869 21586 10935 21589
rect 16573 21586 16639 21589
rect 17217 21586 17283 21589
rect 9998 21584 17283 21586
rect 9998 21528 10874 21584
rect 10930 21528 16578 21584
rect 16634 21528 17222 21584
rect 17278 21528 17283 21584
rect 9998 21526 17283 21528
rect 4613 21523 4679 21526
rect 9857 21523 9923 21526
rect 10869 21523 10935 21526
rect 16573 21523 16639 21526
rect 17217 21523 17283 21526
rect 2129 21450 2195 21453
rect 6085 21450 6151 21453
rect 2129 21448 6151 21450
rect 2129 21392 2134 21448
rect 2190 21392 6090 21448
rect 6146 21392 6151 21448
rect 2129 21390 6151 21392
rect 2129 21387 2195 21390
rect 6085 21387 6151 21390
rect 7833 21450 7899 21453
rect 22185 21450 22251 21453
rect 7833 21448 22251 21450
rect 7833 21392 7838 21448
rect 7894 21392 22190 21448
rect 22246 21392 22251 21448
rect 7833 21390 22251 21392
rect 7833 21387 7899 21390
rect 22185 21387 22251 21390
rect 0 21314 160 21344
rect 1209 21314 1275 21317
rect 0 21312 1275 21314
rect 0 21256 1214 21312
rect 1270 21256 1275 21312
rect 0 21254 1275 21256
rect 0 21224 160 21254
rect 1209 21251 1275 21254
rect 4889 21314 4955 21317
rect 7833 21314 7899 21317
rect 4889 21312 7899 21314
rect 4889 21256 4894 21312
rect 4950 21256 7838 21312
rect 7894 21256 7899 21312
rect 4889 21254 7899 21256
rect 4889 21251 4955 21254
rect 7833 21251 7899 21254
rect 23841 21314 23907 21317
rect 25840 21314 26000 21344
rect 23841 21312 26000 21314
rect 23841 21256 23846 21312
rect 23902 21256 26000 21312
rect 23841 21254 26000 21256
rect 23841 21251 23907 21254
rect 3913 21248 4229 21249
rect 3913 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4229 21248
rect 3913 21183 4229 21184
rect 9847 21248 10163 21249
rect 9847 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10163 21248
rect 9847 21183 10163 21184
rect 15781 21248 16097 21249
rect 15781 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16097 21248
rect 15781 21183 16097 21184
rect 21715 21248 22031 21249
rect 21715 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22031 21248
rect 25840 21224 26000 21254
rect 21715 21183 22031 21184
rect 4429 21178 4495 21181
rect 5073 21178 5139 21181
rect 4429 21176 5139 21178
rect 4429 21120 4434 21176
rect 4490 21120 5078 21176
rect 5134 21120 5139 21176
rect 4429 21118 5139 21120
rect 4429 21115 4495 21118
rect 5073 21115 5139 21118
rect 8293 21178 8359 21181
rect 9581 21178 9647 21181
rect 12525 21178 12591 21181
rect 13445 21178 13511 21181
rect 15377 21178 15443 21181
rect 8293 21176 9647 21178
rect 8293 21120 8298 21176
rect 8354 21120 9586 21176
rect 9642 21120 9647 21176
rect 8293 21118 9647 21120
rect 8293 21115 8359 21118
rect 9581 21115 9647 21118
rect 12390 21176 15443 21178
rect 12390 21120 12530 21176
rect 12586 21120 13450 21176
rect 13506 21120 15382 21176
rect 15438 21120 15443 21176
rect 12390 21118 15443 21120
rect 0 21042 160 21072
rect 1301 21042 1367 21045
rect 0 21040 1367 21042
rect 0 20984 1306 21040
rect 1362 20984 1367 21040
rect 0 20982 1367 20984
rect 0 20952 160 20982
rect 1301 20979 1367 20982
rect 2589 21042 2655 21045
rect 4470 21042 4476 21044
rect 2589 21040 4476 21042
rect 2589 20984 2594 21040
rect 2650 20984 4476 21040
rect 2589 20982 4476 20984
rect 2589 20979 2655 20982
rect 4470 20980 4476 20982
rect 4540 21042 4546 21044
rect 10593 21042 10659 21045
rect 4540 21040 10659 21042
rect 4540 20984 10598 21040
rect 10654 20984 10659 21040
rect 4540 20982 10659 20984
rect 4540 20980 4546 20982
rect 10593 20979 10659 20982
rect 1209 20906 1275 20909
rect 1342 20906 1348 20908
rect 1209 20904 1348 20906
rect 1209 20848 1214 20904
rect 1270 20848 1348 20904
rect 1209 20846 1348 20848
rect 1209 20843 1275 20846
rect 1342 20844 1348 20846
rect 1412 20844 1418 20908
rect 1853 20906 1919 20909
rect 4889 20906 4955 20909
rect 1853 20904 4955 20906
rect 1853 20848 1858 20904
rect 1914 20848 4894 20904
rect 4950 20848 4955 20904
rect 1853 20846 4955 20848
rect 1853 20843 1919 20846
rect 4889 20843 4955 20846
rect 5390 20844 5396 20908
rect 5460 20844 5466 20908
rect 7189 20906 7255 20909
rect 7833 20906 7899 20909
rect 12390 20906 12450 21118
rect 12525 21115 12591 21118
rect 13445 21115 13511 21118
rect 15377 21115 15443 21118
rect 7189 20904 7712 20906
rect 7189 20848 7194 20904
rect 7250 20848 7712 20904
rect 7189 20846 7712 20848
rect 0 20770 160 20800
rect 1301 20770 1367 20773
rect 0 20768 1367 20770
rect 0 20712 1306 20768
rect 1362 20712 1367 20768
rect 0 20710 1367 20712
rect 0 20680 160 20710
rect 1301 20707 1367 20710
rect 2313 20770 2379 20773
rect 4153 20770 4219 20773
rect 5398 20770 5458 20844
rect 7189 20843 7255 20846
rect 2313 20768 5458 20770
rect 2313 20712 2318 20768
rect 2374 20712 4158 20768
rect 4214 20712 5458 20768
rect 2313 20710 5458 20712
rect 7652 20770 7712 20846
rect 7833 20904 12450 20906
rect 7833 20848 7838 20904
rect 7894 20848 12450 20904
rect 7833 20846 12450 20848
rect 12574 20846 13370 20906
rect 7833 20843 7899 20846
rect 8109 20770 8175 20773
rect 12574 20770 12634 20846
rect 7652 20768 12634 20770
rect 7652 20712 8114 20768
rect 8170 20712 12634 20768
rect 7652 20710 12634 20712
rect 13310 20770 13370 20846
rect 14181 20770 14247 20773
rect 14733 20770 14799 20773
rect 13310 20768 14799 20770
rect 13310 20712 14186 20768
rect 14242 20712 14738 20768
rect 14794 20712 14799 20768
rect 13310 20710 14799 20712
rect 2313 20707 2379 20710
rect 4153 20707 4219 20710
rect 8109 20707 8175 20710
rect 14181 20707 14247 20710
rect 14733 20707 14799 20710
rect 25129 20770 25195 20773
rect 25840 20770 26000 20800
rect 25129 20768 26000 20770
rect 25129 20712 25134 20768
rect 25190 20712 26000 20768
rect 25129 20710 26000 20712
rect 25129 20707 25195 20710
rect 6880 20704 7196 20705
rect 6880 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7196 20704
rect 6880 20639 7196 20640
rect 12814 20704 13130 20705
rect 12814 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13130 20704
rect 12814 20639 13130 20640
rect 18748 20704 19064 20705
rect 18748 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19064 20704
rect 18748 20639 19064 20640
rect 24682 20704 24998 20705
rect 24682 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 24998 20704
rect 25840 20680 26000 20710
rect 24682 20639 24998 20640
rect 9765 20634 9831 20637
rect 9765 20632 12634 20634
rect 9765 20576 9770 20632
rect 9826 20576 12634 20632
rect 9765 20574 12634 20576
rect 9765 20571 9831 20574
rect 0 20498 160 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 160 20438
rect 1393 20435 1459 20438
rect 2037 20498 2103 20501
rect 11421 20498 11487 20501
rect 2037 20496 2790 20498
rect 2037 20440 2042 20496
rect 2098 20440 2790 20496
rect 2037 20438 2790 20440
rect 2037 20435 2103 20438
rect 2730 20362 2790 20438
rect 9124 20496 11487 20498
rect 9124 20440 11426 20496
rect 11482 20440 11487 20496
rect 9124 20438 11487 20440
rect 12574 20498 12634 20574
rect 17861 20498 17927 20501
rect 12574 20496 17927 20498
rect 12574 20440 17866 20496
rect 17922 20440 17927 20496
rect 12574 20438 17927 20440
rect 2730 20302 7482 20362
rect 0 20226 160 20256
rect 749 20226 815 20229
rect 2957 20228 3023 20229
rect 2957 20226 3004 20228
rect 0 20224 815 20226
rect 0 20168 754 20224
rect 810 20168 815 20224
rect 0 20166 815 20168
rect 2912 20224 3004 20226
rect 2912 20168 2962 20224
rect 2912 20166 3004 20168
rect 0 20136 160 20166
rect 749 20163 815 20166
rect 2957 20164 3004 20166
rect 3068 20164 3074 20228
rect 7422 20226 7482 20302
rect 8845 20226 8911 20229
rect 9124 20226 9184 20438
rect 11421 20435 11487 20438
rect 17861 20435 17927 20438
rect 9254 20300 9260 20364
rect 9324 20362 9330 20364
rect 9324 20302 12450 20362
rect 9324 20300 9330 20302
rect 7422 20224 9184 20226
rect 7422 20168 8850 20224
rect 8906 20168 9184 20224
rect 7422 20166 9184 20168
rect 2957 20163 3023 20164
rect 8845 20163 8911 20166
rect 3913 20160 4229 20161
rect 3913 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4229 20160
rect 3913 20095 4229 20096
rect 9847 20160 10163 20161
rect 9847 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10163 20160
rect 9847 20095 10163 20096
rect 289 20090 355 20093
rect 4613 20090 4679 20093
rect 9121 20090 9187 20093
rect 11237 20090 11303 20093
rect 289 20088 3802 20090
rect 289 20032 294 20088
rect 350 20032 3802 20088
rect 289 20030 3802 20032
rect 289 20027 355 20030
rect 0 19954 160 19984
rect 841 19954 907 19957
rect 0 19952 907 19954
rect 0 19896 846 19952
rect 902 19896 907 19952
rect 0 19894 907 19896
rect 3742 19954 3802 20030
rect 4613 20088 9187 20090
rect 4613 20032 4618 20088
rect 4674 20032 9126 20088
rect 9182 20032 9187 20088
rect 4613 20030 9187 20032
rect 4613 20027 4679 20030
rect 9121 20027 9187 20030
rect 10366 20088 11303 20090
rect 10366 20032 11242 20088
rect 11298 20032 11303 20088
rect 10366 20030 11303 20032
rect 10366 19954 10426 20030
rect 11237 20027 11303 20030
rect 3742 19894 10426 19954
rect 12390 19954 12450 20302
rect 24025 20226 24091 20229
rect 25840 20226 26000 20256
rect 24025 20224 26000 20226
rect 24025 20168 24030 20224
rect 24086 20168 26000 20224
rect 24025 20166 26000 20168
rect 24025 20163 24091 20166
rect 15781 20160 16097 20161
rect 15781 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16097 20160
rect 15781 20095 16097 20096
rect 21715 20160 22031 20161
rect 21715 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22031 20160
rect 25840 20136 26000 20166
rect 21715 20095 22031 20096
rect 21541 19954 21607 19957
rect 12390 19952 21607 19954
rect 12390 19896 21546 19952
rect 21602 19896 21607 19952
rect 12390 19894 21607 19896
rect 0 19864 160 19894
rect 841 19891 907 19894
rect 21541 19891 21607 19894
rect 22277 19954 22343 19957
rect 22502 19954 22508 19956
rect 22277 19952 22508 19954
rect 22277 19896 22282 19952
rect 22338 19896 22508 19952
rect 22277 19894 22508 19896
rect 22277 19891 22343 19894
rect 22502 19892 22508 19894
rect 22572 19892 22578 19956
rect 1577 19818 1643 19821
rect 3049 19818 3115 19821
rect 6821 19818 6887 19821
rect 1577 19816 6887 19818
rect 1577 19760 1582 19816
rect 1638 19760 3054 19816
rect 3110 19760 6826 19816
rect 6882 19760 6887 19816
rect 1577 19758 6887 19760
rect 1577 19755 1643 19758
rect 3049 19755 3115 19758
rect 6821 19755 6887 19758
rect 7741 19818 7807 19821
rect 12709 19818 12775 19821
rect 22737 19820 22803 19821
rect 7741 19816 12775 19818
rect 7741 19760 7746 19816
rect 7802 19760 12714 19816
rect 12770 19760 12775 19816
rect 7741 19758 12775 19760
rect 7741 19755 7807 19758
rect 12709 19755 12775 19758
rect 22686 19756 22692 19820
rect 22756 19818 22803 19820
rect 22756 19816 22848 19818
rect 22798 19760 22848 19816
rect 22756 19758 22848 19760
rect 22756 19756 22803 19758
rect 22737 19755 22803 19756
rect 0 19682 160 19712
rect 1301 19682 1367 19685
rect 0 19680 1367 19682
rect 0 19624 1306 19680
rect 1362 19624 1367 19680
rect 0 19622 1367 19624
rect 0 19592 160 19622
rect 1301 19619 1367 19622
rect 10358 19620 10364 19684
rect 10428 19620 10434 19684
rect 25497 19682 25563 19685
rect 25840 19682 26000 19712
rect 25497 19680 26000 19682
rect 25497 19624 25502 19680
rect 25558 19624 26000 19680
rect 25497 19622 26000 19624
rect 6880 19616 7196 19617
rect 6880 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7196 19616
rect 6880 19551 7196 19552
rect 0 19410 160 19440
rect 10366 19413 10426 19620
rect 25497 19619 25563 19622
rect 12814 19616 13130 19617
rect 12814 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13130 19616
rect 12814 19551 13130 19552
rect 18748 19616 19064 19617
rect 18748 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19064 19616
rect 18748 19551 19064 19552
rect 24682 19616 24998 19617
rect 24682 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 24998 19616
rect 25840 19592 26000 19622
rect 24682 19551 24998 19552
rect 1761 19410 1827 19413
rect 0 19408 1827 19410
rect 0 19352 1766 19408
rect 1822 19352 1827 19408
rect 0 19350 1827 19352
rect 0 19320 160 19350
rect 1761 19347 1827 19350
rect 1945 19410 2011 19413
rect 8201 19410 8267 19413
rect 10317 19410 10426 19413
rect 13537 19410 13603 19413
rect 1945 19408 9690 19410
rect 1945 19352 1950 19408
rect 2006 19352 8206 19408
rect 8262 19352 9690 19408
rect 1945 19350 9690 19352
rect 10236 19408 13603 19410
rect 10236 19352 10322 19408
rect 10378 19352 13542 19408
rect 13598 19352 13603 19408
rect 10236 19350 13603 19352
rect 1945 19347 2011 19350
rect 8201 19347 8267 19350
rect 1669 19274 1735 19277
rect 5349 19274 5415 19277
rect 5993 19274 6059 19277
rect 1669 19272 6059 19274
rect 1669 19216 1674 19272
rect 1730 19216 5354 19272
rect 5410 19216 5998 19272
rect 6054 19216 6059 19272
rect 1669 19214 6059 19216
rect 1669 19211 1735 19214
rect 5349 19211 5415 19214
rect 5993 19211 6059 19214
rect 0 19138 160 19168
rect 3325 19138 3391 19141
rect 0 19136 3391 19138
rect 0 19080 3330 19136
rect 3386 19080 3391 19136
rect 0 19078 3391 19080
rect 0 19048 160 19078
rect 3325 19075 3391 19078
rect 5349 19138 5415 19141
rect 8017 19138 8083 19141
rect 5349 19136 8083 19138
rect 5349 19080 5354 19136
rect 5410 19080 8022 19136
rect 8078 19080 8083 19136
rect 5349 19078 8083 19080
rect 5349 19075 5415 19078
rect 8017 19075 8083 19078
rect 3913 19072 4229 19073
rect 3913 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4229 19072
rect 3913 19007 4229 19008
rect 0 18866 160 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 160 18806
rect 1393 18803 1459 18806
rect 2446 18804 2452 18868
rect 2516 18866 2522 18868
rect 3969 18866 4035 18869
rect 7557 18866 7623 18869
rect 2516 18864 7623 18866
rect 2516 18808 3974 18864
rect 4030 18808 7562 18864
rect 7618 18808 7623 18864
rect 2516 18806 7623 18808
rect 9630 18866 9690 19350
rect 10317 19347 10383 19350
rect 13537 19347 13603 19350
rect 23841 19138 23907 19141
rect 25840 19138 26000 19168
rect 23841 19136 26000 19138
rect 23841 19080 23846 19136
rect 23902 19080 26000 19136
rect 23841 19078 26000 19080
rect 23841 19075 23907 19078
rect 9847 19072 10163 19073
rect 9847 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10163 19072
rect 9847 19007 10163 19008
rect 15781 19072 16097 19073
rect 15781 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16097 19072
rect 15781 19007 16097 19008
rect 21715 19072 22031 19073
rect 21715 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22031 19072
rect 25840 19048 26000 19078
rect 21715 19007 22031 19008
rect 11605 19004 11671 19005
rect 17125 19004 17191 19005
rect 11605 19002 11652 19004
rect 11560 19000 11652 19002
rect 11560 18944 11610 19000
rect 11560 18942 11652 18944
rect 11605 18940 11652 18942
rect 11716 18940 11722 19004
rect 17125 19002 17172 19004
rect 17080 19000 17172 19002
rect 17080 18944 17130 19000
rect 17080 18942 17172 18944
rect 17125 18940 17172 18942
rect 17236 18940 17242 19004
rect 11605 18939 11671 18940
rect 17125 18939 17191 18940
rect 9857 18866 9923 18869
rect 9630 18864 9923 18866
rect 9630 18808 9862 18864
rect 9918 18808 9923 18864
rect 9630 18806 9923 18808
rect 2516 18804 2522 18806
rect 3969 18803 4035 18806
rect 7557 18803 7623 18806
rect 9857 18803 9923 18806
rect 11881 18866 11947 18869
rect 17033 18866 17099 18869
rect 11881 18864 17099 18866
rect 11881 18808 11886 18864
rect 11942 18808 17038 18864
rect 17094 18808 17099 18864
rect 11881 18806 17099 18808
rect 11881 18803 11947 18806
rect 17033 18803 17099 18806
rect 10593 18730 10659 18733
rect 13629 18732 13695 18733
rect 13629 18730 13676 18732
rect 10593 18728 13676 18730
rect 13740 18730 13746 18732
rect 10593 18672 10598 18728
rect 10654 18672 13634 18728
rect 10593 18670 13676 18672
rect 10593 18667 10659 18670
rect 13629 18668 13676 18670
rect 13740 18670 13786 18730
rect 13740 18668 13746 18670
rect 13629 18667 13695 18668
rect 0 18594 160 18624
rect 1485 18594 1551 18597
rect 0 18592 1551 18594
rect 0 18536 1490 18592
rect 1546 18536 1551 18592
rect 0 18534 1551 18536
rect 0 18504 160 18534
rect 1485 18531 1551 18534
rect 8661 18594 8727 18597
rect 10041 18594 10107 18597
rect 8661 18592 10107 18594
rect 8661 18536 8666 18592
rect 8722 18536 10046 18592
rect 10102 18536 10107 18592
rect 8661 18534 10107 18536
rect 8661 18531 8727 18534
rect 10041 18531 10107 18534
rect 25129 18594 25195 18597
rect 25840 18594 26000 18624
rect 25129 18592 26000 18594
rect 25129 18536 25134 18592
rect 25190 18536 26000 18592
rect 25129 18534 26000 18536
rect 25129 18531 25195 18534
rect 6880 18528 7196 18529
rect 6880 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7196 18528
rect 6880 18463 7196 18464
rect 12814 18528 13130 18529
rect 12814 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13130 18528
rect 12814 18463 13130 18464
rect 18748 18528 19064 18529
rect 18748 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19064 18528
rect 18748 18463 19064 18464
rect 24682 18528 24998 18529
rect 24682 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 24998 18528
rect 25840 18504 26000 18534
rect 24682 18463 24998 18464
rect 2589 18460 2655 18461
rect 2589 18458 2636 18460
rect 2508 18456 2636 18458
rect 2700 18458 2706 18460
rect 4153 18458 4219 18461
rect 5349 18460 5415 18461
rect 5349 18458 5396 18460
rect 2700 18456 4219 18458
rect 2508 18400 2594 18456
rect 2700 18400 4158 18456
rect 4214 18400 4219 18456
rect 2508 18398 2636 18400
rect 2589 18396 2636 18398
rect 2700 18398 4219 18400
rect 5304 18456 5396 18458
rect 5304 18400 5354 18456
rect 5304 18398 5396 18400
rect 2700 18396 2706 18398
rect 2589 18395 2655 18396
rect 4153 18395 4219 18398
rect 5349 18396 5396 18398
rect 5460 18396 5466 18460
rect 5349 18395 5415 18396
rect 0 18322 160 18352
rect 1301 18322 1367 18325
rect 0 18320 1367 18322
rect 0 18264 1306 18320
rect 1362 18264 1367 18320
rect 0 18262 1367 18264
rect 0 18232 160 18262
rect 1301 18259 1367 18262
rect 2589 18322 2655 18325
rect 6361 18322 6427 18325
rect 2589 18320 6427 18322
rect 2589 18264 2594 18320
rect 2650 18264 6366 18320
rect 6422 18264 6427 18320
rect 2589 18262 6427 18264
rect 2589 18259 2655 18262
rect 6361 18259 6427 18262
rect 6729 18322 6795 18325
rect 9489 18322 9555 18325
rect 6729 18320 9555 18322
rect 6729 18264 6734 18320
rect 6790 18264 9494 18320
rect 9550 18264 9555 18320
rect 6729 18262 9555 18264
rect 6729 18259 6795 18262
rect 9489 18259 9555 18262
rect 11789 18322 11855 18325
rect 21633 18322 21699 18325
rect 11789 18320 21699 18322
rect 11789 18264 11794 18320
rect 11850 18264 21638 18320
rect 21694 18264 21699 18320
rect 11789 18262 21699 18264
rect 11789 18259 11855 18262
rect 21633 18259 21699 18262
rect 3969 18186 4035 18189
rect 3969 18184 4354 18186
rect 3969 18128 3974 18184
rect 4030 18128 4354 18184
rect 3969 18126 4354 18128
rect 3969 18123 4035 18126
rect 0 18050 160 18080
rect 1209 18050 1275 18053
rect 0 18048 1275 18050
rect 0 17992 1214 18048
rect 1270 17992 1275 18048
rect 0 17990 1275 17992
rect 4294 18050 4354 18126
rect 4838 18124 4844 18188
rect 4908 18186 4914 18188
rect 4981 18186 5047 18189
rect 4908 18184 5047 18186
rect 4908 18128 4986 18184
rect 5042 18128 5047 18184
rect 4908 18126 5047 18128
rect 4908 18124 4914 18126
rect 4981 18123 5047 18126
rect 16982 18124 16988 18188
rect 17052 18186 17058 18188
rect 20846 18186 20852 18188
rect 17052 18126 20852 18186
rect 17052 18124 17058 18126
rect 20846 18124 20852 18126
rect 20916 18124 20922 18188
rect 8293 18050 8359 18053
rect 4294 18048 8359 18050
rect 4294 17992 8298 18048
rect 8354 17992 8359 18048
rect 4294 17990 8359 17992
rect 0 17960 160 17990
rect 1209 17987 1275 17990
rect 8293 17987 8359 17990
rect 14590 17988 14596 18052
rect 14660 18050 14666 18052
rect 15510 18050 15516 18052
rect 14660 17990 15516 18050
rect 14660 17988 14666 17990
rect 15510 17988 15516 17990
rect 15580 17988 15586 18052
rect 20713 18050 20779 18053
rect 20846 18050 20852 18052
rect 20713 18048 20852 18050
rect 20713 17992 20718 18048
rect 20774 17992 20852 18048
rect 20713 17990 20852 17992
rect 20713 17987 20779 17990
rect 20846 17988 20852 17990
rect 20916 17988 20922 18052
rect 24393 18050 24459 18053
rect 25840 18050 26000 18080
rect 24393 18048 26000 18050
rect 24393 17992 24398 18048
rect 24454 17992 26000 18048
rect 24393 17990 26000 17992
rect 24393 17987 24459 17990
rect 3913 17984 4229 17985
rect 3913 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4229 17984
rect 3913 17919 4229 17920
rect 9847 17984 10163 17985
rect 9847 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10163 17984
rect 9847 17919 10163 17920
rect 15781 17984 16097 17985
rect 15781 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16097 17984
rect 15781 17919 16097 17920
rect 21715 17984 22031 17985
rect 21715 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22031 17984
rect 25840 17960 26000 17990
rect 21715 17919 22031 17920
rect 10726 17852 10732 17916
rect 10796 17852 10802 17916
rect 12014 17852 12020 17916
rect 12084 17914 12090 17916
rect 12433 17914 12499 17917
rect 12084 17912 12499 17914
rect 12084 17856 12438 17912
rect 12494 17856 12499 17912
rect 12084 17854 12499 17856
rect 12084 17852 12090 17854
rect 0 17778 160 17808
rect 1577 17778 1643 17781
rect 3969 17778 4035 17781
rect 5993 17778 6059 17781
rect 10734 17778 10794 17852
rect 12433 17851 12499 17854
rect 13353 17914 13419 17917
rect 16849 17914 16915 17917
rect 19742 17914 19748 17916
rect 13353 17912 13738 17914
rect 13353 17856 13358 17912
rect 13414 17856 13738 17912
rect 13353 17854 13738 17856
rect 13353 17851 13419 17854
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 160 17718
rect 1577 17715 1643 17718
rect 2730 17776 10794 17778
rect 2730 17720 3974 17776
rect 4030 17720 5998 17776
rect 6054 17720 10794 17776
rect 2730 17718 10794 17720
rect 0 17506 160 17536
rect 1761 17506 1827 17509
rect 0 17504 1827 17506
rect 0 17448 1766 17504
rect 1822 17448 1827 17504
rect 0 17446 1827 17448
rect 0 17416 160 17446
rect 1761 17443 1827 17446
rect 2078 17308 2084 17372
rect 2148 17370 2154 17372
rect 2730 17370 2790 17718
rect 3969 17715 4035 17718
rect 5993 17715 6059 17718
rect 13678 17642 13738 17854
rect 16849 17912 19748 17914
rect 16849 17856 16854 17912
rect 16910 17856 19748 17912
rect 16849 17854 19748 17856
rect 16849 17851 16915 17854
rect 19742 17852 19748 17854
rect 19812 17852 19818 17916
rect 17718 17716 17724 17780
rect 17788 17778 17794 17780
rect 22277 17778 22343 17781
rect 17788 17776 22343 17778
rect 17788 17720 22282 17776
rect 22338 17720 22343 17776
rect 17788 17718 22343 17720
rect 17788 17716 17794 17718
rect 22277 17715 22343 17718
rect 13678 17582 23122 17642
rect 21214 17444 21220 17508
rect 21284 17506 21290 17508
rect 21541 17506 21607 17509
rect 21284 17504 21607 17506
rect 21284 17448 21546 17504
rect 21602 17448 21607 17504
rect 21284 17446 21607 17448
rect 21284 17444 21290 17446
rect 21541 17443 21607 17446
rect 6880 17440 7196 17441
rect 6880 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7196 17440
rect 6880 17375 7196 17376
rect 12814 17440 13130 17441
rect 12814 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13130 17440
rect 12814 17375 13130 17376
rect 18748 17440 19064 17441
rect 18748 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19064 17440
rect 18748 17375 19064 17376
rect 2148 17310 2790 17370
rect 2148 17308 2154 17310
rect 0 17234 160 17264
rect 23062 17237 23122 17582
rect 25129 17506 25195 17509
rect 25840 17506 26000 17536
rect 25129 17504 26000 17506
rect 25129 17448 25134 17504
rect 25190 17448 26000 17504
rect 25129 17446 26000 17448
rect 25129 17443 25195 17446
rect 24682 17440 24998 17441
rect 24682 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 24998 17440
rect 25840 17416 26000 17446
rect 24682 17375 24998 17376
rect 3325 17234 3391 17237
rect 0 17232 3391 17234
rect 0 17176 3330 17232
rect 3386 17176 3391 17232
rect 0 17174 3391 17176
rect 0 17144 160 17174
rect 3325 17171 3391 17174
rect 6545 17234 6611 17237
rect 12249 17234 12315 17237
rect 6545 17232 22110 17234
rect 6545 17176 6550 17232
rect 6606 17176 12254 17232
rect 12310 17176 22110 17232
rect 6545 17174 22110 17176
rect 6545 17171 6611 17174
rect 12249 17171 12315 17174
rect 1025 17098 1091 17101
rect 6913 17098 6979 17101
rect 1025 17096 6979 17098
rect 1025 17040 1030 17096
rect 1086 17040 6918 17096
rect 6974 17040 6979 17096
rect 1025 17038 6979 17040
rect 1025 17035 1091 17038
rect 6913 17035 6979 17038
rect 10409 17098 10475 17101
rect 14457 17098 14523 17101
rect 17861 17098 17927 17101
rect 10409 17096 17927 17098
rect 10409 17040 10414 17096
rect 10470 17040 14462 17096
rect 14518 17040 17866 17096
rect 17922 17040 17927 17096
rect 10409 17038 17927 17040
rect 22050 17098 22110 17174
rect 23013 17232 23122 17237
rect 25865 17234 25931 17237
rect 23013 17176 23018 17232
rect 23074 17176 23122 17232
rect 23013 17174 23122 17176
rect 23982 17232 25931 17234
rect 23982 17176 25870 17232
rect 25926 17176 25931 17232
rect 23982 17174 25931 17176
rect 23013 17171 23079 17174
rect 23982 17098 24042 17174
rect 25865 17171 25931 17174
rect 22050 17038 24042 17098
rect 10409 17035 10475 17038
rect 14457 17035 14523 17038
rect 17861 17035 17927 17038
rect 0 16962 160 16992
rect 1025 16962 1091 16965
rect 0 16960 1091 16962
rect 0 16904 1030 16960
rect 1086 16904 1091 16960
rect 0 16902 1091 16904
rect 0 16872 160 16902
rect 1025 16899 1091 16902
rect 5165 16962 5231 16965
rect 7465 16962 7531 16965
rect 5165 16960 7531 16962
rect 5165 16904 5170 16960
rect 5226 16904 7470 16960
rect 7526 16904 7531 16960
rect 5165 16902 7531 16904
rect 5165 16899 5231 16902
rect 7465 16899 7531 16902
rect 24117 16962 24183 16965
rect 25840 16962 26000 16992
rect 24117 16960 26000 16962
rect 24117 16904 24122 16960
rect 24178 16904 26000 16960
rect 24117 16902 26000 16904
rect 24117 16899 24183 16902
rect 3913 16896 4229 16897
rect 3913 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4229 16896
rect 3913 16831 4229 16832
rect 9847 16896 10163 16897
rect 9847 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10163 16896
rect 9847 16831 10163 16832
rect 15781 16896 16097 16897
rect 15781 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16097 16896
rect 15781 16831 16097 16832
rect 21715 16896 22031 16897
rect 21715 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22031 16896
rect 25840 16872 26000 16902
rect 21715 16831 22031 16832
rect 1853 16828 1919 16829
rect 1853 16826 1900 16828
rect 1808 16824 1900 16826
rect 1808 16768 1858 16824
rect 1808 16766 1900 16768
rect 1853 16764 1900 16766
rect 1964 16764 1970 16828
rect 1853 16763 1919 16764
rect 0 16690 160 16720
rect 2865 16690 2931 16693
rect 0 16688 2931 16690
rect 0 16632 2870 16688
rect 2926 16632 2931 16688
rect 0 16630 2931 16632
rect 0 16600 160 16630
rect 2865 16627 2931 16630
rect 7373 16554 7439 16557
rect 7966 16554 7972 16556
rect 7373 16552 7972 16554
rect 7373 16496 7378 16552
rect 7434 16496 7972 16552
rect 7373 16494 7972 16496
rect 7373 16491 7439 16494
rect 7966 16492 7972 16494
rect 8036 16492 8042 16556
rect 9765 16554 9831 16557
rect 15469 16554 15535 16557
rect 9765 16552 15535 16554
rect 9765 16496 9770 16552
rect 9826 16496 15474 16552
rect 15530 16496 15535 16552
rect 9765 16494 15535 16496
rect 9765 16491 9831 16494
rect 15469 16491 15535 16494
rect 23933 16554 23999 16557
rect 23933 16552 25146 16554
rect 23933 16496 23938 16552
rect 23994 16496 25146 16552
rect 23933 16494 25146 16496
rect 23933 16491 23999 16494
rect 0 16418 160 16448
rect 2681 16418 2747 16421
rect 0 16416 2747 16418
rect 0 16360 2686 16416
rect 2742 16360 2747 16416
rect 0 16358 2747 16360
rect 0 16328 160 16358
rect 2681 16355 2747 16358
rect 19977 16418 20043 16421
rect 20294 16418 20300 16420
rect 19977 16416 20300 16418
rect 19977 16360 19982 16416
rect 20038 16360 20300 16416
rect 19977 16358 20300 16360
rect 19977 16355 20043 16358
rect 20294 16356 20300 16358
rect 20364 16356 20370 16420
rect 25086 16418 25146 16494
rect 25840 16418 26000 16448
rect 25086 16358 26000 16418
rect 6880 16352 7196 16353
rect 6880 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7196 16352
rect 6880 16287 7196 16288
rect 12814 16352 13130 16353
rect 12814 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13130 16352
rect 12814 16287 13130 16288
rect 18748 16352 19064 16353
rect 18748 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19064 16352
rect 18748 16287 19064 16288
rect 24682 16352 24998 16353
rect 24682 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 24998 16352
rect 25840 16328 26000 16358
rect 24682 16287 24998 16288
rect 3325 16282 3391 16285
rect 3550 16282 3556 16284
rect 3325 16280 3556 16282
rect 3325 16224 3330 16280
rect 3386 16224 3556 16280
rect 3325 16222 3556 16224
rect 3325 16219 3391 16222
rect 3550 16220 3556 16222
rect 3620 16220 3626 16284
rect 0 16146 160 16176
rect 3049 16146 3115 16149
rect 0 16144 3115 16146
rect 0 16088 3054 16144
rect 3110 16088 3115 16144
rect 0 16086 3115 16088
rect 0 16056 160 16086
rect 3049 16083 3115 16086
rect 4337 16146 4403 16149
rect 6177 16146 6243 16149
rect 7833 16146 7899 16149
rect 4337 16144 7899 16146
rect 4337 16088 4342 16144
rect 4398 16088 6182 16144
rect 6238 16088 7838 16144
rect 7894 16088 7899 16144
rect 4337 16086 7899 16088
rect 4337 16083 4403 16086
rect 6177 16083 6243 16086
rect 7833 16083 7899 16086
rect 15510 15948 15516 16012
rect 15580 16010 15586 16012
rect 15837 16010 15903 16013
rect 15580 16008 15903 16010
rect 15580 15952 15842 16008
rect 15898 15952 15903 16008
rect 15580 15950 15903 15952
rect 15580 15948 15586 15950
rect 15837 15947 15903 15950
rect 0 15874 160 15904
rect 1669 15874 1735 15877
rect 0 15872 1735 15874
rect 0 15816 1674 15872
rect 1730 15816 1735 15872
rect 0 15814 1735 15816
rect 0 15784 160 15814
rect 1669 15811 1735 15814
rect 24117 15874 24183 15877
rect 25840 15874 26000 15904
rect 24117 15872 26000 15874
rect 24117 15816 24122 15872
rect 24178 15816 26000 15872
rect 24117 15814 26000 15816
rect 24117 15811 24183 15814
rect 3913 15808 4229 15809
rect 3913 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4229 15808
rect 3913 15743 4229 15744
rect 9847 15808 10163 15809
rect 9847 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10163 15808
rect 9847 15743 10163 15744
rect 15781 15808 16097 15809
rect 15781 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16097 15808
rect 15781 15743 16097 15744
rect 21715 15808 22031 15809
rect 21715 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22031 15808
rect 25840 15784 26000 15814
rect 21715 15743 22031 15744
rect 0 15602 160 15632
rect 3049 15602 3115 15605
rect 0 15600 3115 15602
rect 0 15544 3054 15600
rect 3110 15544 3115 15600
rect 0 15542 3115 15544
rect 0 15512 160 15542
rect 3049 15539 3115 15542
rect 3366 15540 3372 15604
rect 3436 15602 3442 15604
rect 3509 15602 3575 15605
rect 3436 15600 3575 15602
rect 3436 15544 3514 15600
rect 3570 15544 3575 15600
rect 3436 15542 3575 15544
rect 3436 15540 3442 15542
rect 3509 15539 3575 15542
rect 9857 15602 9923 15605
rect 15193 15602 15259 15605
rect 9857 15600 15259 15602
rect 9857 15544 9862 15600
rect 9918 15544 15198 15600
rect 15254 15544 15259 15600
rect 9857 15542 15259 15544
rect 9857 15539 9923 15542
rect 15193 15539 15259 15542
rect 3969 15466 4035 15469
rect 1396 15464 4035 15466
rect 1396 15408 3974 15464
rect 4030 15408 4035 15464
rect 1396 15406 4035 15408
rect 0 15330 160 15360
rect 1396 15330 1456 15406
rect 3969 15403 4035 15406
rect 12249 15466 12315 15469
rect 14406 15466 14412 15468
rect 12249 15464 14412 15466
rect 12249 15408 12254 15464
rect 12310 15408 14412 15464
rect 12249 15406 14412 15408
rect 12249 15403 12315 15406
rect 14406 15404 14412 15406
rect 14476 15404 14482 15468
rect 0 15270 1456 15330
rect 25497 15330 25563 15333
rect 25840 15330 26000 15360
rect 25497 15328 26000 15330
rect 25497 15272 25502 15328
rect 25558 15272 26000 15328
rect 25497 15270 26000 15272
rect 0 15240 160 15270
rect 25497 15267 25563 15270
rect 6880 15264 7196 15265
rect 6880 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7196 15264
rect 6880 15199 7196 15200
rect 12814 15264 13130 15265
rect 12814 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13130 15264
rect 12814 15199 13130 15200
rect 18748 15264 19064 15265
rect 18748 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19064 15264
rect 18748 15199 19064 15200
rect 24682 15264 24998 15265
rect 24682 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 24998 15264
rect 25840 15240 26000 15270
rect 24682 15199 24998 15200
rect 2313 15194 2379 15197
rect 4613 15196 4679 15197
rect 4613 15194 4660 15196
rect 1166 15192 2379 15194
rect 1166 15136 2318 15192
rect 2374 15136 2379 15192
rect 1166 15134 2379 15136
rect 4568 15192 4660 15194
rect 4568 15136 4618 15192
rect 4568 15134 4660 15136
rect 0 15058 160 15088
rect 1166 15058 1226 15134
rect 2313 15131 2379 15134
rect 4613 15132 4660 15134
rect 4724 15132 4730 15196
rect 11513 15194 11579 15197
rect 16205 15196 16271 15197
rect 11646 15194 11652 15196
rect 11513 15192 11652 15194
rect 11513 15136 11518 15192
rect 11574 15136 11652 15192
rect 11513 15134 11652 15136
rect 4613 15131 4679 15132
rect 11513 15131 11579 15134
rect 11646 15132 11652 15134
rect 11716 15132 11722 15196
rect 16205 15194 16252 15196
rect 16160 15192 16252 15194
rect 16160 15136 16210 15192
rect 16160 15134 16252 15136
rect 16205 15132 16252 15134
rect 16316 15132 16322 15196
rect 16205 15131 16271 15132
rect 0 14998 1226 15058
rect 6545 15058 6611 15061
rect 6821 15058 6887 15061
rect 6545 15056 6887 15058
rect 6545 15000 6550 15056
rect 6606 15000 6826 15056
rect 6882 15000 6887 15056
rect 6545 14998 6887 15000
rect 0 14968 160 14998
rect 6545 14995 6611 14998
rect 6821 14995 6887 14998
rect 17493 15058 17559 15061
rect 20621 15058 20687 15061
rect 17493 15056 20687 15058
rect 17493 15000 17498 15056
rect 17554 15000 20626 15056
rect 20682 15000 20687 15056
rect 17493 14998 20687 15000
rect 17493 14995 17559 14998
rect 20621 14995 20687 14998
rect 10869 14922 10935 14925
rect 20897 14922 20963 14925
rect 10869 14920 20963 14922
rect 10869 14864 10874 14920
rect 10930 14864 20902 14920
rect 20958 14864 20963 14920
rect 10869 14862 20963 14864
rect 10869 14859 10935 14862
rect 20897 14859 20963 14862
rect 0 14786 160 14816
rect 5809 14786 5875 14789
rect 5942 14786 5948 14788
rect 0 14726 858 14786
rect 0 14696 160 14726
rect 798 14650 858 14726
rect 5809 14784 5948 14786
rect 5809 14728 5814 14784
rect 5870 14728 5948 14784
rect 5809 14726 5948 14728
rect 5809 14723 5875 14726
rect 5942 14724 5948 14726
rect 6012 14724 6018 14788
rect 24025 14786 24091 14789
rect 25840 14786 26000 14816
rect 24025 14784 26000 14786
rect 24025 14728 24030 14784
rect 24086 14728 26000 14784
rect 24025 14726 26000 14728
rect 24025 14723 24091 14726
rect 3913 14720 4229 14721
rect 3913 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4229 14720
rect 3913 14655 4229 14656
rect 9847 14720 10163 14721
rect 9847 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10163 14720
rect 9847 14655 10163 14656
rect 15781 14720 16097 14721
rect 15781 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16097 14720
rect 15781 14655 16097 14656
rect 21715 14720 22031 14721
rect 21715 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22031 14720
rect 25840 14696 26000 14726
rect 21715 14655 22031 14656
rect 1853 14650 1919 14653
rect 798 14648 1919 14650
rect 798 14592 1858 14648
rect 1914 14592 1919 14648
rect 798 14590 1919 14592
rect 1853 14587 1919 14590
rect 5625 14650 5691 14653
rect 6126 14650 6132 14652
rect 5625 14648 6132 14650
rect 5625 14592 5630 14648
rect 5686 14592 6132 14648
rect 5625 14590 6132 14592
rect 5625 14587 5691 14590
rect 6126 14588 6132 14590
rect 6196 14588 6202 14652
rect 10961 14650 11027 14653
rect 14273 14650 14339 14653
rect 10961 14648 14339 14650
rect 10961 14592 10966 14648
rect 11022 14592 14278 14648
rect 14334 14592 14339 14648
rect 10961 14590 14339 14592
rect 10961 14587 11027 14590
rect 14273 14587 14339 14590
rect 0 14514 160 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 160 14454
rect 2773 14451 2839 14454
rect 4245 14514 4311 14517
rect 17769 14514 17835 14517
rect 4245 14512 17835 14514
rect 4245 14456 4250 14512
rect 4306 14456 17774 14512
rect 17830 14456 17835 14512
rect 4245 14454 17835 14456
rect 4245 14451 4311 14454
rect 17769 14451 17835 14454
rect 1761 14378 1827 14381
rect 5349 14378 5415 14381
rect 6821 14378 6887 14381
rect 1761 14376 5415 14378
rect 1761 14320 1766 14376
rect 1822 14320 5354 14376
rect 5410 14320 5415 14376
rect 1761 14318 5415 14320
rect 1761 14315 1827 14318
rect 5349 14315 5415 14318
rect 5582 14376 6887 14378
rect 5582 14320 6826 14376
rect 6882 14320 6887 14376
rect 5582 14318 6887 14320
rect 0 14242 160 14272
rect 1761 14242 1827 14245
rect 0 14240 1827 14242
rect 0 14184 1766 14240
rect 1822 14184 1827 14240
rect 0 14182 1827 14184
rect 0 14152 160 14182
rect 1761 14179 1827 14182
rect 1945 14242 2011 14245
rect 5582 14242 5642 14318
rect 6821 14315 6887 14318
rect 11881 14378 11947 14381
rect 16113 14378 16179 14381
rect 11881 14376 16179 14378
rect 11881 14320 11886 14376
rect 11942 14320 16118 14376
rect 16174 14320 16179 14376
rect 11881 14318 16179 14320
rect 11881 14315 11947 14318
rect 16113 14315 16179 14318
rect 1945 14240 5642 14242
rect 1945 14184 1950 14240
rect 2006 14184 5642 14240
rect 1945 14182 5642 14184
rect 25129 14242 25195 14245
rect 25840 14242 26000 14272
rect 25129 14240 26000 14242
rect 25129 14184 25134 14240
rect 25190 14184 26000 14240
rect 25129 14182 26000 14184
rect 1945 14179 2011 14182
rect 25129 14179 25195 14182
rect 6880 14176 7196 14177
rect 6880 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7196 14176
rect 6880 14111 7196 14112
rect 12814 14176 13130 14177
rect 12814 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13130 14176
rect 12814 14111 13130 14112
rect 18748 14176 19064 14177
rect 18748 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19064 14176
rect 18748 14111 19064 14112
rect 24682 14176 24998 14177
rect 24682 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 24998 14176
rect 25840 14152 26000 14182
rect 24682 14111 24998 14112
rect 5441 14106 5507 14109
rect 5901 14106 5967 14109
rect 5441 14104 5967 14106
rect 5441 14048 5446 14104
rect 5502 14048 5906 14104
rect 5962 14048 5967 14104
rect 5441 14046 5967 14048
rect 5441 14043 5507 14046
rect 5901 14043 5967 14046
rect 0 13970 160 14000
rect 1393 13970 1459 13973
rect 0 13968 1459 13970
rect 0 13912 1398 13968
rect 1454 13912 1459 13968
rect 0 13910 1459 13912
rect 0 13880 160 13910
rect 1393 13907 1459 13910
rect 5390 13908 5396 13972
rect 5460 13970 5466 13972
rect 5625 13970 5691 13973
rect 5460 13968 5691 13970
rect 5460 13912 5630 13968
rect 5686 13912 5691 13968
rect 5460 13910 5691 13912
rect 5460 13908 5466 13910
rect 5625 13907 5691 13910
rect 11605 13970 11671 13973
rect 14917 13970 14983 13973
rect 11605 13968 14983 13970
rect 11605 13912 11610 13968
rect 11666 13912 14922 13968
rect 14978 13912 14983 13968
rect 11605 13910 14983 13912
rect 11605 13907 11671 13910
rect 14917 13907 14983 13910
rect 12157 13834 12223 13837
rect 16941 13834 17007 13837
rect 12157 13832 17007 13834
rect 12157 13776 12162 13832
rect 12218 13776 16946 13832
rect 17002 13776 17007 13832
rect 12157 13774 17007 13776
rect 12157 13771 12223 13774
rect 16941 13771 17007 13774
rect 0 13698 160 13728
rect 3785 13698 3851 13701
rect 0 13696 3851 13698
rect 0 13640 3790 13696
rect 3846 13640 3851 13696
rect 0 13638 3851 13640
rect 0 13608 160 13638
rect 3785 13635 3851 13638
rect 10593 13698 10659 13701
rect 10910 13698 10916 13700
rect 10593 13696 10916 13698
rect 10593 13640 10598 13696
rect 10654 13640 10916 13696
rect 10593 13638 10916 13640
rect 10593 13635 10659 13638
rect 10910 13636 10916 13638
rect 10980 13636 10986 13700
rect 22185 13698 22251 13701
rect 22318 13698 22324 13700
rect 22185 13696 22324 13698
rect 22185 13640 22190 13696
rect 22246 13640 22324 13696
rect 22185 13638 22324 13640
rect 22185 13635 22251 13638
rect 22318 13636 22324 13638
rect 22388 13636 22394 13700
rect 24393 13698 24459 13701
rect 25840 13698 26000 13728
rect 24393 13696 26000 13698
rect 24393 13640 24398 13696
rect 24454 13640 26000 13696
rect 24393 13638 26000 13640
rect 24393 13635 24459 13638
rect 3913 13632 4229 13633
rect 3913 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4229 13632
rect 3913 13567 4229 13568
rect 9847 13632 10163 13633
rect 9847 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10163 13632
rect 9847 13567 10163 13568
rect 15781 13632 16097 13633
rect 15781 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16097 13632
rect 15781 13567 16097 13568
rect 21715 13632 22031 13633
rect 21715 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22031 13632
rect 25840 13608 26000 13638
rect 21715 13567 22031 13568
rect 5901 13564 5967 13565
rect 5901 13562 5948 13564
rect 5856 13560 5948 13562
rect 5856 13504 5906 13560
rect 5856 13502 5948 13504
rect 5901 13500 5948 13502
rect 6012 13500 6018 13564
rect 5901 13499 5967 13500
rect 0 13426 160 13456
rect 3785 13426 3851 13429
rect 4797 13426 4863 13429
rect 6085 13426 6151 13429
rect 6637 13426 6703 13429
rect 0 13366 1410 13426
rect 0 13336 160 13366
rect 0 13154 160 13184
rect 1209 13154 1275 13157
rect 0 13152 1275 13154
rect 0 13096 1214 13152
rect 1270 13096 1275 13152
rect 0 13094 1275 13096
rect 0 13064 160 13094
rect 1209 13091 1275 13094
rect 1350 13018 1410 13366
rect 3785 13424 6703 13426
rect 3785 13368 3790 13424
rect 3846 13368 4802 13424
rect 4858 13368 6090 13424
rect 6146 13368 6642 13424
rect 6698 13368 6703 13424
rect 3785 13366 6703 13368
rect 3785 13363 3851 13366
rect 4797 13363 4863 13366
rect 6085 13363 6151 13366
rect 6637 13363 6703 13366
rect 19517 13426 19583 13429
rect 23473 13426 23539 13429
rect 19517 13424 23539 13426
rect 19517 13368 19522 13424
rect 19578 13368 23478 13424
rect 23534 13368 23539 13424
rect 19517 13366 23539 13368
rect 19517 13363 19583 13366
rect 23473 13363 23539 13366
rect 3325 13290 3391 13293
rect 3550 13290 3556 13292
rect 3325 13288 3556 13290
rect 3325 13232 3330 13288
rect 3386 13232 3556 13288
rect 3325 13230 3556 13232
rect 3325 13227 3391 13230
rect 3550 13228 3556 13230
rect 3620 13290 3626 13292
rect 4061 13290 4127 13293
rect 12433 13292 12499 13293
rect 12382 13290 12388 13292
rect 3620 13288 4127 13290
rect 3620 13232 4066 13288
rect 4122 13232 4127 13288
rect 3620 13230 4127 13232
rect 12346 13230 12388 13290
rect 12452 13290 12499 13292
rect 12452 13288 12544 13290
rect 12494 13232 12544 13288
rect 3620 13228 3626 13230
rect 4061 13227 4127 13230
rect 12382 13228 12388 13230
rect 12452 13230 12544 13232
rect 12452 13228 12499 13230
rect 12433 13227 12499 13228
rect 25840 13154 26000 13184
rect 25454 13094 26000 13154
rect 6880 13088 7196 13089
rect 6880 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7196 13088
rect 6880 13023 7196 13024
rect 12814 13088 13130 13089
rect 12814 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13130 13088
rect 12814 13023 13130 13024
rect 18748 13088 19064 13089
rect 18748 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19064 13088
rect 18748 13023 19064 13024
rect 24682 13088 24998 13089
rect 24682 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 24998 13088
rect 24682 13023 24998 13024
rect 3509 13018 3575 13021
rect 1350 13016 3575 13018
rect 1350 12960 3514 13016
rect 3570 12960 3575 13016
rect 1350 12958 3575 12960
rect 3509 12955 3575 12958
rect 0 12882 160 12912
rect 2313 12882 2379 12885
rect 0 12880 2379 12882
rect 0 12824 2318 12880
rect 2374 12824 2379 12880
rect 0 12822 2379 12824
rect 0 12792 160 12822
rect 2313 12819 2379 12822
rect 3877 12882 3943 12885
rect 6269 12882 6335 12885
rect 3877 12880 6335 12882
rect 3877 12824 3882 12880
rect 3938 12824 6274 12880
rect 6330 12824 6335 12880
rect 3877 12822 6335 12824
rect 3877 12819 3943 12822
rect 6269 12819 6335 12822
rect 11237 12882 11303 12885
rect 13813 12882 13879 12885
rect 11237 12880 13879 12882
rect 11237 12824 11242 12880
rect 11298 12824 13818 12880
rect 13874 12824 13879 12880
rect 11237 12822 13879 12824
rect 11237 12819 11303 12822
rect 13813 12819 13879 12822
rect 4061 12746 4127 12749
rect 8937 12746 9003 12749
rect 4061 12744 9003 12746
rect 4061 12688 4066 12744
rect 4122 12688 8942 12744
rect 8998 12688 9003 12744
rect 4061 12686 9003 12688
rect 4061 12683 4127 12686
rect 0 12610 160 12640
rect 657 12610 723 12613
rect 0 12608 723 12610
rect 0 12552 662 12608
rect 718 12552 723 12608
rect 0 12550 723 12552
rect 0 12520 160 12550
rect 657 12547 723 12550
rect 3913 12544 4229 12545
rect 3913 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4229 12544
rect 3913 12479 4229 12480
rect 0 12338 160 12368
rect 4294 12341 4354 12686
rect 8937 12683 9003 12686
rect 10409 12746 10475 12749
rect 10542 12746 10548 12748
rect 10409 12744 10548 12746
rect 10409 12688 10414 12744
rect 10470 12688 10548 12744
rect 10409 12686 10548 12688
rect 10409 12683 10475 12686
rect 10542 12684 10548 12686
rect 10612 12684 10618 12748
rect 11646 12684 11652 12748
rect 11716 12746 11722 12748
rect 11881 12746 11947 12749
rect 11716 12744 11947 12746
rect 11716 12688 11886 12744
rect 11942 12688 11947 12744
rect 11716 12686 11947 12688
rect 11716 12684 11722 12686
rect 11881 12683 11947 12686
rect 21265 12746 21331 12749
rect 24485 12746 24551 12749
rect 21265 12744 24551 12746
rect 21265 12688 21270 12744
rect 21326 12688 24490 12744
rect 24546 12688 24551 12744
rect 21265 12686 24551 12688
rect 21265 12683 21331 12686
rect 24485 12683 24551 12686
rect 25129 12746 25195 12749
rect 25454 12746 25514 13094
rect 25840 13064 26000 13094
rect 25129 12744 25514 12746
rect 25129 12688 25134 12744
rect 25190 12688 25514 12744
rect 25129 12686 25514 12688
rect 25129 12683 25195 12686
rect 5073 12608 5139 12613
rect 5073 12552 5078 12608
rect 5134 12552 5139 12608
rect 5073 12547 5139 12552
rect 22553 12610 22619 12613
rect 23013 12610 23079 12613
rect 22553 12608 23079 12610
rect 22553 12552 22558 12608
rect 22614 12552 23018 12608
rect 23074 12552 23079 12608
rect 22553 12550 23079 12552
rect 22553 12547 22619 12550
rect 23013 12547 23079 12550
rect 24209 12610 24275 12613
rect 25840 12610 26000 12640
rect 24209 12608 26000 12610
rect 24209 12552 24214 12608
rect 24270 12552 26000 12608
rect 24209 12550 26000 12552
rect 24209 12547 24275 12550
rect 4797 12474 4863 12477
rect 5076 12474 5136 12547
rect 9847 12544 10163 12545
rect 9847 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10163 12544
rect 9847 12479 10163 12480
rect 15781 12544 16097 12545
rect 15781 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16097 12544
rect 15781 12479 16097 12480
rect 21715 12544 22031 12545
rect 21715 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22031 12544
rect 25840 12520 26000 12550
rect 21715 12479 22031 12480
rect 4797 12472 5136 12474
rect 4797 12416 4802 12472
rect 4858 12416 5136 12472
rect 4797 12414 5136 12416
rect 4797 12411 4863 12414
rect 3693 12338 3759 12341
rect 0 12336 3759 12338
rect 0 12280 3698 12336
rect 3754 12280 3759 12336
rect 0 12278 3759 12280
rect 0 12248 160 12278
rect 3693 12275 3759 12278
rect 4245 12336 4354 12341
rect 4245 12280 4250 12336
rect 4306 12280 4354 12336
rect 4245 12278 4354 12280
rect 5901 12338 5967 12341
rect 7833 12338 7899 12341
rect 5901 12336 7899 12338
rect 5901 12280 5906 12336
rect 5962 12280 7838 12336
rect 7894 12280 7899 12336
rect 5901 12278 7899 12280
rect 4245 12275 4311 12278
rect 5901 12275 5967 12278
rect 7833 12275 7899 12278
rect 21173 12340 21239 12341
rect 21173 12336 21220 12340
rect 21284 12338 21290 12340
rect 21173 12280 21178 12336
rect 21173 12276 21220 12280
rect 21284 12278 21330 12338
rect 21284 12276 21290 12278
rect 21173 12275 21239 12276
rect 2957 12202 3023 12205
rect 3366 12202 3372 12204
rect 2957 12200 3372 12202
rect 2957 12144 2962 12200
rect 3018 12144 3372 12200
rect 2957 12142 3372 12144
rect 2957 12139 3023 12142
rect 3366 12140 3372 12142
rect 3436 12202 3442 12204
rect 3877 12202 3943 12205
rect 3436 12200 3943 12202
rect 3436 12144 3882 12200
rect 3938 12144 3943 12200
rect 3436 12142 3943 12144
rect 3436 12140 3442 12142
rect 3877 12139 3943 12142
rect 0 12066 160 12096
rect 1393 12066 1459 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 160 12006
rect 1393 12003 1459 12006
rect 2865 12066 2931 12069
rect 4153 12066 4219 12069
rect 2865 12064 4219 12066
rect 2865 12008 2870 12064
rect 2926 12008 4158 12064
rect 4214 12008 4219 12064
rect 2865 12006 4219 12008
rect 2865 12003 2931 12006
rect 4153 12003 4219 12006
rect 25221 12066 25287 12069
rect 25840 12066 26000 12096
rect 25221 12064 26000 12066
rect 25221 12008 25226 12064
rect 25282 12008 26000 12064
rect 25221 12006 26000 12008
rect 25221 12003 25287 12006
rect 6880 12000 7196 12001
rect 6880 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7196 12000
rect 6880 11935 7196 11936
rect 12814 12000 13130 12001
rect 12814 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13130 12000
rect 12814 11935 13130 11936
rect 18748 12000 19064 12001
rect 18748 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19064 12000
rect 18748 11935 19064 11936
rect 24682 12000 24998 12001
rect 24682 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 24998 12000
rect 25840 11976 26000 12006
rect 24682 11935 24998 11936
rect 2773 11930 2839 11933
rect 2773 11928 6746 11930
rect 2773 11872 2778 11928
rect 2834 11872 6746 11928
rect 2773 11870 6746 11872
rect 2773 11867 2839 11870
rect 0 11794 160 11824
rect 3141 11794 3207 11797
rect 0 11792 3207 11794
rect 0 11736 3146 11792
rect 3202 11736 3207 11792
rect 0 11734 3207 11736
rect 0 11704 160 11734
rect 3141 11731 3207 11734
rect 3509 11794 3575 11797
rect 4705 11794 4771 11797
rect 3509 11792 4771 11794
rect 3509 11736 3514 11792
rect 3570 11736 4710 11792
rect 4766 11736 4771 11792
rect 3509 11734 4771 11736
rect 3509 11731 3575 11734
rect 4705 11731 4771 11734
rect 5022 11732 5028 11796
rect 5092 11794 5098 11796
rect 5257 11794 5323 11797
rect 5092 11792 5323 11794
rect 5092 11736 5262 11792
rect 5318 11736 5323 11792
rect 5092 11734 5323 11736
rect 6686 11794 6746 11870
rect 7557 11794 7623 11797
rect 6686 11792 7623 11794
rect 6686 11736 7562 11792
rect 7618 11736 7623 11792
rect 6686 11734 7623 11736
rect 5092 11732 5098 11734
rect 5257 11731 5323 11734
rect 7557 11731 7623 11734
rect 14733 11794 14799 11797
rect 19425 11794 19491 11797
rect 14733 11792 19491 11794
rect 14733 11736 14738 11792
rect 14794 11736 19430 11792
rect 19486 11736 19491 11792
rect 14733 11734 19491 11736
rect 14733 11731 14799 11734
rect 19425 11731 19491 11734
rect 3325 11658 3391 11661
rect 16573 11658 16639 11661
rect 3325 11656 16639 11658
rect 3325 11600 3330 11656
rect 3386 11600 16578 11656
rect 16634 11600 16639 11656
rect 3325 11598 16639 11600
rect 3325 11595 3391 11598
rect 16573 11595 16639 11598
rect 0 11522 160 11552
rect 1853 11522 1919 11525
rect 0 11520 1919 11522
rect 0 11464 1858 11520
rect 1914 11464 1919 11520
rect 0 11462 1919 11464
rect 0 11432 160 11462
rect 1853 11459 1919 11462
rect 3233 11522 3299 11525
rect 3601 11522 3667 11525
rect 3233 11520 3667 11522
rect 3233 11464 3238 11520
rect 3294 11464 3606 11520
rect 3662 11464 3667 11520
rect 3233 11462 3667 11464
rect 3233 11459 3299 11462
rect 3601 11459 3667 11462
rect 23841 11522 23907 11525
rect 25840 11522 26000 11552
rect 23841 11520 26000 11522
rect 23841 11464 23846 11520
rect 23902 11464 26000 11520
rect 23841 11462 26000 11464
rect 23841 11459 23907 11462
rect 3913 11456 4229 11457
rect 3913 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4229 11456
rect 3913 11391 4229 11392
rect 9847 11456 10163 11457
rect 9847 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10163 11456
rect 9847 11391 10163 11392
rect 15781 11456 16097 11457
rect 15781 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16097 11456
rect 15781 11391 16097 11392
rect 21715 11456 22031 11457
rect 21715 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22031 11456
rect 25840 11432 26000 11462
rect 21715 11391 22031 11392
rect 17217 11386 17283 11389
rect 20846 11386 20852 11388
rect 17217 11384 20852 11386
rect 17217 11328 17222 11384
rect 17278 11328 20852 11384
rect 17217 11326 20852 11328
rect 17217 11323 17283 11326
rect 20846 11324 20852 11326
rect 20916 11324 20922 11388
rect 0 11250 160 11280
rect 3601 11250 3667 11253
rect 0 11248 3667 11250
rect 0 11192 3606 11248
rect 3662 11192 3667 11248
rect 0 11190 3667 11192
rect 0 11160 160 11190
rect 3601 11187 3667 11190
rect 5441 11250 5507 11253
rect 7005 11250 7071 11253
rect 17953 11250 18019 11253
rect 5441 11248 18019 11250
rect 5441 11192 5446 11248
rect 5502 11192 7010 11248
rect 7066 11192 17958 11248
rect 18014 11192 18019 11248
rect 5441 11190 18019 11192
rect 5441 11187 5507 11190
rect 7005 11187 7071 11190
rect 17953 11187 18019 11190
rect 2037 11114 2103 11117
rect 7414 11114 7420 11116
rect 2037 11112 7420 11114
rect 2037 11056 2042 11112
rect 2098 11056 7420 11112
rect 2037 11054 7420 11056
rect 2037 11051 2103 11054
rect 7414 11052 7420 11054
rect 7484 11052 7490 11116
rect 9029 11114 9095 11117
rect 10041 11114 10107 11117
rect 9029 11112 10107 11114
rect 9029 11056 9034 11112
rect 9090 11056 10046 11112
rect 10102 11056 10107 11112
rect 9029 11054 10107 11056
rect 9029 11051 9095 11054
rect 10041 11051 10107 11054
rect 10910 11052 10916 11116
rect 10980 11114 10986 11116
rect 11830 11114 11836 11116
rect 10980 11054 11836 11114
rect 10980 11052 10986 11054
rect 11830 11052 11836 11054
rect 11900 11052 11906 11116
rect 14917 11114 14983 11117
rect 17033 11114 17099 11117
rect 14917 11112 17099 11114
rect 14917 11056 14922 11112
rect 14978 11056 17038 11112
rect 17094 11056 17099 11112
rect 14917 11054 17099 11056
rect 14917 11051 14983 11054
rect 17033 11051 17099 11054
rect 19241 11114 19307 11117
rect 19374 11114 19380 11116
rect 19241 11112 19380 11114
rect 19241 11056 19246 11112
rect 19302 11056 19380 11112
rect 19241 11054 19380 11056
rect 19241 11051 19307 11054
rect 19374 11052 19380 11054
rect 19444 11052 19450 11116
rect 0 10978 160 11008
rect 1669 10978 1735 10981
rect 0 10976 1735 10978
rect 0 10920 1674 10976
rect 1730 10920 1735 10976
rect 0 10918 1735 10920
rect 0 10888 160 10918
rect 1669 10915 1735 10918
rect 7557 10978 7623 10981
rect 9489 10978 9555 10981
rect 7557 10976 9555 10978
rect 7557 10920 7562 10976
rect 7618 10920 9494 10976
rect 9550 10920 9555 10976
rect 7557 10918 9555 10920
rect 7557 10915 7623 10918
rect 9489 10915 9555 10918
rect 15101 10978 15167 10981
rect 16246 10978 16252 10980
rect 15101 10976 16252 10978
rect 15101 10920 15106 10976
rect 15162 10920 16252 10976
rect 15101 10918 16252 10920
rect 15101 10915 15167 10918
rect 16246 10916 16252 10918
rect 16316 10916 16322 10980
rect 25221 10978 25287 10981
rect 25840 10978 26000 11008
rect 25221 10976 26000 10978
rect 25221 10920 25226 10976
rect 25282 10920 26000 10976
rect 25221 10918 26000 10920
rect 25221 10915 25287 10918
rect 6880 10912 7196 10913
rect 6880 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7196 10912
rect 6880 10847 7196 10848
rect 12814 10912 13130 10913
rect 12814 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13130 10912
rect 12814 10847 13130 10848
rect 18748 10912 19064 10913
rect 18748 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19064 10912
rect 18748 10847 19064 10848
rect 24682 10912 24998 10913
rect 24682 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 24998 10912
rect 25840 10888 26000 10918
rect 24682 10847 24998 10848
rect 15469 10844 15535 10845
rect 15469 10842 15516 10844
rect 15424 10840 15516 10842
rect 15424 10784 15474 10840
rect 15424 10782 15516 10784
rect 15469 10780 15516 10782
rect 15580 10780 15586 10844
rect 19425 10842 19491 10845
rect 19701 10842 19767 10845
rect 19425 10840 19767 10842
rect 19425 10784 19430 10840
rect 19486 10784 19706 10840
rect 19762 10784 19767 10840
rect 19425 10782 19767 10784
rect 15469 10779 15535 10780
rect 19425 10779 19491 10782
rect 19701 10779 19767 10782
rect 0 10706 160 10736
rect 3969 10706 4035 10709
rect 0 10704 4035 10706
rect 0 10648 3974 10704
rect 4030 10648 4035 10704
rect 0 10646 4035 10648
rect 0 10616 160 10646
rect 3969 10643 4035 10646
rect 5993 10706 6059 10709
rect 11462 10706 11468 10708
rect 5993 10704 11468 10706
rect 5993 10648 5998 10704
rect 6054 10648 11468 10704
rect 5993 10646 11468 10648
rect 5993 10643 6059 10646
rect 11462 10644 11468 10646
rect 11532 10644 11538 10708
rect 11697 10706 11763 10709
rect 16481 10706 16547 10709
rect 11697 10704 16547 10706
rect 11697 10648 11702 10704
rect 11758 10648 16486 10704
rect 16542 10648 16547 10704
rect 11697 10646 16547 10648
rect 11697 10643 11763 10646
rect 16481 10643 16547 10646
rect 19333 10706 19399 10709
rect 20805 10706 20871 10709
rect 19333 10704 20871 10706
rect 19333 10648 19338 10704
rect 19394 10648 20810 10704
rect 20866 10648 20871 10704
rect 19333 10646 20871 10648
rect 19333 10643 19399 10646
rect 20805 10643 20871 10646
rect 4061 10570 4127 10573
rect 3788 10568 4127 10570
rect 3788 10512 4066 10568
rect 4122 10512 4127 10568
rect 3788 10510 4127 10512
rect 0 10434 160 10464
rect 3325 10434 3391 10437
rect 0 10432 3391 10434
rect 0 10376 3330 10432
rect 3386 10376 3391 10432
rect 0 10374 3391 10376
rect 0 10344 160 10374
rect 3325 10371 3391 10374
rect 0 10162 160 10192
rect 3049 10162 3115 10165
rect 0 10160 3115 10162
rect 0 10104 3054 10160
rect 3110 10104 3115 10160
rect 0 10102 3115 10104
rect 3788 10162 3848 10510
rect 4061 10507 4127 10510
rect 6821 10570 6887 10573
rect 12566 10570 12572 10572
rect 6821 10568 12572 10570
rect 6821 10512 6826 10568
rect 6882 10512 12572 10568
rect 6821 10510 12572 10512
rect 6821 10507 6887 10510
rect 12566 10508 12572 10510
rect 12636 10508 12642 10572
rect 23381 10434 23447 10437
rect 25840 10434 26000 10464
rect 23381 10432 26000 10434
rect 23381 10376 23386 10432
rect 23442 10376 26000 10432
rect 23381 10374 26000 10376
rect 23381 10371 23447 10374
rect 3913 10368 4229 10369
rect 3913 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4229 10368
rect 3913 10303 4229 10304
rect 9847 10368 10163 10369
rect 9847 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10163 10368
rect 9847 10303 10163 10304
rect 15781 10368 16097 10369
rect 15781 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16097 10368
rect 15781 10303 16097 10304
rect 21715 10368 22031 10369
rect 21715 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22031 10368
rect 25840 10344 26000 10374
rect 21715 10303 22031 10304
rect 3969 10162 4035 10165
rect 3788 10160 4035 10162
rect 3788 10104 3974 10160
rect 4030 10104 4035 10160
rect 3788 10102 4035 10104
rect 0 10072 160 10102
rect 3049 10099 3115 10102
rect 3969 10099 4035 10102
rect 1894 9964 1900 10028
rect 1964 10026 1970 10028
rect 2037 10026 2103 10029
rect 2681 10026 2747 10029
rect 3969 10026 4035 10029
rect 1964 10024 4035 10026
rect 1964 9968 2042 10024
rect 2098 9968 2686 10024
rect 2742 9968 3974 10024
rect 4030 9968 4035 10024
rect 1964 9966 4035 9968
rect 1964 9964 1970 9966
rect 2037 9963 2103 9966
rect 2681 9963 2747 9966
rect 3969 9963 4035 9966
rect 6310 9964 6316 10028
rect 6380 10026 6386 10028
rect 7925 10026 7991 10029
rect 6380 10024 7991 10026
rect 6380 9968 7930 10024
rect 7986 9968 7991 10024
rect 6380 9966 7991 9968
rect 6380 9964 6386 9966
rect 7925 9963 7991 9966
rect 0 9890 160 9920
rect 1761 9890 1827 9893
rect 0 9888 1827 9890
rect 0 9832 1766 9888
rect 1822 9832 1827 9888
rect 0 9830 1827 9832
rect 0 9800 160 9830
rect 1761 9827 1827 9830
rect 20294 9828 20300 9892
rect 20364 9890 20370 9892
rect 20805 9890 20871 9893
rect 20364 9888 20871 9890
rect 20364 9832 20810 9888
rect 20866 9832 20871 9888
rect 20364 9830 20871 9832
rect 20364 9828 20370 9830
rect 20805 9827 20871 9830
rect 25313 9890 25379 9893
rect 25840 9890 26000 9920
rect 25313 9888 26000 9890
rect 25313 9832 25318 9888
rect 25374 9832 26000 9888
rect 25313 9830 26000 9832
rect 25313 9827 25379 9830
rect 6880 9824 7196 9825
rect 6880 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7196 9824
rect 6880 9759 7196 9760
rect 12814 9824 13130 9825
rect 12814 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13130 9824
rect 12814 9759 13130 9760
rect 18748 9824 19064 9825
rect 18748 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19064 9824
rect 18748 9759 19064 9760
rect 24682 9824 24998 9825
rect 24682 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 24998 9824
rect 25840 9800 26000 9830
rect 24682 9759 24998 9760
rect 12249 9756 12315 9757
rect 12198 9754 12204 9756
rect 12158 9694 12204 9754
rect 12268 9752 12315 9756
rect 16205 9756 16271 9757
rect 16205 9754 16252 9756
rect 12310 9696 12315 9752
rect 12198 9692 12204 9694
rect 12268 9692 12315 9696
rect 16160 9752 16252 9754
rect 16160 9696 16210 9752
rect 16160 9694 16252 9696
rect 12249 9691 12315 9692
rect 16205 9692 16252 9694
rect 16316 9692 16322 9756
rect 16205 9691 16271 9692
rect 0 9618 160 9648
rect 1209 9618 1275 9621
rect 0 9616 1275 9618
rect 0 9560 1214 9616
rect 1270 9560 1275 9616
rect 0 9558 1275 9560
rect 0 9528 160 9558
rect 1209 9555 1275 9558
rect 2998 9556 3004 9620
rect 3068 9618 3074 9620
rect 3325 9618 3391 9621
rect 3068 9616 3391 9618
rect 3068 9560 3330 9616
rect 3386 9560 3391 9616
rect 3068 9558 3391 9560
rect 3068 9556 3074 9558
rect 3325 9555 3391 9558
rect 1577 9482 1643 9485
rect 5993 9482 6059 9485
rect 1577 9480 6059 9482
rect 1577 9424 1582 9480
rect 1638 9424 5998 9480
rect 6054 9424 6059 9480
rect 1577 9422 6059 9424
rect 1577 9419 1643 9422
rect 5993 9419 6059 9422
rect 11881 9482 11947 9485
rect 17769 9482 17835 9485
rect 11881 9480 17835 9482
rect 11881 9424 11886 9480
rect 11942 9424 17774 9480
rect 17830 9424 17835 9480
rect 11881 9422 17835 9424
rect 11881 9419 11947 9422
rect 17769 9419 17835 9422
rect 0 9346 160 9376
rect 841 9346 907 9349
rect 0 9344 907 9346
rect 0 9288 846 9344
rect 902 9288 907 9344
rect 0 9286 907 9288
rect 0 9256 160 9286
rect 841 9283 907 9286
rect 1025 9346 1091 9349
rect 2037 9346 2103 9349
rect 1025 9344 2103 9346
rect 1025 9288 1030 9344
rect 1086 9288 2042 9344
rect 2098 9288 2103 9344
rect 1025 9286 2103 9288
rect 1025 9283 1091 9286
rect 2037 9283 2103 9286
rect 24025 9346 24091 9349
rect 25840 9346 26000 9376
rect 24025 9344 26000 9346
rect 24025 9288 24030 9344
rect 24086 9288 26000 9344
rect 24025 9286 26000 9288
rect 24025 9283 24091 9286
rect 3913 9280 4229 9281
rect 3913 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4229 9280
rect 3913 9215 4229 9216
rect 9847 9280 10163 9281
rect 9847 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10163 9280
rect 9847 9215 10163 9216
rect 15781 9280 16097 9281
rect 15781 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16097 9280
rect 15781 9215 16097 9216
rect 21715 9280 22031 9281
rect 21715 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22031 9280
rect 25840 9256 26000 9286
rect 21715 9215 22031 9216
rect 24301 9210 24367 9213
rect 23246 9208 24367 9210
rect 23246 9152 24306 9208
rect 24362 9152 24367 9208
rect 23246 9150 24367 9152
rect 0 9074 160 9104
rect 1025 9074 1091 9077
rect 0 9072 1091 9074
rect 0 9016 1030 9072
rect 1086 9016 1091 9072
rect 0 9014 1091 9016
rect 0 8984 160 9014
rect 1025 9011 1091 9014
rect 11053 8938 11119 8941
rect 23246 8938 23306 9150
rect 24301 9147 24367 9150
rect 11053 8936 23306 8938
rect 11053 8880 11058 8936
rect 11114 8880 23306 8936
rect 11053 8878 23306 8880
rect 23565 8938 23631 8941
rect 23565 8936 25146 8938
rect 23565 8880 23570 8936
rect 23626 8880 25146 8936
rect 23565 8878 25146 8880
rect 11053 8875 11119 8878
rect 23565 8875 23631 8878
rect 0 8802 160 8832
rect 1577 8802 1643 8805
rect 0 8800 1643 8802
rect 0 8744 1582 8800
rect 1638 8744 1643 8800
rect 0 8742 1643 8744
rect 25086 8802 25146 8878
rect 25840 8802 26000 8832
rect 25086 8742 26000 8802
rect 0 8712 160 8742
rect 1577 8739 1643 8742
rect 6880 8736 7196 8737
rect 6880 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7196 8736
rect 6880 8671 7196 8672
rect 12814 8736 13130 8737
rect 12814 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13130 8736
rect 12814 8671 13130 8672
rect 18748 8736 19064 8737
rect 18748 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19064 8736
rect 18748 8671 19064 8672
rect 24682 8736 24998 8737
rect 24682 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 24998 8736
rect 25840 8712 26000 8742
rect 24682 8671 24998 8672
rect 0 8530 160 8560
rect 1301 8530 1367 8533
rect 0 8528 1367 8530
rect 0 8472 1306 8528
rect 1362 8472 1367 8528
rect 0 8470 1367 8472
rect 0 8440 160 8470
rect 1301 8467 1367 8470
rect 9673 8530 9739 8533
rect 18689 8530 18755 8533
rect 9673 8528 18755 8530
rect 9673 8472 9678 8528
rect 9734 8472 18694 8528
rect 18750 8472 18755 8528
rect 9673 8470 18755 8472
rect 9673 8467 9739 8470
rect 18689 8467 18755 8470
rect 2313 8394 2379 8397
rect 4889 8394 4955 8397
rect 2313 8392 4955 8394
rect 2313 8336 2318 8392
rect 2374 8336 4894 8392
rect 4950 8336 4955 8392
rect 2313 8334 4955 8336
rect 2313 8331 2379 8334
rect 4889 8331 4955 8334
rect 11789 8394 11855 8397
rect 12709 8394 12775 8397
rect 18137 8394 18203 8397
rect 11789 8392 18203 8394
rect 11789 8336 11794 8392
rect 11850 8336 12714 8392
rect 12770 8336 18142 8392
rect 18198 8336 18203 8392
rect 11789 8334 18203 8336
rect 11789 8331 11855 8334
rect 12709 8331 12775 8334
rect 18137 8331 18203 8334
rect 0 8258 160 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 160 8198
rect 1393 8195 1459 8198
rect 11789 8258 11855 8261
rect 13854 8258 13860 8260
rect 11789 8256 13860 8258
rect 11789 8200 11794 8256
rect 11850 8200 13860 8256
rect 11789 8198 13860 8200
rect 11789 8195 11855 8198
rect 13854 8196 13860 8198
rect 13924 8196 13930 8260
rect 24485 8258 24551 8261
rect 25840 8258 26000 8288
rect 24485 8256 26000 8258
rect 24485 8200 24490 8256
rect 24546 8200 26000 8256
rect 24485 8198 26000 8200
rect 24485 8195 24551 8198
rect 3913 8192 4229 8193
rect 3913 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4229 8192
rect 3913 8127 4229 8128
rect 9847 8192 10163 8193
rect 9847 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10163 8192
rect 9847 8127 10163 8128
rect 15781 8192 16097 8193
rect 15781 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16097 8192
rect 15781 8127 16097 8128
rect 21715 8192 22031 8193
rect 21715 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22031 8192
rect 25840 8168 26000 8198
rect 21715 8127 22031 8128
rect 7189 8122 7255 8125
rect 8293 8122 8359 8125
rect 7189 8120 8359 8122
rect 7189 8064 7194 8120
rect 7250 8064 8298 8120
rect 8354 8064 8359 8120
rect 7189 8062 8359 8064
rect 7189 8059 7255 8062
rect 8293 8059 8359 8062
rect 0 7986 160 8016
rect 3325 7986 3391 7989
rect 0 7984 3391 7986
rect 0 7928 3330 7984
rect 3386 7928 3391 7984
rect 0 7926 3391 7928
rect 0 7896 160 7926
rect 3325 7923 3391 7926
rect 10961 7986 11027 7989
rect 16205 7986 16271 7989
rect 10961 7984 16271 7986
rect 10961 7928 10966 7984
rect 11022 7928 16210 7984
rect 16266 7928 16271 7984
rect 10961 7926 16271 7928
rect 10961 7923 11027 7926
rect 16205 7923 16271 7926
rect 2129 7850 2195 7853
rect 8293 7850 8359 7853
rect 2129 7848 8359 7850
rect 2129 7792 2134 7848
rect 2190 7792 8298 7848
rect 8354 7792 8359 7848
rect 2129 7790 8359 7792
rect 2129 7787 2195 7790
rect 8293 7787 8359 7790
rect 0 7714 160 7744
rect 1669 7714 1735 7717
rect 0 7712 1735 7714
rect 0 7656 1674 7712
rect 1730 7656 1735 7712
rect 0 7654 1735 7656
rect 0 7624 160 7654
rect 1669 7651 1735 7654
rect 25221 7714 25287 7717
rect 25840 7714 26000 7744
rect 25221 7712 26000 7714
rect 25221 7656 25226 7712
rect 25282 7656 26000 7712
rect 25221 7654 26000 7656
rect 25221 7651 25287 7654
rect 6880 7648 7196 7649
rect 6880 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7196 7648
rect 6880 7583 7196 7584
rect 12814 7648 13130 7649
rect 12814 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13130 7648
rect 12814 7583 13130 7584
rect 18748 7648 19064 7649
rect 18748 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19064 7648
rect 18748 7583 19064 7584
rect 24682 7648 24998 7649
rect 24682 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 24998 7648
rect 25840 7624 26000 7654
rect 24682 7583 24998 7584
rect 13629 7578 13695 7581
rect 17902 7578 17908 7580
rect 13629 7576 17908 7578
rect 13629 7520 13634 7576
rect 13690 7520 17908 7576
rect 13629 7518 17908 7520
rect 13629 7515 13695 7518
rect 17902 7516 17908 7518
rect 17972 7516 17978 7580
rect 0 7442 160 7472
rect 1761 7442 1827 7445
rect 0 7440 1827 7442
rect 0 7384 1766 7440
rect 1822 7384 1827 7440
rect 0 7382 1827 7384
rect 0 7352 160 7382
rect 1761 7379 1827 7382
rect 12157 7306 12223 7309
rect 14958 7306 14964 7308
rect 12157 7304 14964 7306
rect 12157 7248 12162 7304
rect 12218 7248 14964 7304
rect 12157 7246 14964 7248
rect 12157 7243 12223 7246
rect 14958 7244 14964 7246
rect 15028 7244 15034 7308
rect 0 7170 160 7200
rect 3509 7170 3575 7173
rect 0 7168 3575 7170
rect 0 7112 3514 7168
rect 3570 7112 3575 7168
rect 0 7110 3575 7112
rect 0 7080 160 7110
rect 3509 7107 3575 7110
rect 23749 7170 23815 7173
rect 25840 7170 26000 7200
rect 23749 7168 26000 7170
rect 23749 7112 23754 7168
rect 23810 7112 26000 7168
rect 23749 7110 26000 7112
rect 23749 7107 23815 7110
rect 3913 7104 4229 7105
rect 3913 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4229 7104
rect 3913 7039 4229 7040
rect 9847 7104 10163 7105
rect 9847 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10163 7104
rect 9847 7039 10163 7040
rect 15781 7104 16097 7105
rect 15781 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16097 7104
rect 15781 7039 16097 7040
rect 21715 7104 22031 7105
rect 21715 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22031 7104
rect 25840 7080 26000 7110
rect 21715 7039 22031 7040
rect 0 6898 160 6928
rect 1209 6898 1275 6901
rect 0 6896 1275 6898
rect 0 6840 1214 6896
rect 1270 6840 1275 6896
rect 0 6838 1275 6840
rect 0 6808 160 6838
rect 1209 6835 1275 6838
rect 4245 6898 4311 6901
rect 4654 6898 4660 6900
rect 4245 6896 4660 6898
rect 4245 6840 4250 6896
rect 4306 6840 4660 6896
rect 4245 6838 4660 6840
rect 4245 6835 4311 6838
rect 4654 6836 4660 6838
rect 4724 6836 4730 6900
rect 7833 6898 7899 6901
rect 12801 6898 12867 6901
rect 20713 6898 20779 6901
rect 7833 6896 20779 6898
rect 7833 6840 7838 6896
rect 7894 6840 12806 6896
rect 12862 6840 20718 6896
rect 20774 6840 20779 6896
rect 7833 6838 20779 6840
rect 7833 6835 7899 6838
rect 12801 6835 12867 6838
rect 20713 6835 20779 6838
rect 21449 6898 21515 6901
rect 23657 6898 23723 6901
rect 21449 6896 23723 6898
rect 21449 6840 21454 6896
rect 21510 6840 23662 6896
rect 23718 6840 23723 6896
rect 21449 6838 23723 6840
rect 21449 6835 21515 6838
rect 23657 6835 23723 6838
rect 2589 6762 2655 6765
rect 9305 6762 9371 6765
rect 2589 6760 9371 6762
rect 2589 6704 2594 6760
rect 2650 6704 9310 6760
rect 9366 6704 9371 6760
rect 2589 6702 9371 6704
rect 2589 6699 2655 6702
rect 9305 6699 9371 6702
rect 17953 6762 18019 6765
rect 18137 6762 18203 6765
rect 17953 6760 18203 6762
rect 17953 6704 17958 6760
rect 18014 6704 18142 6760
rect 18198 6704 18203 6760
rect 17953 6702 18203 6704
rect 17953 6699 18019 6702
rect 18137 6699 18203 6702
rect 19425 6762 19491 6765
rect 21817 6762 21883 6765
rect 19425 6760 21883 6762
rect 19425 6704 19430 6760
rect 19486 6704 21822 6760
rect 21878 6704 21883 6760
rect 19425 6702 21883 6704
rect 19425 6699 19491 6702
rect 21817 6699 21883 6702
rect 22134 6700 22140 6764
rect 22204 6762 22210 6764
rect 23197 6762 23263 6765
rect 22204 6760 23263 6762
rect 22204 6704 23202 6760
rect 23258 6704 23263 6760
rect 22204 6702 23263 6704
rect 22204 6700 22210 6702
rect 23197 6699 23263 6702
rect 24534 6702 25146 6762
rect 0 6626 160 6656
rect 1025 6626 1091 6629
rect 24534 6626 24594 6702
rect 0 6624 1091 6626
rect 0 6568 1030 6624
rect 1086 6568 1091 6624
rect 0 6566 1091 6568
rect 0 6536 160 6566
rect 1025 6563 1091 6566
rect 20854 6566 24594 6626
rect 25086 6626 25146 6702
rect 25840 6626 26000 6656
rect 25086 6566 26000 6626
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 20854 6493 20914 6566
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 25840 6536 26000 6566
rect 24682 6495 24998 6496
rect 20854 6488 20963 6493
rect 20854 6432 20902 6488
rect 20958 6432 20963 6488
rect 20854 6430 20963 6432
rect 20897 6427 20963 6430
rect 21081 6490 21147 6493
rect 23381 6490 23447 6493
rect 21081 6488 23447 6490
rect 21081 6432 21086 6488
rect 21142 6432 23386 6488
rect 23442 6432 23447 6488
rect 21081 6430 23447 6432
rect 21081 6427 21147 6430
rect 23381 6427 23447 6430
rect 0 6354 160 6384
rect 1301 6354 1367 6357
rect 0 6352 1367 6354
rect 0 6296 1306 6352
rect 1362 6296 1367 6352
rect 0 6294 1367 6296
rect 0 6264 160 6294
rect 1301 6291 1367 6294
rect 3233 6354 3299 6357
rect 23381 6354 23447 6357
rect 3233 6352 23447 6354
rect 3233 6296 3238 6352
rect 3294 6296 23386 6352
rect 23442 6296 23447 6352
rect 3233 6294 23447 6296
rect 3233 6291 3299 6294
rect 23381 6291 23447 6294
rect 8201 6218 8267 6221
rect 17953 6218 18019 6221
rect 21357 6220 21423 6221
rect 21357 6218 21404 6220
rect 8201 6216 18019 6218
rect 8201 6160 8206 6216
rect 8262 6160 17958 6216
rect 18014 6160 18019 6216
rect 8201 6158 18019 6160
rect 21312 6216 21404 6218
rect 21312 6160 21362 6216
rect 21312 6158 21404 6160
rect 8201 6155 8267 6158
rect 17953 6155 18019 6158
rect 21357 6156 21404 6158
rect 21468 6156 21474 6220
rect 21909 6218 21975 6221
rect 22277 6218 22343 6221
rect 21909 6216 22343 6218
rect 21909 6160 21914 6216
rect 21970 6160 22282 6216
rect 22338 6160 22343 6216
rect 21909 6158 22343 6160
rect 21357 6155 21423 6156
rect 21909 6155 21975 6158
rect 22277 6155 22343 6158
rect 0 6082 160 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 160 6022
rect 1577 6019 1643 6022
rect 10542 6020 10548 6084
rect 10612 6082 10618 6084
rect 13353 6082 13419 6085
rect 10612 6080 13419 6082
rect 10612 6024 13358 6080
rect 13414 6024 13419 6080
rect 10612 6022 13419 6024
rect 10612 6020 10618 6022
rect 13353 6019 13419 6022
rect 20897 6082 20963 6085
rect 21541 6082 21607 6085
rect 20897 6080 21607 6082
rect 20897 6024 20902 6080
rect 20958 6024 21546 6080
rect 21602 6024 21607 6080
rect 20897 6022 21607 6024
rect 20897 6019 20963 6022
rect 21541 6019 21607 6022
rect 23657 6082 23723 6085
rect 25840 6082 26000 6112
rect 23657 6080 26000 6082
rect 23657 6024 23662 6080
rect 23718 6024 26000 6080
rect 23657 6022 26000 6024
rect 23657 6019 23723 6022
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 25840 5992 26000 6022
rect 21715 5951 22031 5952
rect 9305 5946 9371 5949
rect 4294 5944 9371 5946
rect 4294 5888 9310 5944
rect 9366 5888 9371 5944
rect 4294 5886 9371 5888
rect 0 5810 160 5840
rect 1301 5810 1367 5813
rect 0 5808 1367 5810
rect 0 5752 1306 5808
rect 1362 5752 1367 5808
rect 0 5750 1367 5752
rect 0 5720 160 5750
rect 1301 5747 1367 5750
rect 3550 5748 3556 5812
rect 3620 5810 3626 5812
rect 4061 5810 4127 5813
rect 4294 5810 4354 5886
rect 9305 5883 9371 5886
rect 11513 5946 11579 5949
rect 11646 5946 11652 5948
rect 11513 5944 11652 5946
rect 11513 5888 11518 5944
rect 11574 5888 11652 5944
rect 11513 5886 11652 5888
rect 11513 5883 11579 5886
rect 11646 5884 11652 5886
rect 11716 5884 11722 5948
rect 3620 5808 4354 5810
rect 3620 5752 4066 5808
rect 4122 5752 4354 5808
rect 3620 5750 4354 5752
rect 7465 5810 7531 5813
rect 12157 5810 12223 5813
rect 17493 5810 17559 5813
rect 7465 5808 12223 5810
rect 7465 5752 7470 5808
rect 7526 5752 12162 5808
rect 12218 5752 12223 5808
rect 7465 5750 12223 5752
rect 3620 5748 3626 5750
rect 4061 5747 4127 5750
rect 7465 5747 7531 5750
rect 12157 5747 12223 5750
rect 12390 5808 17559 5810
rect 12390 5752 17498 5808
rect 17554 5752 17559 5808
rect 12390 5750 17559 5752
rect 2313 5674 2379 5677
rect 6913 5674 6979 5677
rect 2313 5672 6979 5674
rect 2313 5616 2318 5672
rect 2374 5616 6918 5672
rect 6974 5616 6979 5672
rect 2313 5614 6979 5616
rect 2313 5611 2379 5614
rect 6913 5611 6979 5614
rect 7281 5674 7347 5677
rect 10041 5674 10107 5677
rect 12390 5674 12450 5750
rect 17493 5747 17559 5750
rect 22093 5810 22159 5813
rect 25681 5810 25747 5813
rect 22093 5808 25747 5810
rect 22093 5752 22098 5808
rect 22154 5752 25686 5808
rect 25742 5752 25747 5808
rect 22093 5750 25747 5752
rect 22093 5747 22159 5750
rect 25681 5747 25747 5750
rect 16389 5674 16455 5677
rect 17953 5674 18019 5677
rect 7281 5672 10107 5674
rect 7281 5616 7286 5672
rect 7342 5616 10046 5672
rect 10102 5616 10107 5672
rect 7281 5614 10107 5616
rect 7281 5611 7347 5614
rect 10041 5611 10107 5614
rect 10182 5614 12450 5674
rect 12620 5672 18019 5674
rect 12620 5616 16394 5672
rect 16450 5616 17958 5672
rect 18014 5616 18019 5672
rect 12620 5614 18019 5616
rect 0 5538 160 5568
rect 9305 5538 9371 5541
rect 10182 5538 10242 5614
rect 0 5478 1042 5538
rect 0 5448 160 5478
rect 982 5402 1042 5478
rect 9305 5536 10242 5538
rect 9305 5480 9310 5536
rect 9366 5480 10242 5536
rect 9305 5478 10242 5480
rect 11053 5538 11119 5541
rect 12620 5538 12680 5614
rect 16389 5611 16455 5614
rect 17953 5611 18019 5614
rect 22737 5540 22803 5541
rect 22686 5538 22692 5540
rect 11053 5536 12680 5538
rect 11053 5480 11058 5536
rect 11114 5480 12680 5536
rect 11053 5478 12680 5480
rect 22646 5478 22692 5538
rect 22756 5536 22803 5540
rect 22798 5480 22803 5536
rect 9305 5475 9371 5478
rect 11053 5475 11119 5478
rect 22686 5476 22692 5478
rect 22756 5476 22803 5480
rect 22870 5476 22876 5540
rect 22940 5538 22946 5540
rect 23381 5538 23447 5541
rect 22940 5536 23447 5538
rect 22940 5480 23386 5536
rect 23442 5480 23447 5536
rect 22940 5478 23447 5480
rect 22940 5476 22946 5478
rect 22737 5475 22803 5476
rect 23381 5475 23447 5478
rect 25681 5538 25747 5541
rect 25840 5538 26000 5568
rect 25681 5536 26000 5538
rect 25681 5480 25686 5536
rect 25742 5480 26000 5536
rect 25681 5478 26000 5480
rect 25681 5475 25747 5478
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 25840 5448 26000 5478
rect 24682 5407 24998 5408
rect 1761 5402 1827 5405
rect 982 5400 1827 5402
rect 982 5344 1766 5400
rect 1822 5344 1827 5400
rect 982 5342 1827 5344
rect 1761 5339 1827 5342
rect 20253 5402 20319 5405
rect 23657 5402 23723 5405
rect 20253 5400 23723 5402
rect 20253 5344 20258 5400
rect 20314 5344 23662 5400
rect 23718 5344 23723 5400
rect 20253 5342 23723 5344
rect 20253 5339 20319 5342
rect 23657 5339 23723 5342
rect 0 5266 160 5296
rect 2865 5266 2931 5269
rect 0 5264 2931 5266
rect 0 5208 2870 5264
rect 2926 5208 2931 5264
rect 0 5206 2931 5208
rect 0 5176 160 5206
rect 2865 5203 2931 5206
rect 4889 5266 4955 5269
rect 20713 5266 20779 5269
rect 4889 5264 20779 5266
rect 4889 5208 4894 5264
rect 4950 5208 20718 5264
rect 20774 5208 20779 5264
rect 4889 5206 20779 5208
rect 4889 5203 4955 5206
rect 20713 5203 20779 5206
rect 5901 5130 5967 5133
rect 12617 5130 12683 5133
rect 16205 5130 16271 5133
rect 5901 5128 12683 5130
rect 5901 5072 5906 5128
rect 5962 5072 12622 5128
rect 12678 5072 12683 5128
rect 5901 5070 12683 5072
rect 5901 5067 5967 5070
rect 12617 5067 12683 5070
rect 15564 5128 16271 5130
rect 15564 5072 16210 5128
rect 16266 5072 16271 5128
rect 15564 5070 16271 5072
rect 0 4994 160 5024
rect 15564 4997 15624 5070
rect 16205 5067 16271 5070
rect 16982 5068 16988 5132
rect 17052 5130 17058 5132
rect 19057 5130 19123 5133
rect 17052 5128 19123 5130
rect 17052 5072 19062 5128
rect 19118 5072 19123 5128
rect 17052 5070 19123 5072
rect 17052 5068 17058 5070
rect 19057 5067 19123 5070
rect 22001 5130 22067 5133
rect 22001 5128 24042 5130
rect 22001 5072 22006 5128
rect 22062 5072 24042 5128
rect 22001 5070 24042 5072
rect 22001 5067 22067 5070
rect 1393 4994 1459 4997
rect 0 4992 1459 4994
rect 0 4936 1398 4992
rect 1454 4936 1459 4992
rect 0 4934 1459 4936
rect 0 4904 160 4934
rect 1393 4931 1459 4934
rect 4521 4994 4587 4997
rect 5993 4994 6059 4997
rect 4521 4992 6059 4994
rect 4521 4936 4526 4992
rect 4582 4936 5998 4992
rect 6054 4936 6059 4992
rect 4521 4934 6059 4936
rect 4521 4931 4587 4934
rect 5993 4931 6059 4934
rect 12157 4994 12223 4997
rect 15561 4994 15627 4997
rect 12157 4992 15627 4994
rect 12157 4936 12162 4992
rect 12218 4936 15566 4992
rect 15622 4936 15627 4992
rect 12157 4934 15627 4936
rect 23982 4994 24042 5070
rect 25840 4994 26000 5024
rect 23982 4934 26000 4994
rect 12157 4931 12223 4934
rect 15561 4931 15627 4934
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 25840 4904 26000 4934
rect 21715 4863 22031 4864
rect 16573 4722 16639 4725
rect 2132 4720 16639 4722
rect 2132 4664 16578 4720
rect 16634 4664 16639 4720
rect 2132 4662 16639 4664
rect 2132 4453 2192 4662
rect 16573 4659 16639 4662
rect 17585 4722 17651 4725
rect 21541 4722 21607 4725
rect 17585 4720 21607 4722
rect 17585 4664 17590 4720
rect 17646 4664 21546 4720
rect 21602 4664 21607 4720
rect 17585 4662 21607 4664
rect 17585 4659 17651 4662
rect 21541 4659 21607 4662
rect 3969 4586 4035 4589
rect 6821 4586 6887 4589
rect 3969 4584 6887 4586
rect 3969 4528 3974 4584
rect 4030 4528 6826 4584
rect 6882 4528 6887 4584
rect 3969 4526 6887 4528
rect 3969 4523 4035 4526
rect 6821 4523 6887 4526
rect 11421 4586 11487 4589
rect 15561 4586 15627 4589
rect 11421 4584 15627 4586
rect 11421 4528 11426 4584
rect 11482 4528 15566 4584
rect 15622 4528 15627 4584
rect 11421 4526 15627 4528
rect 11421 4523 11487 4526
rect 15561 4523 15627 4526
rect 2129 4448 2195 4453
rect 2129 4392 2134 4448
rect 2190 4392 2195 4448
rect 2129 4387 2195 4392
rect 25221 4450 25287 4453
rect 25840 4450 26000 4480
rect 25221 4448 26000 4450
rect 25221 4392 25226 4448
rect 25282 4392 26000 4448
rect 25221 4390 26000 4392
rect 25221 4387 25287 4390
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 25840 4360 26000 4390
rect 24682 4319 24998 4320
rect 381 4314 447 4317
rect 4429 4314 4495 4317
rect 381 4312 4495 4314
rect 381 4256 386 4312
rect 442 4256 4434 4312
rect 4490 4256 4495 4312
rect 381 4254 4495 4256
rect 381 4251 447 4254
rect 4429 4251 4495 4254
rect 10225 4178 10291 4181
rect 13353 4178 13419 4181
rect 10225 4176 13419 4178
rect 10225 4120 10230 4176
rect 10286 4120 13358 4176
rect 13414 4120 13419 4176
rect 10225 4118 13419 4120
rect 10225 4115 10291 4118
rect 13353 4115 13419 4118
rect 17953 4178 18019 4181
rect 22645 4178 22711 4181
rect 17953 4176 22711 4178
rect 17953 4120 17958 4176
rect 18014 4120 22650 4176
rect 22706 4120 22711 4176
rect 17953 4118 22711 4120
rect 17953 4115 18019 4118
rect 22645 4115 22711 4118
rect 974 3980 980 4044
rect 1044 4042 1050 4044
rect 3325 4042 3391 4045
rect 1044 4040 3391 4042
rect 1044 3984 3330 4040
rect 3386 3984 3391 4040
rect 1044 3982 3391 3984
rect 1044 3980 1050 3982
rect 3325 3979 3391 3982
rect 10133 4042 10199 4045
rect 10685 4042 10751 4045
rect 12249 4044 12315 4045
rect 10133 4040 10751 4042
rect 10133 3984 10138 4040
rect 10194 3984 10690 4040
rect 10746 3984 10751 4040
rect 10133 3982 10751 3984
rect 10133 3979 10199 3982
rect 10685 3979 10751 3982
rect 12198 3980 12204 4044
rect 12268 4042 12315 4044
rect 13721 4042 13787 4045
rect 18321 4044 18387 4045
rect 14590 4042 14596 4044
rect 12268 4040 12360 4042
rect 12310 3984 12360 4040
rect 12268 3982 12360 3984
rect 13721 4040 14596 4042
rect 13721 3984 13726 4040
rect 13782 3984 14596 4040
rect 13721 3982 14596 3984
rect 12268 3980 12315 3982
rect 12249 3979 12315 3980
rect 13721 3979 13787 3982
rect 14590 3980 14596 3982
rect 14660 3980 14666 4044
rect 18270 4042 18276 4044
rect 18230 3982 18276 4042
rect 18340 4040 18387 4044
rect 18382 3984 18387 4040
rect 18270 3980 18276 3982
rect 18340 3980 18387 3984
rect 18321 3979 18387 3980
rect 19517 4042 19583 4045
rect 20897 4042 20963 4045
rect 19517 4040 20963 4042
rect 19517 3984 19522 4040
rect 19578 3984 20902 4040
rect 20958 3984 20963 4040
rect 19517 3982 20963 3984
rect 19517 3979 19583 3982
rect 20897 3979 20963 3982
rect 21449 4042 21515 4045
rect 21449 4040 24042 4042
rect 21449 3984 21454 4040
rect 21510 3984 24042 4040
rect 21449 3982 24042 3984
rect 21449 3979 21515 3982
rect 18229 3906 18295 3909
rect 20529 3906 20595 3909
rect 18229 3904 20595 3906
rect 18229 3848 18234 3904
rect 18290 3848 20534 3904
rect 20590 3848 20595 3904
rect 18229 3846 20595 3848
rect 23982 3906 24042 3982
rect 25840 3906 26000 3936
rect 23982 3846 26000 3906
rect 18229 3843 18295 3846
rect 20529 3843 20595 3846
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 25840 3816 26000 3846
rect 21715 3775 22031 3776
rect 5073 3770 5139 3773
rect 9489 3770 9555 3773
rect 5073 3768 9555 3770
rect 5073 3712 5078 3768
rect 5134 3712 9494 3768
rect 9550 3712 9555 3768
rect 5073 3710 9555 3712
rect 5073 3707 5139 3710
rect 9489 3707 9555 3710
rect 10501 3770 10567 3773
rect 10501 3768 12450 3770
rect 10501 3712 10506 3768
rect 10562 3712 12450 3768
rect 10501 3710 12450 3712
rect 10501 3707 10567 3710
rect 6545 3634 6611 3637
rect 12065 3634 12131 3637
rect 6545 3632 12131 3634
rect 6545 3576 6550 3632
rect 6606 3576 12070 3632
rect 12126 3576 12131 3632
rect 6545 3574 12131 3576
rect 12390 3634 12450 3710
rect 17534 3708 17540 3772
rect 17604 3770 17610 3772
rect 18689 3770 18755 3773
rect 17604 3768 18755 3770
rect 17604 3712 18694 3768
rect 18750 3712 18755 3768
rect 17604 3710 18755 3712
rect 17604 3708 17610 3710
rect 18689 3707 18755 3710
rect 19149 3772 19215 3773
rect 19149 3768 19196 3772
rect 19260 3770 19266 3772
rect 19149 3712 19154 3768
rect 19149 3708 19196 3712
rect 19260 3710 19306 3770
rect 19260 3708 19266 3710
rect 19149 3707 19215 3708
rect 20805 3634 20871 3637
rect 12390 3632 20871 3634
rect 12390 3576 20810 3632
rect 20866 3576 20871 3632
rect 12390 3574 20871 3576
rect 6545 3571 6611 3574
rect 12065 3571 12131 3574
rect 20805 3571 20871 3574
rect 2681 3498 2747 3501
rect 9765 3498 9831 3501
rect 10501 3498 10567 3501
rect 2681 3496 9831 3498
rect 2681 3440 2686 3496
rect 2742 3440 9770 3496
rect 9826 3440 9831 3496
rect 2681 3438 9831 3440
rect 2681 3435 2747 3438
rect 9765 3435 9831 3438
rect 9998 3496 10567 3498
rect 9998 3440 10506 3496
rect 10562 3440 10567 3496
rect 9998 3438 10567 3440
rect 790 3300 796 3364
rect 860 3362 866 3364
rect 4889 3362 4955 3365
rect 860 3360 4955 3362
rect 860 3304 4894 3360
rect 4950 3304 4955 3360
rect 860 3302 4955 3304
rect 860 3300 866 3302
rect 4889 3299 4955 3302
rect 9121 3362 9187 3365
rect 9998 3362 10058 3438
rect 10501 3435 10567 3438
rect 18229 3498 18295 3501
rect 21265 3498 21331 3501
rect 18229 3496 20178 3498
rect 18229 3440 18234 3496
rect 18290 3440 20178 3496
rect 18229 3438 20178 3440
rect 18229 3435 18295 3438
rect 9121 3360 10058 3362
rect 9121 3304 9126 3360
rect 9182 3304 10058 3360
rect 9121 3302 10058 3304
rect 10133 3362 10199 3365
rect 12617 3364 12683 3365
rect 10910 3362 10916 3364
rect 10133 3360 10916 3362
rect 10133 3304 10138 3360
rect 10194 3304 10916 3360
rect 10133 3302 10916 3304
rect 9121 3299 9187 3302
rect 10133 3299 10199 3302
rect 10910 3300 10916 3302
rect 10980 3300 10986 3364
rect 12566 3362 12572 3364
rect 12526 3302 12572 3362
rect 12636 3360 12683 3364
rect 12678 3304 12683 3360
rect 12566 3300 12572 3302
rect 12636 3300 12683 3304
rect 12617 3299 12683 3300
rect 18137 3362 18203 3365
rect 18597 3362 18663 3365
rect 18137 3360 18663 3362
rect 18137 3304 18142 3360
rect 18198 3304 18602 3360
rect 18658 3304 18663 3360
rect 18137 3302 18663 3304
rect 20118 3362 20178 3438
rect 21265 3496 25146 3498
rect 21265 3440 21270 3496
rect 21326 3440 25146 3496
rect 21265 3438 25146 3440
rect 21265 3435 21331 3438
rect 25086 3362 25146 3438
rect 25840 3362 26000 3392
rect 20118 3302 24042 3362
rect 25086 3302 26000 3362
rect 18137 3299 18203 3302
rect 18597 3299 18663 3302
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 9949 3226 10015 3229
rect 10869 3226 10935 3229
rect 12157 3226 12223 3229
rect 9949 3224 12223 3226
rect 9949 3168 9954 3224
rect 10010 3168 10874 3224
rect 10930 3168 12162 3224
rect 12218 3168 12223 3224
rect 9949 3166 12223 3168
rect 9949 3163 10015 3166
rect 10869 3163 10935 3166
rect 12157 3163 12223 3166
rect 19149 3226 19215 3229
rect 22134 3226 22140 3228
rect 19149 3224 22140 3226
rect 19149 3168 19154 3224
rect 19210 3168 22140 3224
rect 19149 3166 22140 3168
rect 19149 3163 19215 3166
rect 22134 3164 22140 3166
rect 22204 3164 22210 3228
rect 1853 3090 1919 3093
rect 22645 3090 22711 3093
rect 1853 3088 22711 3090
rect 1853 3032 1858 3088
rect 1914 3032 22650 3088
rect 22706 3032 22711 3088
rect 1853 3030 22711 3032
rect 23982 3090 24042 3302
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 25840 3272 26000 3302
rect 24682 3231 24998 3232
rect 25681 3226 25747 3229
rect 25086 3224 25747 3226
rect 25086 3168 25686 3224
rect 25742 3168 25747 3224
rect 25086 3166 25747 3168
rect 25086 3090 25146 3166
rect 25681 3163 25747 3166
rect 23982 3030 25146 3090
rect 1853 3027 1919 3030
rect 22645 3027 22711 3030
rect 4061 2954 4127 2957
rect 11053 2954 11119 2957
rect 4061 2952 11119 2954
rect 4061 2896 4066 2952
rect 4122 2896 11058 2952
rect 11114 2896 11119 2952
rect 4061 2894 11119 2896
rect 4061 2891 4127 2894
rect 11053 2891 11119 2894
rect 17953 2954 18019 2957
rect 18689 2954 18755 2957
rect 17953 2952 18755 2954
rect 17953 2896 17958 2952
rect 18014 2896 18694 2952
rect 18750 2896 18755 2952
rect 17953 2894 18755 2896
rect 17953 2891 18019 2894
rect 18689 2891 18755 2894
rect 20713 2954 20779 2957
rect 20713 2952 22708 2954
rect 20713 2896 20718 2952
rect 20774 2896 22708 2952
rect 20713 2894 22708 2896
rect 20713 2891 20779 2894
rect 17033 2818 17099 2821
rect 20713 2818 20779 2821
rect 17033 2816 20779 2818
rect 17033 2760 17038 2816
rect 17094 2760 20718 2816
rect 20774 2760 20779 2816
rect 17033 2758 20779 2760
rect 22648 2818 22708 2894
rect 25840 2818 26000 2848
rect 22648 2758 26000 2818
rect 17033 2755 17099 2758
rect 20713 2755 20779 2758
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 25840 2728 26000 2758
rect 21715 2687 22031 2688
rect 2129 2684 2195 2685
rect 9489 2684 9555 2685
rect 2078 2620 2084 2684
rect 2148 2682 2195 2684
rect 2148 2680 2240 2682
rect 2190 2624 2240 2680
rect 2148 2622 2240 2624
rect 2148 2620 2195 2622
rect 9438 2620 9444 2684
rect 9508 2682 9555 2684
rect 12893 2682 12959 2685
rect 13302 2682 13308 2684
rect 9508 2680 9600 2682
rect 9550 2624 9600 2680
rect 9508 2622 9600 2624
rect 12893 2680 13308 2682
rect 12893 2624 12898 2680
rect 12954 2624 13308 2680
rect 12893 2622 13308 2624
rect 9508 2620 9555 2622
rect 2129 2619 2195 2620
rect 9489 2619 9555 2620
rect 12893 2619 12959 2622
rect 13302 2620 13308 2622
rect 13372 2620 13378 2684
rect 17217 2682 17283 2685
rect 17350 2682 17356 2684
rect 17217 2680 17356 2682
rect 17217 2624 17222 2680
rect 17278 2624 17356 2680
rect 17217 2622 17356 2624
rect 17217 2619 17283 2622
rect 17350 2620 17356 2622
rect 17420 2620 17426 2684
rect 17493 2682 17559 2685
rect 17953 2682 18019 2685
rect 18505 2684 18571 2685
rect 18454 2682 18460 2684
rect 17493 2680 18019 2682
rect 17493 2624 17498 2680
rect 17554 2624 17958 2680
rect 18014 2624 18019 2680
rect 17493 2622 18019 2624
rect 18414 2622 18460 2682
rect 18524 2680 18571 2684
rect 18566 2624 18571 2680
rect 17493 2619 17559 2622
rect 17953 2619 18019 2622
rect 18454 2620 18460 2622
rect 18524 2620 18571 2624
rect 18505 2619 18571 2620
rect 18689 2682 18755 2685
rect 19190 2682 19196 2684
rect 18689 2680 19196 2682
rect 18689 2624 18694 2680
rect 18750 2624 19196 2680
rect 18689 2622 19196 2624
rect 18689 2619 18755 2622
rect 19190 2620 19196 2622
rect 19260 2620 19266 2684
rect 19425 2682 19491 2685
rect 19558 2682 19564 2684
rect 19425 2680 19564 2682
rect 19425 2624 19430 2680
rect 19486 2624 19564 2680
rect 19425 2622 19564 2624
rect 19425 2619 19491 2622
rect 19558 2620 19564 2622
rect 19628 2620 19634 2684
rect 19793 2682 19859 2685
rect 19926 2682 19932 2684
rect 19793 2680 19932 2682
rect 19793 2624 19798 2680
rect 19854 2624 19932 2680
rect 19793 2622 19932 2624
rect 19793 2619 19859 2622
rect 19926 2620 19932 2622
rect 19996 2620 20002 2684
rect 2630 2484 2636 2548
rect 2700 2546 2706 2548
rect 6545 2546 6611 2549
rect 15561 2546 15627 2549
rect 2700 2544 6611 2546
rect 2700 2488 6550 2544
rect 6606 2488 6611 2544
rect 2700 2486 6611 2488
rect 2700 2484 2706 2486
rect 6545 2483 6611 2486
rect 6686 2486 12450 2546
rect 1158 2348 1164 2412
rect 1228 2410 1234 2412
rect 6177 2410 6243 2413
rect 1228 2408 6243 2410
rect 1228 2352 6182 2408
rect 6238 2352 6243 2408
rect 1228 2350 6243 2352
rect 1228 2348 1234 2350
rect 6177 2347 6243 2350
rect 1117 2274 1183 2277
rect 6686 2274 6746 2486
rect 7189 2410 7255 2413
rect 8477 2410 8543 2413
rect 7189 2408 8543 2410
rect 7189 2352 7194 2408
rect 7250 2352 8482 2408
rect 8538 2352 8543 2408
rect 7189 2350 8543 2352
rect 7189 2347 7255 2350
rect 8477 2347 8543 2350
rect 9213 2410 9279 2413
rect 10542 2410 10548 2412
rect 9213 2408 10548 2410
rect 9213 2352 9218 2408
rect 9274 2352 10548 2408
rect 9213 2350 10548 2352
rect 9213 2347 9279 2350
rect 10542 2348 10548 2350
rect 10612 2348 10618 2412
rect 11789 2410 11855 2413
rect 12014 2410 12020 2412
rect 11789 2408 12020 2410
rect 11789 2352 11794 2408
rect 11850 2352 12020 2408
rect 11789 2350 12020 2352
rect 11789 2347 11855 2350
rect 12014 2348 12020 2350
rect 12084 2348 12090 2412
rect 12390 2410 12450 2486
rect 15561 2544 21098 2546
rect 15561 2488 15566 2544
rect 15622 2488 21098 2544
rect 15561 2486 21098 2488
rect 15561 2483 15627 2486
rect 13261 2410 13327 2413
rect 12390 2408 13327 2410
rect 12390 2352 13266 2408
rect 13322 2352 13327 2408
rect 12390 2350 13327 2352
rect 13261 2347 13327 2350
rect 16389 2410 16455 2413
rect 17718 2410 17724 2412
rect 16389 2408 17724 2410
rect 16389 2352 16394 2408
rect 16450 2352 17724 2408
rect 16389 2350 17724 2352
rect 16389 2347 16455 2350
rect 17718 2348 17724 2350
rect 17788 2348 17794 2412
rect 18137 2410 18203 2413
rect 18597 2410 18663 2413
rect 18137 2408 18663 2410
rect 18137 2352 18142 2408
rect 18198 2352 18602 2408
rect 18658 2352 18663 2408
rect 18137 2350 18663 2352
rect 21038 2410 21098 2486
rect 25589 2410 25655 2413
rect 21038 2408 25655 2410
rect 21038 2352 25594 2408
rect 25650 2352 25655 2408
rect 21038 2350 25655 2352
rect 18137 2347 18203 2350
rect 18597 2347 18663 2350
rect 25589 2347 25655 2350
rect 7741 2276 7807 2277
rect 8109 2276 8175 2277
rect 7741 2274 7788 2276
rect 1117 2272 6746 2274
rect 1117 2216 1122 2272
rect 1178 2216 6746 2272
rect 1117 2214 6746 2216
rect 7696 2272 7788 2274
rect 7696 2216 7746 2272
rect 7696 2214 7788 2216
rect 1117 2211 1183 2214
rect 7741 2212 7788 2214
rect 7852 2212 7858 2276
rect 8109 2274 8156 2276
rect 8064 2272 8156 2274
rect 8064 2216 8114 2272
rect 8064 2214 8156 2216
rect 8109 2212 8156 2214
rect 8220 2212 8226 2276
rect 8385 2274 8451 2277
rect 8845 2276 8911 2277
rect 8518 2274 8524 2276
rect 8385 2272 8524 2274
rect 8385 2216 8390 2272
rect 8446 2216 8524 2272
rect 8385 2214 8524 2216
rect 7741 2211 7807 2212
rect 8109 2211 8175 2212
rect 8385 2211 8451 2214
rect 8518 2212 8524 2214
rect 8588 2212 8594 2276
rect 8845 2274 8892 2276
rect 8800 2272 8892 2274
rect 8800 2216 8850 2272
rect 8800 2214 8892 2216
rect 8845 2212 8892 2214
rect 8956 2212 8962 2276
rect 25681 2274 25747 2277
rect 25840 2274 26000 2304
rect 25681 2272 26000 2274
rect 25681 2216 25686 2272
rect 25742 2216 26000 2272
rect 25681 2214 26000 2216
rect 8845 2211 8911 2212
rect 25681 2211 25747 2214
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 25840 2184 26000 2214
rect 24682 2143 24998 2144
rect 7649 2138 7715 2141
rect 12617 2138 12683 2141
rect 7649 2136 12683 2138
rect 7649 2080 7654 2136
rect 7710 2080 12622 2136
rect 12678 2080 12683 2136
rect 7649 2078 12683 2080
rect 7649 2075 7715 2078
rect 12617 2075 12683 2078
rect 933 2002 999 2005
rect 12065 2002 12131 2005
rect 933 2000 12131 2002
rect 933 1944 938 2000
rect 994 1944 12070 2000
rect 12126 1944 12131 2000
rect 933 1942 12131 1944
rect 933 1939 999 1942
rect 12065 1939 12131 1942
rect 13537 2002 13603 2005
rect 20662 2002 20668 2004
rect 13537 2000 20668 2002
rect 13537 1944 13542 2000
rect 13598 1944 20668 2000
rect 13537 1942 20668 1944
rect 13537 1939 13603 1942
rect 20662 1940 20668 1942
rect 20732 1940 20738 2004
rect 5533 1866 5599 1869
rect 9673 1866 9739 1869
rect 5533 1864 9739 1866
rect 5533 1808 5538 1864
rect 5594 1808 9678 1864
rect 9734 1808 9739 1864
rect 5533 1806 9739 1808
rect 5533 1803 5599 1806
rect 9673 1803 9739 1806
rect 25840 1730 26000 1760
rect 23982 1670 26000 1730
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 21357 1458 21423 1461
rect 23982 1458 24042 1670
rect 25840 1640 26000 1670
rect 21357 1456 24042 1458
rect 21357 1400 21362 1456
rect 21418 1400 24042 1456
rect 21357 1398 24042 1400
rect 21357 1395 21423 1398
rect 3969 1322 4035 1325
rect 5533 1324 5599 1325
rect 6545 1324 6611 1325
rect 4838 1322 4844 1324
rect 3969 1320 4844 1322
rect 3969 1264 3974 1320
rect 4030 1264 4844 1320
rect 3969 1262 4844 1264
rect 3969 1259 4035 1262
rect 4838 1260 4844 1262
rect 4908 1260 4914 1324
rect 5533 1320 5580 1324
rect 5644 1322 5650 1324
rect 5533 1264 5538 1320
rect 5533 1260 5580 1264
rect 5644 1262 5690 1322
rect 5644 1260 5650 1262
rect 6494 1260 6500 1324
rect 6564 1322 6611 1324
rect 7925 1324 7991 1325
rect 8661 1324 8727 1325
rect 16481 1324 16547 1325
rect 7925 1322 7972 1324
rect 6564 1320 6656 1322
rect 6606 1264 6656 1320
rect 6564 1262 6656 1264
rect 7880 1320 7972 1322
rect 7880 1264 7930 1320
rect 7880 1262 7972 1264
rect 6564 1260 6611 1262
rect 5533 1259 5599 1260
rect 6545 1259 6611 1260
rect 7925 1260 7972 1262
rect 8036 1260 8042 1324
rect 8661 1322 8708 1324
rect 8616 1320 8708 1322
rect 8616 1264 8666 1320
rect 8616 1262 8708 1264
rect 8661 1260 8708 1262
rect 8772 1260 8778 1324
rect 16430 1322 16436 1324
rect 16390 1262 16436 1322
rect 16500 1320 16547 1324
rect 16542 1264 16547 1320
rect 16430 1260 16436 1262
rect 16500 1260 16547 1264
rect 7925 1259 7991 1260
rect 8661 1259 8727 1260
rect 16481 1259 16547 1260
rect 21081 1322 21147 1325
rect 21081 1320 25146 1322
rect 21081 1264 21086 1320
rect 21142 1264 25146 1320
rect 21081 1262 25146 1264
rect 21081 1259 21147 1262
rect 606 1124 612 1188
rect 676 1186 682 1188
rect 4061 1186 4127 1189
rect 676 1184 4127 1186
rect 676 1128 4066 1184
rect 4122 1128 4127 1184
rect 676 1126 4127 1128
rect 676 1124 682 1126
rect 4061 1123 4127 1126
rect 6126 1124 6132 1188
rect 6196 1186 6202 1188
rect 6729 1186 6795 1189
rect 6196 1184 6795 1186
rect 6196 1128 6734 1184
rect 6790 1128 6795 1184
rect 6196 1126 6795 1128
rect 25086 1186 25146 1262
rect 25840 1186 26000 1216
rect 25086 1126 26000 1186
rect 6196 1124 6202 1126
rect 6729 1123 6795 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 25840 1096 26000 1126
rect 24682 1055 24998 1056
rect 20437 642 20503 645
rect 25840 642 26000 672
rect 20437 640 26000 642
rect 20437 584 20442 640
rect 20498 584 26000 640
rect 20437 582 26000 584
rect 20437 579 20503 582
rect 25840 552 26000 582
<< via3 >>
rect 6886 43548 6950 43552
rect 6886 43492 6890 43548
rect 6890 43492 6946 43548
rect 6946 43492 6950 43548
rect 6886 43488 6950 43492
rect 6966 43548 7030 43552
rect 6966 43492 6970 43548
rect 6970 43492 7026 43548
rect 7026 43492 7030 43548
rect 6966 43488 7030 43492
rect 7046 43548 7110 43552
rect 7046 43492 7050 43548
rect 7050 43492 7106 43548
rect 7106 43492 7110 43548
rect 7046 43488 7110 43492
rect 7126 43548 7190 43552
rect 7126 43492 7130 43548
rect 7130 43492 7186 43548
rect 7186 43492 7190 43548
rect 7126 43488 7190 43492
rect 12820 43548 12884 43552
rect 12820 43492 12824 43548
rect 12824 43492 12880 43548
rect 12880 43492 12884 43548
rect 12820 43488 12884 43492
rect 12900 43548 12964 43552
rect 12900 43492 12904 43548
rect 12904 43492 12960 43548
rect 12960 43492 12964 43548
rect 12900 43488 12964 43492
rect 12980 43548 13044 43552
rect 12980 43492 12984 43548
rect 12984 43492 13040 43548
rect 13040 43492 13044 43548
rect 12980 43488 13044 43492
rect 13060 43548 13124 43552
rect 13060 43492 13064 43548
rect 13064 43492 13120 43548
rect 13120 43492 13124 43548
rect 13060 43488 13124 43492
rect 18754 43548 18818 43552
rect 18754 43492 18758 43548
rect 18758 43492 18814 43548
rect 18814 43492 18818 43548
rect 18754 43488 18818 43492
rect 18834 43548 18898 43552
rect 18834 43492 18838 43548
rect 18838 43492 18894 43548
rect 18894 43492 18898 43548
rect 18834 43488 18898 43492
rect 18914 43548 18978 43552
rect 18914 43492 18918 43548
rect 18918 43492 18974 43548
rect 18974 43492 18978 43548
rect 18914 43488 18978 43492
rect 18994 43548 19058 43552
rect 18994 43492 18998 43548
rect 18998 43492 19054 43548
rect 19054 43492 19058 43548
rect 18994 43488 19058 43492
rect 24688 43548 24752 43552
rect 24688 43492 24692 43548
rect 24692 43492 24748 43548
rect 24748 43492 24752 43548
rect 24688 43488 24752 43492
rect 24768 43548 24832 43552
rect 24768 43492 24772 43548
rect 24772 43492 24828 43548
rect 24828 43492 24832 43548
rect 24768 43488 24832 43492
rect 24848 43548 24912 43552
rect 24848 43492 24852 43548
rect 24852 43492 24908 43548
rect 24908 43492 24912 43548
rect 24848 43488 24912 43492
rect 24928 43548 24992 43552
rect 24928 43492 24932 43548
rect 24932 43492 24988 43548
rect 24988 43492 24992 43548
rect 24928 43488 24992 43492
rect 3919 43004 3983 43008
rect 3919 42948 3923 43004
rect 3923 42948 3979 43004
rect 3979 42948 3983 43004
rect 3919 42944 3983 42948
rect 3999 43004 4063 43008
rect 3999 42948 4003 43004
rect 4003 42948 4059 43004
rect 4059 42948 4063 43004
rect 3999 42944 4063 42948
rect 4079 43004 4143 43008
rect 4079 42948 4083 43004
rect 4083 42948 4139 43004
rect 4139 42948 4143 43004
rect 4079 42944 4143 42948
rect 4159 43004 4223 43008
rect 4159 42948 4163 43004
rect 4163 42948 4219 43004
rect 4219 42948 4223 43004
rect 4159 42944 4223 42948
rect 9853 43004 9917 43008
rect 9853 42948 9857 43004
rect 9857 42948 9913 43004
rect 9913 42948 9917 43004
rect 9853 42944 9917 42948
rect 9933 43004 9997 43008
rect 9933 42948 9937 43004
rect 9937 42948 9993 43004
rect 9993 42948 9997 43004
rect 9933 42944 9997 42948
rect 10013 43004 10077 43008
rect 10013 42948 10017 43004
rect 10017 42948 10073 43004
rect 10073 42948 10077 43004
rect 10013 42944 10077 42948
rect 10093 43004 10157 43008
rect 10093 42948 10097 43004
rect 10097 42948 10153 43004
rect 10153 42948 10157 43004
rect 10093 42944 10157 42948
rect 15787 43004 15851 43008
rect 15787 42948 15791 43004
rect 15791 42948 15847 43004
rect 15847 42948 15851 43004
rect 15787 42944 15851 42948
rect 15867 43004 15931 43008
rect 15867 42948 15871 43004
rect 15871 42948 15927 43004
rect 15927 42948 15931 43004
rect 15867 42944 15931 42948
rect 15947 43004 16011 43008
rect 15947 42948 15951 43004
rect 15951 42948 16007 43004
rect 16007 42948 16011 43004
rect 15947 42944 16011 42948
rect 16027 43004 16091 43008
rect 16027 42948 16031 43004
rect 16031 42948 16087 43004
rect 16087 42948 16091 43004
rect 16027 42944 16091 42948
rect 21721 43004 21785 43008
rect 21721 42948 21725 43004
rect 21725 42948 21781 43004
rect 21781 42948 21785 43004
rect 21721 42944 21785 42948
rect 21801 43004 21865 43008
rect 21801 42948 21805 43004
rect 21805 42948 21861 43004
rect 21861 42948 21865 43004
rect 21801 42944 21865 42948
rect 21881 43004 21945 43008
rect 21881 42948 21885 43004
rect 21885 42948 21941 43004
rect 21941 42948 21945 43004
rect 21881 42944 21945 42948
rect 21961 43004 22025 43008
rect 21961 42948 21965 43004
rect 21965 42948 22021 43004
rect 22021 42948 22025 43004
rect 21961 42944 22025 42948
rect 11836 42876 11900 42940
rect 12204 42936 12268 42940
rect 12204 42880 12254 42936
rect 12254 42880 12268 42936
rect 12204 42876 12268 42880
rect 12572 42936 12636 42940
rect 12572 42880 12586 42936
rect 12586 42880 12636 42936
rect 12572 42876 12636 42880
rect 13860 42936 13924 42940
rect 13860 42880 13874 42936
rect 13874 42880 13924 42936
rect 13860 42876 13924 42880
rect 14412 42876 14476 42940
rect 14964 42936 15028 42940
rect 14964 42880 14978 42936
rect 14978 42880 15028 42936
rect 14964 42876 15028 42880
rect 15516 42876 15580 42940
rect 6886 42460 6950 42464
rect 6886 42404 6890 42460
rect 6890 42404 6946 42460
rect 6946 42404 6950 42460
rect 6886 42400 6950 42404
rect 6966 42460 7030 42464
rect 6966 42404 6970 42460
rect 6970 42404 7026 42460
rect 7026 42404 7030 42460
rect 6966 42400 7030 42404
rect 7046 42460 7110 42464
rect 7046 42404 7050 42460
rect 7050 42404 7106 42460
rect 7106 42404 7110 42460
rect 7046 42400 7110 42404
rect 7126 42460 7190 42464
rect 7126 42404 7130 42460
rect 7130 42404 7186 42460
rect 7186 42404 7190 42460
rect 7126 42400 7190 42404
rect 12820 42460 12884 42464
rect 12820 42404 12824 42460
rect 12824 42404 12880 42460
rect 12880 42404 12884 42460
rect 12820 42400 12884 42404
rect 12900 42460 12964 42464
rect 12900 42404 12904 42460
rect 12904 42404 12960 42460
rect 12960 42404 12964 42460
rect 12900 42400 12964 42404
rect 12980 42460 13044 42464
rect 12980 42404 12984 42460
rect 12984 42404 13040 42460
rect 13040 42404 13044 42460
rect 12980 42400 13044 42404
rect 13060 42460 13124 42464
rect 13060 42404 13064 42460
rect 13064 42404 13120 42460
rect 13120 42404 13124 42460
rect 13060 42400 13124 42404
rect 18754 42460 18818 42464
rect 18754 42404 18758 42460
rect 18758 42404 18814 42460
rect 18814 42404 18818 42460
rect 18754 42400 18818 42404
rect 18834 42460 18898 42464
rect 18834 42404 18838 42460
rect 18838 42404 18894 42460
rect 18894 42404 18898 42460
rect 18834 42400 18898 42404
rect 18914 42460 18978 42464
rect 18914 42404 18918 42460
rect 18918 42404 18974 42460
rect 18974 42404 18978 42460
rect 18914 42400 18978 42404
rect 18994 42460 19058 42464
rect 18994 42404 18998 42460
rect 18998 42404 19054 42460
rect 19054 42404 19058 42460
rect 18994 42400 19058 42404
rect 24688 42460 24752 42464
rect 24688 42404 24692 42460
rect 24692 42404 24748 42460
rect 24748 42404 24752 42460
rect 24688 42400 24752 42404
rect 24768 42460 24832 42464
rect 24768 42404 24772 42460
rect 24772 42404 24828 42460
rect 24828 42404 24832 42460
rect 24768 42400 24832 42404
rect 24848 42460 24912 42464
rect 24848 42404 24852 42460
rect 24852 42404 24908 42460
rect 24908 42404 24912 42460
rect 24848 42400 24912 42404
rect 24928 42460 24992 42464
rect 24928 42404 24932 42460
rect 24932 42404 24988 42460
rect 24988 42404 24992 42460
rect 24928 42400 24992 42404
rect 7604 42196 7668 42260
rect 7788 42060 7852 42124
rect 8708 42060 8772 42124
rect 3919 41916 3983 41920
rect 3919 41860 3923 41916
rect 3923 41860 3979 41916
rect 3979 41860 3983 41916
rect 3919 41856 3983 41860
rect 3999 41916 4063 41920
rect 3999 41860 4003 41916
rect 4003 41860 4059 41916
rect 4059 41860 4063 41916
rect 3999 41856 4063 41860
rect 4079 41916 4143 41920
rect 4079 41860 4083 41916
rect 4083 41860 4139 41916
rect 4139 41860 4143 41916
rect 4079 41856 4143 41860
rect 4159 41916 4223 41920
rect 4159 41860 4163 41916
rect 4163 41860 4219 41916
rect 4219 41860 4223 41916
rect 4159 41856 4223 41860
rect 9853 41916 9917 41920
rect 9853 41860 9857 41916
rect 9857 41860 9913 41916
rect 9913 41860 9917 41916
rect 9853 41856 9917 41860
rect 9933 41916 9997 41920
rect 9933 41860 9937 41916
rect 9937 41860 9993 41916
rect 9993 41860 9997 41916
rect 9933 41856 9997 41860
rect 10013 41916 10077 41920
rect 10013 41860 10017 41916
rect 10017 41860 10073 41916
rect 10073 41860 10077 41916
rect 10013 41856 10077 41860
rect 10093 41916 10157 41920
rect 10093 41860 10097 41916
rect 10097 41860 10153 41916
rect 10153 41860 10157 41916
rect 10093 41856 10157 41860
rect 15787 41916 15851 41920
rect 15787 41860 15791 41916
rect 15791 41860 15847 41916
rect 15847 41860 15851 41916
rect 15787 41856 15851 41860
rect 15867 41916 15931 41920
rect 15867 41860 15871 41916
rect 15871 41860 15927 41916
rect 15927 41860 15931 41916
rect 15867 41856 15931 41860
rect 15947 41916 16011 41920
rect 15947 41860 15951 41916
rect 15951 41860 16007 41916
rect 16007 41860 16011 41916
rect 15947 41856 16011 41860
rect 16027 41916 16091 41920
rect 16027 41860 16031 41916
rect 16031 41860 16087 41916
rect 16087 41860 16091 41916
rect 16027 41856 16091 41860
rect 21721 41916 21785 41920
rect 21721 41860 21725 41916
rect 21725 41860 21781 41916
rect 21781 41860 21785 41916
rect 21721 41856 21785 41860
rect 21801 41916 21865 41920
rect 21801 41860 21805 41916
rect 21805 41860 21861 41916
rect 21861 41860 21865 41916
rect 21801 41856 21865 41860
rect 21881 41916 21945 41920
rect 21881 41860 21885 41916
rect 21885 41860 21941 41916
rect 21941 41860 21945 41916
rect 21881 41856 21945 41860
rect 21961 41916 22025 41920
rect 21961 41860 21965 41916
rect 21965 41860 22021 41916
rect 22021 41860 22025 41916
rect 21961 41856 22025 41860
rect 6316 41788 6380 41852
rect 8156 41788 8220 41852
rect 9444 41848 9508 41852
rect 9444 41792 9458 41848
rect 9458 41792 9508 41848
rect 9444 41788 9508 41792
rect 17540 41788 17604 41852
rect 1164 41652 1228 41716
rect 8524 41652 8588 41716
rect 16436 41712 16500 41716
rect 16436 41656 16450 41712
rect 16450 41656 16500 41712
rect 16436 41652 16500 41656
rect 17356 41652 17420 41716
rect 18460 41712 18524 41716
rect 18460 41656 18474 41712
rect 18474 41656 18524 41712
rect 18460 41652 18524 41656
rect 19380 41712 19444 41716
rect 19380 41656 19430 41712
rect 19430 41656 19444 41712
rect 19380 41652 19444 41656
rect 796 41516 860 41580
rect 4660 41576 4724 41580
rect 4660 41520 4674 41576
rect 4674 41520 4724 41576
rect 4660 41516 4724 41520
rect 6132 41516 6196 41580
rect 980 41380 1044 41444
rect 18276 41380 18340 41444
rect 6886 41372 6950 41376
rect 6886 41316 6890 41372
rect 6890 41316 6946 41372
rect 6946 41316 6950 41372
rect 6886 41312 6950 41316
rect 6966 41372 7030 41376
rect 6966 41316 6970 41372
rect 6970 41316 7026 41372
rect 7026 41316 7030 41372
rect 6966 41312 7030 41316
rect 7046 41372 7110 41376
rect 7046 41316 7050 41372
rect 7050 41316 7106 41372
rect 7106 41316 7110 41372
rect 7046 41312 7110 41316
rect 7126 41372 7190 41376
rect 7126 41316 7130 41372
rect 7130 41316 7186 41372
rect 7186 41316 7190 41372
rect 7126 41312 7190 41316
rect 12820 41372 12884 41376
rect 12820 41316 12824 41372
rect 12824 41316 12880 41372
rect 12880 41316 12884 41372
rect 12820 41312 12884 41316
rect 12900 41372 12964 41376
rect 12900 41316 12904 41372
rect 12904 41316 12960 41372
rect 12960 41316 12964 41372
rect 12900 41312 12964 41316
rect 12980 41372 13044 41376
rect 12980 41316 12984 41372
rect 12984 41316 13040 41372
rect 13040 41316 13044 41372
rect 12980 41312 13044 41316
rect 13060 41372 13124 41376
rect 13060 41316 13064 41372
rect 13064 41316 13120 41372
rect 13120 41316 13124 41372
rect 13060 41312 13124 41316
rect 18754 41372 18818 41376
rect 18754 41316 18758 41372
rect 18758 41316 18814 41372
rect 18814 41316 18818 41372
rect 18754 41312 18818 41316
rect 18834 41372 18898 41376
rect 18834 41316 18838 41372
rect 18838 41316 18894 41372
rect 18894 41316 18898 41372
rect 18834 41312 18898 41316
rect 18914 41372 18978 41376
rect 18914 41316 18918 41372
rect 18918 41316 18974 41372
rect 18974 41316 18978 41372
rect 18914 41312 18978 41316
rect 18994 41372 19058 41376
rect 18994 41316 18998 41372
rect 18998 41316 19054 41372
rect 19054 41316 19058 41372
rect 18994 41312 19058 41316
rect 24688 41372 24752 41376
rect 24688 41316 24692 41372
rect 24692 41316 24748 41372
rect 24748 41316 24752 41372
rect 24688 41312 24752 41316
rect 24768 41372 24832 41376
rect 24768 41316 24772 41372
rect 24772 41316 24828 41372
rect 24828 41316 24832 41372
rect 24768 41312 24832 41316
rect 24848 41372 24912 41376
rect 24848 41316 24852 41372
rect 24852 41316 24908 41372
rect 24908 41316 24912 41372
rect 24848 41312 24912 41316
rect 24928 41372 24992 41376
rect 24928 41316 24932 41372
rect 24932 41316 24988 41372
rect 24988 41316 24992 41372
rect 24928 41312 24992 41316
rect 3919 40828 3983 40832
rect 3919 40772 3923 40828
rect 3923 40772 3979 40828
rect 3979 40772 3983 40828
rect 3919 40768 3983 40772
rect 3999 40828 4063 40832
rect 3999 40772 4003 40828
rect 4003 40772 4059 40828
rect 4059 40772 4063 40828
rect 3999 40768 4063 40772
rect 4079 40828 4143 40832
rect 4079 40772 4083 40828
rect 4083 40772 4139 40828
rect 4139 40772 4143 40828
rect 4079 40768 4143 40772
rect 4159 40828 4223 40832
rect 4159 40772 4163 40828
rect 4163 40772 4219 40828
rect 4219 40772 4223 40828
rect 4159 40768 4223 40772
rect 9853 40828 9917 40832
rect 9853 40772 9857 40828
rect 9857 40772 9913 40828
rect 9913 40772 9917 40828
rect 9853 40768 9917 40772
rect 9933 40828 9997 40832
rect 9933 40772 9937 40828
rect 9937 40772 9993 40828
rect 9993 40772 9997 40828
rect 9933 40768 9997 40772
rect 10013 40828 10077 40832
rect 10013 40772 10017 40828
rect 10017 40772 10073 40828
rect 10073 40772 10077 40828
rect 10013 40768 10077 40772
rect 10093 40828 10157 40832
rect 10093 40772 10097 40828
rect 10097 40772 10153 40828
rect 10153 40772 10157 40828
rect 10093 40768 10157 40772
rect 15787 40828 15851 40832
rect 15787 40772 15791 40828
rect 15791 40772 15847 40828
rect 15847 40772 15851 40828
rect 15787 40768 15851 40772
rect 15867 40828 15931 40832
rect 15867 40772 15871 40828
rect 15871 40772 15927 40828
rect 15927 40772 15931 40828
rect 15867 40768 15931 40772
rect 15947 40828 16011 40832
rect 15947 40772 15951 40828
rect 15951 40772 16007 40828
rect 16007 40772 16011 40828
rect 15947 40768 16011 40772
rect 16027 40828 16091 40832
rect 16027 40772 16031 40828
rect 16031 40772 16087 40828
rect 16087 40772 16091 40828
rect 16027 40768 16091 40772
rect 21721 40828 21785 40832
rect 21721 40772 21725 40828
rect 21725 40772 21781 40828
rect 21781 40772 21785 40828
rect 21721 40768 21785 40772
rect 21801 40828 21865 40832
rect 21801 40772 21805 40828
rect 21805 40772 21861 40828
rect 21861 40772 21865 40828
rect 21801 40768 21865 40772
rect 21881 40828 21945 40832
rect 21881 40772 21885 40828
rect 21885 40772 21941 40828
rect 21941 40772 21945 40828
rect 21881 40768 21945 40772
rect 21961 40828 22025 40832
rect 21961 40772 21965 40828
rect 21965 40772 22021 40828
rect 22021 40772 22025 40828
rect 21961 40768 22025 40772
rect 6886 40284 6950 40288
rect 6886 40228 6890 40284
rect 6890 40228 6946 40284
rect 6946 40228 6950 40284
rect 6886 40224 6950 40228
rect 6966 40284 7030 40288
rect 6966 40228 6970 40284
rect 6970 40228 7026 40284
rect 7026 40228 7030 40284
rect 6966 40224 7030 40228
rect 7046 40284 7110 40288
rect 7046 40228 7050 40284
rect 7050 40228 7106 40284
rect 7106 40228 7110 40284
rect 7046 40224 7110 40228
rect 7126 40284 7190 40288
rect 7126 40228 7130 40284
rect 7130 40228 7186 40284
rect 7186 40228 7190 40284
rect 7126 40224 7190 40228
rect 12820 40284 12884 40288
rect 12820 40228 12824 40284
rect 12824 40228 12880 40284
rect 12880 40228 12884 40284
rect 12820 40224 12884 40228
rect 12900 40284 12964 40288
rect 12900 40228 12904 40284
rect 12904 40228 12960 40284
rect 12960 40228 12964 40284
rect 12900 40224 12964 40228
rect 12980 40284 13044 40288
rect 12980 40228 12984 40284
rect 12984 40228 13040 40284
rect 13040 40228 13044 40284
rect 12980 40224 13044 40228
rect 13060 40284 13124 40288
rect 13060 40228 13064 40284
rect 13064 40228 13120 40284
rect 13120 40228 13124 40284
rect 13060 40224 13124 40228
rect 18754 40284 18818 40288
rect 18754 40228 18758 40284
rect 18758 40228 18814 40284
rect 18814 40228 18818 40284
rect 18754 40224 18818 40228
rect 18834 40284 18898 40288
rect 18834 40228 18838 40284
rect 18838 40228 18894 40284
rect 18894 40228 18898 40284
rect 18834 40224 18898 40228
rect 18914 40284 18978 40288
rect 18914 40228 18918 40284
rect 18918 40228 18974 40284
rect 18974 40228 18978 40284
rect 18914 40224 18978 40228
rect 18994 40284 19058 40288
rect 18994 40228 18998 40284
rect 18998 40228 19054 40284
rect 19054 40228 19058 40284
rect 18994 40224 19058 40228
rect 24688 40284 24752 40288
rect 24688 40228 24692 40284
rect 24692 40228 24748 40284
rect 24748 40228 24752 40284
rect 24688 40224 24752 40228
rect 24768 40284 24832 40288
rect 24768 40228 24772 40284
rect 24772 40228 24828 40284
rect 24828 40228 24832 40284
rect 24768 40224 24832 40228
rect 24848 40284 24912 40288
rect 24848 40228 24852 40284
rect 24852 40228 24908 40284
rect 24908 40228 24912 40284
rect 24848 40224 24912 40228
rect 24928 40284 24992 40288
rect 24928 40228 24932 40284
rect 24932 40228 24988 40284
rect 24988 40228 24992 40284
rect 24928 40224 24992 40228
rect 22876 40156 22940 40220
rect 3919 39740 3983 39744
rect 3919 39684 3923 39740
rect 3923 39684 3979 39740
rect 3979 39684 3983 39740
rect 3919 39680 3983 39684
rect 3999 39740 4063 39744
rect 3999 39684 4003 39740
rect 4003 39684 4059 39740
rect 4059 39684 4063 39740
rect 3999 39680 4063 39684
rect 4079 39740 4143 39744
rect 4079 39684 4083 39740
rect 4083 39684 4139 39740
rect 4139 39684 4143 39740
rect 4079 39680 4143 39684
rect 4159 39740 4223 39744
rect 4159 39684 4163 39740
rect 4163 39684 4219 39740
rect 4219 39684 4223 39740
rect 4159 39680 4223 39684
rect 9853 39740 9917 39744
rect 9853 39684 9857 39740
rect 9857 39684 9913 39740
rect 9913 39684 9917 39740
rect 9853 39680 9917 39684
rect 9933 39740 9997 39744
rect 9933 39684 9937 39740
rect 9937 39684 9993 39740
rect 9993 39684 9997 39740
rect 9933 39680 9997 39684
rect 10013 39740 10077 39744
rect 10013 39684 10017 39740
rect 10017 39684 10073 39740
rect 10073 39684 10077 39740
rect 10013 39680 10077 39684
rect 10093 39740 10157 39744
rect 10093 39684 10097 39740
rect 10097 39684 10153 39740
rect 10153 39684 10157 39740
rect 10093 39680 10157 39684
rect 15787 39740 15851 39744
rect 15787 39684 15791 39740
rect 15791 39684 15847 39740
rect 15847 39684 15851 39740
rect 15787 39680 15851 39684
rect 15867 39740 15931 39744
rect 15867 39684 15871 39740
rect 15871 39684 15927 39740
rect 15927 39684 15931 39740
rect 15867 39680 15931 39684
rect 15947 39740 16011 39744
rect 15947 39684 15951 39740
rect 15951 39684 16007 39740
rect 16007 39684 16011 39740
rect 15947 39680 16011 39684
rect 16027 39740 16091 39744
rect 16027 39684 16031 39740
rect 16031 39684 16087 39740
rect 16087 39684 16091 39740
rect 16027 39680 16091 39684
rect 21721 39740 21785 39744
rect 21721 39684 21725 39740
rect 21725 39684 21781 39740
rect 21781 39684 21785 39740
rect 21721 39680 21785 39684
rect 21801 39740 21865 39744
rect 21801 39684 21805 39740
rect 21805 39684 21861 39740
rect 21861 39684 21865 39740
rect 21801 39680 21865 39684
rect 21881 39740 21945 39744
rect 21881 39684 21885 39740
rect 21885 39684 21941 39740
rect 21941 39684 21945 39740
rect 21881 39680 21945 39684
rect 21961 39740 22025 39744
rect 21961 39684 21965 39740
rect 21965 39684 22021 39740
rect 22021 39684 22025 39740
rect 21961 39680 22025 39684
rect 6886 39196 6950 39200
rect 6886 39140 6890 39196
rect 6890 39140 6946 39196
rect 6946 39140 6950 39196
rect 6886 39136 6950 39140
rect 6966 39196 7030 39200
rect 6966 39140 6970 39196
rect 6970 39140 7026 39196
rect 7026 39140 7030 39196
rect 6966 39136 7030 39140
rect 7046 39196 7110 39200
rect 7046 39140 7050 39196
rect 7050 39140 7106 39196
rect 7106 39140 7110 39196
rect 7046 39136 7110 39140
rect 7126 39196 7190 39200
rect 7126 39140 7130 39196
rect 7130 39140 7186 39196
rect 7186 39140 7190 39196
rect 7126 39136 7190 39140
rect 12820 39196 12884 39200
rect 12820 39140 12824 39196
rect 12824 39140 12880 39196
rect 12880 39140 12884 39196
rect 12820 39136 12884 39140
rect 12900 39196 12964 39200
rect 12900 39140 12904 39196
rect 12904 39140 12960 39196
rect 12960 39140 12964 39196
rect 12900 39136 12964 39140
rect 12980 39196 13044 39200
rect 12980 39140 12984 39196
rect 12984 39140 13040 39196
rect 13040 39140 13044 39196
rect 12980 39136 13044 39140
rect 13060 39196 13124 39200
rect 13060 39140 13064 39196
rect 13064 39140 13120 39196
rect 13120 39140 13124 39196
rect 13060 39136 13124 39140
rect 18754 39196 18818 39200
rect 18754 39140 18758 39196
rect 18758 39140 18814 39196
rect 18814 39140 18818 39196
rect 18754 39136 18818 39140
rect 18834 39196 18898 39200
rect 18834 39140 18838 39196
rect 18838 39140 18894 39196
rect 18894 39140 18898 39196
rect 18834 39136 18898 39140
rect 18914 39196 18978 39200
rect 18914 39140 18918 39196
rect 18918 39140 18974 39196
rect 18974 39140 18978 39196
rect 18914 39136 18978 39140
rect 18994 39196 19058 39200
rect 18994 39140 18998 39196
rect 18998 39140 19054 39196
rect 19054 39140 19058 39196
rect 18994 39136 19058 39140
rect 24688 39196 24752 39200
rect 24688 39140 24692 39196
rect 24692 39140 24748 39196
rect 24748 39140 24752 39196
rect 24688 39136 24752 39140
rect 24768 39196 24832 39200
rect 24768 39140 24772 39196
rect 24772 39140 24828 39196
rect 24828 39140 24832 39196
rect 24768 39136 24832 39140
rect 24848 39196 24912 39200
rect 24848 39140 24852 39196
rect 24852 39140 24908 39196
rect 24908 39140 24912 39196
rect 24848 39136 24912 39140
rect 24928 39196 24992 39200
rect 24928 39140 24932 39196
rect 24932 39140 24988 39196
rect 24988 39140 24992 39196
rect 24928 39136 24992 39140
rect 2636 39068 2700 39132
rect 22508 38932 22572 38996
rect 9628 38660 9692 38724
rect 19564 38660 19628 38724
rect 3919 38652 3983 38656
rect 3919 38596 3923 38652
rect 3923 38596 3979 38652
rect 3979 38596 3983 38652
rect 3919 38592 3983 38596
rect 3999 38652 4063 38656
rect 3999 38596 4003 38652
rect 4003 38596 4059 38652
rect 4059 38596 4063 38652
rect 3999 38592 4063 38596
rect 4079 38652 4143 38656
rect 4079 38596 4083 38652
rect 4083 38596 4139 38652
rect 4139 38596 4143 38652
rect 4079 38592 4143 38596
rect 4159 38652 4223 38656
rect 4159 38596 4163 38652
rect 4163 38596 4219 38652
rect 4219 38596 4223 38652
rect 4159 38592 4223 38596
rect 9853 38652 9917 38656
rect 9853 38596 9857 38652
rect 9857 38596 9913 38652
rect 9913 38596 9917 38652
rect 9853 38592 9917 38596
rect 9933 38652 9997 38656
rect 9933 38596 9937 38652
rect 9937 38596 9993 38652
rect 9993 38596 9997 38652
rect 9933 38592 9997 38596
rect 10013 38652 10077 38656
rect 10013 38596 10017 38652
rect 10017 38596 10073 38652
rect 10073 38596 10077 38652
rect 10013 38592 10077 38596
rect 10093 38652 10157 38656
rect 10093 38596 10097 38652
rect 10097 38596 10153 38652
rect 10153 38596 10157 38652
rect 10093 38592 10157 38596
rect 15787 38652 15851 38656
rect 15787 38596 15791 38652
rect 15791 38596 15847 38652
rect 15847 38596 15851 38652
rect 15787 38592 15851 38596
rect 15867 38652 15931 38656
rect 15867 38596 15871 38652
rect 15871 38596 15927 38652
rect 15927 38596 15931 38652
rect 15867 38592 15931 38596
rect 15947 38652 16011 38656
rect 15947 38596 15951 38652
rect 15951 38596 16007 38652
rect 16007 38596 16011 38652
rect 15947 38592 16011 38596
rect 16027 38652 16091 38656
rect 16027 38596 16031 38652
rect 16031 38596 16087 38652
rect 16087 38596 16091 38652
rect 16027 38592 16091 38596
rect 21721 38652 21785 38656
rect 21721 38596 21725 38652
rect 21725 38596 21781 38652
rect 21781 38596 21785 38652
rect 21721 38592 21785 38596
rect 21801 38652 21865 38656
rect 21801 38596 21805 38652
rect 21805 38596 21861 38652
rect 21861 38596 21865 38652
rect 21801 38592 21865 38596
rect 21881 38652 21945 38656
rect 21881 38596 21885 38652
rect 21885 38596 21941 38652
rect 21941 38596 21945 38652
rect 21881 38592 21945 38596
rect 21961 38652 22025 38656
rect 21961 38596 21965 38652
rect 21965 38596 22021 38652
rect 22021 38596 22025 38652
rect 21961 38592 22025 38596
rect 2820 38116 2884 38180
rect 6886 38108 6950 38112
rect 6886 38052 6890 38108
rect 6890 38052 6946 38108
rect 6946 38052 6950 38108
rect 6886 38048 6950 38052
rect 6966 38108 7030 38112
rect 6966 38052 6970 38108
rect 6970 38052 7026 38108
rect 7026 38052 7030 38108
rect 6966 38048 7030 38052
rect 7046 38108 7110 38112
rect 7046 38052 7050 38108
rect 7050 38052 7106 38108
rect 7106 38052 7110 38108
rect 7046 38048 7110 38052
rect 7126 38108 7190 38112
rect 7126 38052 7130 38108
rect 7130 38052 7186 38108
rect 7186 38052 7190 38108
rect 7126 38048 7190 38052
rect 12820 38108 12884 38112
rect 12820 38052 12824 38108
rect 12824 38052 12880 38108
rect 12880 38052 12884 38108
rect 12820 38048 12884 38052
rect 12900 38108 12964 38112
rect 12900 38052 12904 38108
rect 12904 38052 12960 38108
rect 12960 38052 12964 38108
rect 12900 38048 12964 38052
rect 12980 38108 13044 38112
rect 12980 38052 12984 38108
rect 12984 38052 13040 38108
rect 13040 38052 13044 38108
rect 12980 38048 13044 38052
rect 13060 38108 13124 38112
rect 13060 38052 13064 38108
rect 13064 38052 13120 38108
rect 13120 38052 13124 38108
rect 13060 38048 13124 38052
rect 18754 38108 18818 38112
rect 18754 38052 18758 38108
rect 18758 38052 18814 38108
rect 18814 38052 18818 38108
rect 18754 38048 18818 38052
rect 18834 38108 18898 38112
rect 18834 38052 18838 38108
rect 18838 38052 18894 38108
rect 18894 38052 18898 38108
rect 18834 38048 18898 38052
rect 18914 38108 18978 38112
rect 18914 38052 18918 38108
rect 18918 38052 18974 38108
rect 18974 38052 18978 38108
rect 18914 38048 18978 38052
rect 18994 38108 19058 38112
rect 18994 38052 18998 38108
rect 18998 38052 19054 38108
rect 19054 38052 19058 38108
rect 18994 38048 19058 38052
rect 24688 38108 24752 38112
rect 24688 38052 24692 38108
rect 24692 38052 24748 38108
rect 24748 38052 24752 38108
rect 24688 38048 24752 38052
rect 24768 38108 24832 38112
rect 24768 38052 24772 38108
rect 24772 38052 24828 38108
rect 24828 38052 24832 38108
rect 24768 38048 24832 38052
rect 24848 38108 24912 38112
rect 24848 38052 24852 38108
rect 24852 38052 24908 38108
rect 24908 38052 24912 38108
rect 24848 38048 24912 38052
rect 24928 38108 24992 38112
rect 24928 38052 24932 38108
rect 24932 38052 24988 38108
rect 24988 38052 24992 38108
rect 24928 38048 24992 38052
rect 17908 37844 17972 37908
rect 11100 37708 11164 37772
rect 3919 37564 3983 37568
rect 3919 37508 3923 37564
rect 3923 37508 3979 37564
rect 3979 37508 3983 37564
rect 3919 37504 3983 37508
rect 3999 37564 4063 37568
rect 3999 37508 4003 37564
rect 4003 37508 4059 37564
rect 4059 37508 4063 37564
rect 3999 37504 4063 37508
rect 4079 37564 4143 37568
rect 4079 37508 4083 37564
rect 4083 37508 4139 37564
rect 4139 37508 4143 37564
rect 4079 37504 4143 37508
rect 4159 37564 4223 37568
rect 4159 37508 4163 37564
rect 4163 37508 4219 37564
rect 4219 37508 4223 37564
rect 4159 37504 4223 37508
rect 9853 37564 9917 37568
rect 9853 37508 9857 37564
rect 9857 37508 9913 37564
rect 9913 37508 9917 37564
rect 9853 37504 9917 37508
rect 9933 37564 9997 37568
rect 9933 37508 9937 37564
rect 9937 37508 9993 37564
rect 9993 37508 9997 37564
rect 9933 37504 9997 37508
rect 10013 37564 10077 37568
rect 10013 37508 10017 37564
rect 10017 37508 10073 37564
rect 10073 37508 10077 37564
rect 10013 37504 10077 37508
rect 10093 37564 10157 37568
rect 10093 37508 10097 37564
rect 10097 37508 10153 37564
rect 10153 37508 10157 37564
rect 10093 37504 10157 37508
rect 15787 37564 15851 37568
rect 15787 37508 15791 37564
rect 15791 37508 15847 37564
rect 15847 37508 15851 37564
rect 15787 37504 15851 37508
rect 15867 37564 15931 37568
rect 15867 37508 15871 37564
rect 15871 37508 15927 37564
rect 15927 37508 15931 37564
rect 15867 37504 15931 37508
rect 15947 37564 16011 37568
rect 15947 37508 15951 37564
rect 15951 37508 16007 37564
rect 16007 37508 16011 37564
rect 15947 37504 16011 37508
rect 16027 37564 16091 37568
rect 16027 37508 16031 37564
rect 16031 37508 16087 37564
rect 16087 37508 16091 37564
rect 16027 37504 16091 37508
rect 21721 37564 21785 37568
rect 21721 37508 21725 37564
rect 21725 37508 21781 37564
rect 21781 37508 21785 37564
rect 21721 37504 21785 37508
rect 21801 37564 21865 37568
rect 21801 37508 21805 37564
rect 21805 37508 21861 37564
rect 21861 37508 21865 37564
rect 21801 37504 21865 37508
rect 21881 37564 21945 37568
rect 21881 37508 21885 37564
rect 21885 37508 21941 37564
rect 21941 37508 21945 37564
rect 21881 37504 21945 37508
rect 21961 37564 22025 37568
rect 21961 37508 21965 37564
rect 21965 37508 22021 37564
rect 22021 37508 22025 37564
rect 21961 37504 22025 37508
rect 3004 37496 3068 37500
rect 3004 37440 3018 37496
rect 3018 37440 3068 37496
rect 3004 37436 3068 37440
rect 6684 37300 6748 37364
rect 8892 37300 8956 37364
rect 6886 37020 6950 37024
rect 6886 36964 6890 37020
rect 6890 36964 6946 37020
rect 6946 36964 6950 37020
rect 6886 36960 6950 36964
rect 6966 37020 7030 37024
rect 6966 36964 6970 37020
rect 6970 36964 7026 37020
rect 7026 36964 7030 37020
rect 6966 36960 7030 36964
rect 7046 37020 7110 37024
rect 7046 36964 7050 37020
rect 7050 36964 7106 37020
rect 7106 36964 7110 37020
rect 7046 36960 7110 36964
rect 7126 37020 7190 37024
rect 7126 36964 7130 37020
rect 7130 36964 7186 37020
rect 7186 36964 7190 37020
rect 7126 36960 7190 36964
rect 12820 37020 12884 37024
rect 12820 36964 12824 37020
rect 12824 36964 12880 37020
rect 12880 36964 12884 37020
rect 12820 36960 12884 36964
rect 12900 37020 12964 37024
rect 12900 36964 12904 37020
rect 12904 36964 12960 37020
rect 12960 36964 12964 37020
rect 12900 36960 12964 36964
rect 12980 37020 13044 37024
rect 12980 36964 12984 37020
rect 12984 36964 13040 37020
rect 13040 36964 13044 37020
rect 12980 36960 13044 36964
rect 13060 37020 13124 37024
rect 13060 36964 13064 37020
rect 13064 36964 13120 37020
rect 13120 36964 13124 37020
rect 13060 36960 13124 36964
rect 18754 37020 18818 37024
rect 18754 36964 18758 37020
rect 18758 36964 18814 37020
rect 18814 36964 18818 37020
rect 18754 36960 18818 36964
rect 18834 37020 18898 37024
rect 18834 36964 18838 37020
rect 18838 36964 18894 37020
rect 18894 36964 18898 37020
rect 18834 36960 18898 36964
rect 18914 37020 18978 37024
rect 18914 36964 18918 37020
rect 18918 36964 18974 37020
rect 18974 36964 18978 37020
rect 18914 36960 18978 36964
rect 18994 37020 19058 37024
rect 18994 36964 18998 37020
rect 18998 36964 19054 37020
rect 19054 36964 19058 37020
rect 18994 36960 19058 36964
rect 24688 37020 24752 37024
rect 24688 36964 24692 37020
rect 24692 36964 24748 37020
rect 24748 36964 24752 37020
rect 24688 36960 24752 36964
rect 24768 37020 24832 37024
rect 24768 36964 24772 37020
rect 24772 36964 24828 37020
rect 24828 36964 24832 37020
rect 24768 36960 24832 36964
rect 24848 37020 24912 37024
rect 24848 36964 24852 37020
rect 24852 36964 24908 37020
rect 24908 36964 24912 37020
rect 24848 36960 24912 36964
rect 24928 37020 24992 37024
rect 24928 36964 24932 37020
rect 24932 36964 24988 37020
rect 24988 36964 24992 37020
rect 24928 36960 24992 36964
rect 3919 36476 3983 36480
rect 3919 36420 3923 36476
rect 3923 36420 3979 36476
rect 3979 36420 3983 36476
rect 3919 36416 3983 36420
rect 3999 36476 4063 36480
rect 3999 36420 4003 36476
rect 4003 36420 4059 36476
rect 4059 36420 4063 36476
rect 3999 36416 4063 36420
rect 4079 36476 4143 36480
rect 4079 36420 4083 36476
rect 4083 36420 4139 36476
rect 4139 36420 4143 36476
rect 4079 36416 4143 36420
rect 4159 36476 4223 36480
rect 4159 36420 4163 36476
rect 4163 36420 4219 36476
rect 4219 36420 4223 36476
rect 4159 36416 4223 36420
rect 9853 36476 9917 36480
rect 9853 36420 9857 36476
rect 9857 36420 9913 36476
rect 9913 36420 9917 36476
rect 9853 36416 9917 36420
rect 9933 36476 9997 36480
rect 9933 36420 9937 36476
rect 9937 36420 9993 36476
rect 9993 36420 9997 36476
rect 9933 36416 9997 36420
rect 10013 36476 10077 36480
rect 10013 36420 10017 36476
rect 10017 36420 10073 36476
rect 10073 36420 10077 36476
rect 10013 36416 10077 36420
rect 10093 36476 10157 36480
rect 10093 36420 10097 36476
rect 10097 36420 10153 36476
rect 10153 36420 10157 36476
rect 10093 36416 10157 36420
rect 15787 36476 15851 36480
rect 15787 36420 15791 36476
rect 15791 36420 15847 36476
rect 15847 36420 15851 36476
rect 15787 36416 15851 36420
rect 15867 36476 15931 36480
rect 15867 36420 15871 36476
rect 15871 36420 15927 36476
rect 15927 36420 15931 36476
rect 15867 36416 15931 36420
rect 15947 36476 16011 36480
rect 15947 36420 15951 36476
rect 15951 36420 16007 36476
rect 16007 36420 16011 36476
rect 15947 36416 16011 36420
rect 16027 36476 16091 36480
rect 16027 36420 16031 36476
rect 16031 36420 16087 36476
rect 16087 36420 16091 36476
rect 16027 36416 16091 36420
rect 21721 36476 21785 36480
rect 21721 36420 21725 36476
rect 21725 36420 21781 36476
rect 21781 36420 21785 36476
rect 21721 36416 21785 36420
rect 21801 36476 21865 36480
rect 21801 36420 21805 36476
rect 21805 36420 21861 36476
rect 21861 36420 21865 36476
rect 21801 36416 21865 36420
rect 21881 36476 21945 36480
rect 21881 36420 21885 36476
rect 21885 36420 21941 36476
rect 21941 36420 21945 36476
rect 21881 36416 21945 36420
rect 21961 36476 22025 36480
rect 21961 36420 21965 36476
rect 21965 36420 22021 36476
rect 22021 36420 22025 36476
rect 21961 36416 22025 36420
rect 2452 36076 2516 36140
rect 3004 36076 3068 36140
rect 3740 35940 3804 36004
rect 22876 35940 22940 36004
rect 6886 35932 6950 35936
rect 6886 35876 6890 35932
rect 6890 35876 6946 35932
rect 6946 35876 6950 35932
rect 6886 35872 6950 35876
rect 6966 35932 7030 35936
rect 6966 35876 6970 35932
rect 6970 35876 7026 35932
rect 7026 35876 7030 35932
rect 6966 35872 7030 35876
rect 7046 35932 7110 35936
rect 7046 35876 7050 35932
rect 7050 35876 7106 35932
rect 7106 35876 7110 35932
rect 7046 35872 7110 35876
rect 7126 35932 7190 35936
rect 7126 35876 7130 35932
rect 7130 35876 7186 35932
rect 7186 35876 7190 35932
rect 7126 35872 7190 35876
rect 12820 35932 12884 35936
rect 12820 35876 12824 35932
rect 12824 35876 12880 35932
rect 12880 35876 12884 35932
rect 12820 35872 12884 35876
rect 12900 35932 12964 35936
rect 12900 35876 12904 35932
rect 12904 35876 12960 35932
rect 12960 35876 12964 35932
rect 12900 35872 12964 35876
rect 12980 35932 13044 35936
rect 12980 35876 12984 35932
rect 12984 35876 13040 35932
rect 13040 35876 13044 35932
rect 12980 35872 13044 35876
rect 13060 35932 13124 35936
rect 13060 35876 13064 35932
rect 13064 35876 13120 35932
rect 13120 35876 13124 35932
rect 13060 35872 13124 35876
rect 18754 35932 18818 35936
rect 18754 35876 18758 35932
rect 18758 35876 18814 35932
rect 18814 35876 18818 35932
rect 18754 35872 18818 35876
rect 18834 35932 18898 35936
rect 18834 35876 18838 35932
rect 18838 35876 18894 35932
rect 18894 35876 18898 35932
rect 18834 35872 18898 35876
rect 18914 35932 18978 35936
rect 18914 35876 18918 35932
rect 18918 35876 18974 35932
rect 18974 35876 18978 35932
rect 18914 35872 18978 35876
rect 18994 35932 19058 35936
rect 18994 35876 18998 35932
rect 18998 35876 19054 35932
rect 19054 35876 19058 35932
rect 18994 35872 19058 35876
rect 24688 35932 24752 35936
rect 24688 35876 24692 35932
rect 24692 35876 24748 35932
rect 24748 35876 24752 35932
rect 24688 35872 24752 35876
rect 24768 35932 24832 35936
rect 24768 35876 24772 35932
rect 24772 35876 24828 35932
rect 24828 35876 24832 35932
rect 24768 35872 24832 35876
rect 24848 35932 24912 35936
rect 24848 35876 24852 35932
rect 24852 35876 24908 35932
rect 24908 35876 24912 35932
rect 24848 35872 24912 35876
rect 24928 35932 24992 35936
rect 24928 35876 24932 35932
rect 24932 35876 24988 35932
rect 24988 35876 24992 35932
rect 24928 35872 24992 35876
rect 10548 35804 10612 35868
rect 6684 35396 6748 35460
rect 3919 35388 3983 35392
rect 3919 35332 3923 35388
rect 3923 35332 3979 35388
rect 3979 35332 3983 35388
rect 3919 35328 3983 35332
rect 3999 35388 4063 35392
rect 3999 35332 4003 35388
rect 4003 35332 4059 35388
rect 4059 35332 4063 35388
rect 3999 35328 4063 35332
rect 4079 35388 4143 35392
rect 4079 35332 4083 35388
rect 4083 35332 4139 35388
rect 4139 35332 4143 35388
rect 4079 35328 4143 35332
rect 4159 35388 4223 35392
rect 4159 35332 4163 35388
rect 4163 35332 4219 35388
rect 4219 35332 4223 35388
rect 4159 35328 4223 35332
rect 9853 35388 9917 35392
rect 9853 35332 9857 35388
rect 9857 35332 9913 35388
rect 9913 35332 9917 35388
rect 9853 35328 9917 35332
rect 9933 35388 9997 35392
rect 9933 35332 9937 35388
rect 9937 35332 9993 35388
rect 9993 35332 9997 35388
rect 9933 35328 9997 35332
rect 10013 35388 10077 35392
rect 10013 35332 10017 35388
rect 10017 35332 10073 35388
rect 10073 35332 10077 35388
rect 10013 35328 10077 35332
rect 10093 35388 10157 35392
rect 10093 35332 10097 35388
rect 10097 35332 10153 35388
rect 10153 35332 10157 35388
rect 10093 35328 10157 35332
rect 15787 35388 15851 35392
rect 15787 35332 15791 35388
rect 15791 35332 15847 35388
rect 15847 35332 15851 35388
rect 15787 35328 15851 35332
rect 15867 35388 15931 35392
rect 15867 35332 15871 35388
rect 15871 35332 15927 35388
rect 15927 35332 15931 35388
rect 15867 35328 15931 35332
rect 15947 35388 16011 35392
rect 15947 35332 15951 35388
rect 15951 35332 16007 35388
rect 16007 35332 16011 35388
rect 15947 35328 16011 35332
rect 16027 35388 16091 35392
rect 16027 35332 16031 35388
rect 16031 35332 16087 35388
rect 16087 35332 16091 35388
rect 16027 35328 16091 35332
rect 21721 35388 21785 35392
rect 21721 35332 21725 35388
rect 21725 35332 21781 35388
rect 21781 35332 21785 35388
rect 21721 35328 21785 35332
rect 21801 35388 21865 35392
rect 21801 35332 21805 35388
rect 21805 35332 21861 35388
rect 21861 35332 21865 35388
rect 21801 35328 21865 35332
rect 21881 35388 21945 35392
rect 21881 35332 21885 35388
rect 21885 35332 21941 35388
rect 21941 35332 21945 35388
rect 21881 35328 21945 35332
rect 21961 35388 22025 35392
rect 21961 35332 21965 35388
rect 21965 35332 22021 35388
rect 22021 35332 22025 35388
rect 21961 35328 22025 35332
rect 11468 35260 11532 35324
rect 5580 35124 5644 35188
rect 13308 34988 13372 35052
rect 6886 34844 6950 34848
rect 6886 34788 6890 34844
rect 6890 34788 6946 34844
rect 6946 34788 6950 34844
rect 6886 34784 6950 34788
rect 6966 34844 7030 34848
rect 6966 34788 6970 34844
rect 6970 34788 7026 34844
rect 7026 34788 7030 34844
rect 6966 34784 7030 34788
rect 7046 34844 7110 34848
rect 7046 34788 7050 34844
rect 7050 34788 7106 34844
rect 7106 34788 7110 34844
rect 7046 34784 7110 34788
rect 7126 34844 7190 34848
rect 7126 34788 7130 34844
rect 7130 34788 7186 34844
rect 7186 34788 7190 34844
rect 7126 34784 7190 34788
rect 12820 34844 12884 34848
rect 12820 34788 12824 34844
rect 12824 34788 12880 34844
rect 12880 34788 12884 34844
rect 12820 34784 12884 34788
rect 12900 34844 12964 34848
rect 12900 34788 12904 34844
rect 12904 34788 12960 34844
rect 12960 34788 12964 34844
rect 12900 34784 12964 34788
rect 12980 34844 13044 34848
rect 12980 34788 12984 34844
rect 12984 34788 13040 34844
rect 13040 34788 13044 34844
rect 12980 34784 13044 34788
rect 13060 34844 13124 34848
rect 13060 34788 13064 34844
rect 13064 34788 13120 34844
rect 13120 34788 13124 34844
rect 13060 34784 13124 34788
rect 18754 34844 18818 34848
rect 18754 34788 18758 34844
rect 18758 34788 18814 34844
rect 18814 34788 18818 34844
rect 18754 34784 18818 34788
rect 18834 34844 18898 34848
rect 18834 34788 18838 34844
rect 18838 34788 18894 34844
rect 18894 34788 18898 34844
rect 18834 34784 18898 34788
rect 18914 34844 18978 34848
rect 18914 34788 18918 34844
rect 18918 34788 18974 34844
rect 18974 34788 18978 34844
rect 18914 34784 18978 34788
rect 18994 34844 19058 34848
rect 18994 34788 18998 34844
rect 18998 34788 19054 34844
rect 19054 34788 19058 34844
rect 18994 34784 19058 34788
rect 24688 34844 24752 34848
rect 24688 34788 24692 34844
rect 24692 34788 24748 34844
rect 24748 34788 24752 34844
rect 24688 34784 24752 34788
rect 24768 34844 24832 34848
rect 24768 34788 24772 34844
rect 24772 34788 24828 34844
rect 24828 34788 24832 34844
rect 24768 34784 24832 34788
rect 24848 34844 24912 34848
rect 24848 34788 24852 34844
rect 24852 34788 24908 34844
rect 24908 34788 24912 34844
rect 24848 34784 24912 34788
rect 24928 34844 24992 34848
rect 24928 34788 24932 34844
rect 24932 34788 24988 34844
rect 24988 34788 24992 34844
rect 24928 34784 24992 34788
rect 2084 34640 2148 34644
rect 2084 34584 2098 34640
rect 2098 34584 2148 34640
rect 2084 34580 2148 34584
rect 4476 34580 4540 34644
rect 5396 34444 5460 34508
rect 3919 34300 3983 34304
rect 3919 34244 3923 34300
rect 3923 34244 3979 34300
rect 3979 34244 3983 34300
rect 3919 34240 3983 34244
rect 3999 34300 4063 34304
rect 3999 34244 4003 34300
rect 4003 34244 4059 34300
rect 4059 34244 4063 34300
rect 3999 34240 4063 34244
rect 4079 34300 4143 34304
rect 4079 34244 4083 34300
rect 4083 34244 4139 34300
rect 4139 34244 4143 34300
rect 4079 34240 4143 34244
rect 4159 34300 4223 34304
rect 4159 34244 4163 34300
rect 4163 34244 4219 34300
rect 4219 34244 4223 34300
rect 4159 34240 4223 34244
rect 9853 34300 9917 34304
rect 9853 34244 9857 34300
rect 9857 34244 9913 34300
rect 9913 34244 9917 34300
rect 9853 34240 9917 34244
rect 9933 34300 9997 34304
rect 9933 34244 9937 34300
rect 9937 34244 9993 34300
rect 9993 34244 9997 34300
rect 9933 34240 9997 34244
rect 10013 34300 10077 34304
rect 10013 34244 10017 34300
rect 10017 34244 10073 34300
rect 10073 34244 10077 34300
rect 10013 34240 10077 34244
rect 10093 34300 10157 34304
rect 10093 34244 10097 34300
rect 10097 34244 10153 34300
rect 10153 34244 10157 34300
rect 10093 34240 10157 34244
rect 15787 34300 15851 34304
rect 15787 34244 15791 34300
rect 15791 34244 15847 34300
rect 15847 34244 15851 34300
rect 15787 34240 15851 34244
rect 15867 34300 15931 34304
rect 15867 34244 15871 34300
rect 15871 34244 15927 34300
rect 15927 34244 15931 34300
rect 15867 34240 15931 34244
rect 15947 34300 16011 34304
rect 15947 34244 15951 34300
rect 15951 34244 16007 34300
rect 16007 34244 16011 34300
rect 15947 34240 16011 34244
rect 16027 34300 16091 34304
rect 16027 34244 16031 34300
rect 16031 34244 16087 34300
rect 16087 34244 16091 34300
rect 16027 34240 16091 34244
rect 21721 34300 21785 34304
rect 21721 34244 21725 34300
rect 21725 34244 21781 34300
rect 21781 34244 21785 34300
rect 21721 34240 21785 34244
rect 21801 34300 21865 34304
rect 21801 34244 21805 34300
rect 21805 34244 21861 34300
rect 21861 34244 21865 34300
rect 21801 34240 21865 34244
rect 21881 34300 21945 34304
rect 21881 34244 21885 34300
rect 21885 34244 21941 34300
rect 21941 34244 21945 34300
rect 21881 34240 21945 34244
rect 21961 34300 22025 34304
rect 21961 34244 21965 34300
rect 21965 34244 22021 34300
rect 22021 34244 22025 34300
rect 21961 34240 22025 34244
rect 4660 34036 4724 34100
rect 3004 33764 3068 33828
rect 6886 33756 6950 33760
rect 6886 33700 6890 33756
rect 6890 33700 6946 33756
rect 6946 33700 6950 33756
rect 6886 33696 6950 33700
rect 6966 33756 7030 33760
rect 6966 33700 6970 33756
rect 6970 33700 7026 33756
rect 7026 33700 7030 33756
rect 6966 33696 7030 33700
rect 7046 33756 7110 33760
rect 7046 33700 7050 33756
rect 7050 33700 7106 33756
rect 7106 33700 7110 33756
rect 7046 33696 7110 33700
rect 7126 33756 7190 33760
rect 7126 33700 7130 33756
rect 7130 33700 7186 33756
rect 7186 33700 7190 33756
rect 7126 33696 7190 33700
rect 12820 33756 12884 33760
rect 12820 33700 12824 33756
rect 12824 33700 12880 33756
rect 12880 33700 12884 33756
rect 12820 33696 12884 33700
rect 12900 33756 12964 33760
rect 12900 33700 12904 33756
rect 12904 33700 12960 33756
rect 12960 33700 12964 33756
rect 12900 33696 12964 33700
rect 12980 33756 13044 33760
rect 12980 33700 12984 33756
rect 12984 33700 13040 33756
rect 13040 33700 13044 33756
rect 12980 33696 13044 33700
rect 13060 33756 13124 33760
rect 13060 33700 13064 33756
rect 13064 33700 13120 33756
rect 13120 33700 13124 33756
rect 13060 33696 13124 33700
rect 18754 33756 18818 33760
rect 18754 33700 18758 33756
rect 18758 33700 18814 33756
rect 18814 33700 18818 33756
rect 18754 33696 18818 33700
rect 18834 33756 18898 33760
rect 18834 33700 18838 33756
rect 18838 33700 18894 33756
rect 18894 33700 18898 33756
rect 18834 33696 18898 33700
rect 18914 33756 18978 33760
rect 18914 33700 18918 33756
rect 18918 33700 18974 33756
rect 18974 33700 18978 33756
rect 18914 33696 18978 33700
rect 18994 33756 19058 33760
rect 18994 33700 18998 33756
rect 18998 33700 19054 33756
rect 19054 33700 19058 33756
rect 18994 33696 19058 33700
rect 24688 33756 24752 33760
rect 24688 33700 24692 33756
rect 24692 33700 24748 33756
rect 24748 33700 24752 33756
rect 24688 33696 24752 33700
rect 24768 33756 24832 33760
rect 24768 33700 24772 33756
rect 24772 33700 24828 33756
rect 24828 33700 24832 33756
rect 24768 33696 24832 33700
rect 24848 33756 24912 33760
rect 24848 33700 24852 33756
rect 24852 33700 24908 33756
rect 24908 33700 24912 33756
rect 24848 33696 24912 33700
rect 24928 33756 24992 33760
rect 24928 33700 24932 33756
rect 24932 33700 24988 33756
rect 24988 33700 24992 33756
rect 24928 33696 24992 33700
rect 3740 33628 3804 33692
rect 10916 33492 10980 33556
rect 2452 33356 2516 33420
rect 19932 33356 19996 33420
rect 19748 33220 19812 33284
rect 3919 33212 3983 33216
rect 3919 33156 3923 33212
rect 3923 33156 3979 33212
rect 3979 33156 3983 33212
rect 3919 33152 3983 33156
rect 3999 33212 4063 33216
rect 3999 33156 4003 33212
rect 4003 33156 4059 33212
rect 4059 33156 4063 33212
rect 3999 33152 4063 33156
rect 4079 33212 4143 33216
rect 4079 33156 4083 33212
rect 4083 33156 4139 33212
rect 4139 33156 4143 33212
rect 4079 33152 4143 33156
rect 4159 33212 4223 33216
rect 4159 33156 4163 33212
rect 4163 33156 4219 33212
rect 4219 33156 4223 33212
rect 4159 33152 4223 33156
rect 9853 33212 9917 33216
rect 9853 33156 9857 33212
rect 9857 33156 9913 33212
rect 9913 33156 9917 33212
rect 9853 33152 9917 33156
rect 9933 33212 9997 33216
rect 9933 33156 9937 33212
rect 9937 33156 9993 33212
rect 9993 33156 9997 33212
rect 9933 33152 9997 33156
rect 10013 33212 10077 33216
rect 10013 33156 10017 33212
rect 10017 33156 10073 33212
rect 10073 33156 10077 33212
rect 10013 33152 10077 33156
rect 10093 33212 10157 33216
rect 10093 33156 10097 33212
rect 10097 33156 10153 33212
rect 10153 33156 10157 33212
rect 10093 33152 10157 33156
rect 15787 33212 15851 33216
rect 15787 33156 15791 33212
rect 15791 33156 15847 33212
rect 15847 33156 15851 33212
rect 15787 33152 15851 33156
rect 15867 33212 15931 33216
rect 15867 33156 15871 33212
rect 15871 33156 15927 33212
rect 15927 33156 15931 33212
rect 15867 33152 15931 33156
rect 15947 33212 16011 33216
rect 15947 33156 15951 33212
rect 15951 33156 16007 33212
rect 16007 33156 16011 33212
rect 15947 33152 16011 33156
rect 16027 33212 16091 33216
rect 16027 33156 16031 33212
rect 16031 33156 16087 33212
rect 16087 33156 16091 33212
rect 16027 33152 16091 33156
rect 21721 33212 21785 33216
rect 21721 33156 21725 33212
rect 21725 33156 21781 33212
rect 21781 33156 21785 33212
rect 21721 33152 21785 33156
rect 21801 33212 21865 33216
rect 21801 33156 21805 33212
rect 21805 33156 21861 33212
rect 21861 33156 21865 33212
rect 21801 33152 21865 33156
rect 21881 33212 21945 33216
rect 21881 33156 21885 33212
rect 21885 33156 21941 33212
rect 21941 33156 21945 33212
rect 21881 33152 21945 33156
rect 21961 33212 22025 33216
rect 21961 33156 21965 33212
rect 21965 33156 22021 33212
rect 22021 33156 22025 33212
rect 21961 33152 22025 33156
rect 9628 32948 9692 33012
rect 10364 32812 10428 32876
rect 6886 32668 6950 32672
rect 6886 32612 6890 32668
rect 6890 32612 6946 32668
rect 6946 32612 6950 32668
rect 6886 32608 6950 32612
rect 6966 32668 7030 32672
rect 6966 32612 6970 32668
rect 6970 32612 7026 32668
rect 7026 32612 7030 32668
rect 6966 32608 7030 32612
rect 7046 32668 7110 32672
rect 7046 32612 7050 32668
rect 7050 32612 7106 32668
rect 7106 32612 7110 32668
rect 7046 32608 7110 32612
rect 7126 32668 7190 32672
rect 7126 32612 7130 32668
rect 7130 32612 7186 32668
rect 7186 32612 7190 32668
rect 7126 32608 7190 32612
rect 12820 32668 12884 32672
rect 12820 32612 12824 32668
rect 12824 32612 12880 32668
rect 12880 32612 12884 32668
rect 12820 32608 12884 32612
rect 12900 32668 12964 32672
rect 12900 32612 12904 32668
rect 12904 32612 12960 32668
rect 12960 32612 12964 32668
rect 12900 32608 12964 32612
rect 12980 32668 13044 32672
rect 12980 32612 12984 32668
rect 12984 32612 13040 32668
rect 13040 32612 13044 32668
rect 12980 32608 13044 32612
rect 13060 32668 13124 32672
rect 13060 32612 13064 32668
rect 13064 32612 13120 32668
rect 13120 32612 13124 32668
rect 13060 32608 13124 32612
rect 18754 32668 18818 32672
rect 18754 32612 18758 32668
rect 18758 32612 18814 32668
rect 18814 32612 18818 32668
rect 18754 32608 18818 32612
rect 18834 32668 18898 32672
rect 18834 32612 18838 32668
rect 18838 32612 18894 32668
rect 18894 32612 18898 32668
rect 18834 32608 18898 32612
rect 18914 32668 18978 32672
rect 18914 32612 18918 32668
rect 18918 32612 18974 32668
rect 18974 32612 18978 32668
rect 18914 32608 18978 32612
rect 18994 32668 19058 32672
rect 18994 32612 18998 32668
rect 18998 32612 19054 32668
rect 19054 32612 19058 32668
rect 18994 32608 19058 32612
rect 24688 32668 24752 32672
rect 24688 32612 24692 32668
rect 24692 32612 24748 32668
rect 24748 32612 24752 32668
rect 24688 32608 24752 32612
rect 24768 32668 24832 32672
rect 24768 32612 24772 32668
rect 24772 32612 24828 32668
rect 24828 32612 24832 32668
rect 24768 32608 24832 32612
rect 24848 32668 24912 32672
rect 24848 32612 24852 32668
rect 24852 32612 24908 32668
rect 24908 32612 24912 32668
rect 24848 32608 24912 32612
rect 24928 32668 24992 32672
rect 24928 32612 24932 32668
rect 24932 32612 24988 32668
rect 24988 32612 24992 32668
rect 24928 32608 24992 32612
rect 3556 32268 3620 32332
rect 3919 32124 3983 32128
rect 3919 32068 3923 32124
rect 3923 32068 3979 32124
rect 3979 32068 3983 32124
rect 3919 32064 3983 32068
rect 3999 32124 4063 32128
rect 3999 32068 4003 32124
rect 4003 32068 4059 32124
rect 4059 32068 4063 32124
rect 3999 32064 4063 32068
rect 4079 32124 4143 32128
rect 4079 32068 4083 32124
rect 4083 32068 4139 32124
rect 4139 32068 4143 32124
rect 4079 32064 4143 32068
rect 4159 32124 4223 32128
rect 4159 32068 4163 32124
rect 4163 32068 4219 32124
rect 4219 32068 4223 32124
rect 4159 32064 4223 32068
rect 9853 32124 9917 32128
rect 9853 32068 9857 32124
rect 9857 32068 9913 32124
rect 9913 32068 9917 32124
rect 9853 32064 9917 32068
rect 9933 32124 9997 32128
rect 9933 32068 9937 32124
rect 9937 32068 9993 32124
rect 9993 32068 9997 32124
rect 9933 32064 9997 32068
rect 10013 32124 10077 32128
rect 10013 32068 10017 32124
rect 10017 32068 10073 32124
rect 10073 32068 10077 32124
rect 10013 32064 10077 32068
rect 10093 32124 10157 32128
rect 10093 32068 10097 32124
rect 10097 32068 10153 32124
rect 10153 32068 10157 32124
rect 10093 32064 10157 32068
rect 15787 32124 15851 32128
rect 15787 32068 15791 32124
rect 15791 32068 15847 32124
rect 15847 32068 15851 32124
rect 15787 32064 15851 32068
rect 15867 32124 15931 32128
rect 15867 32068 15871 32124
rect 15871 32068 15927 32124
rect 15927 32068 15931 32124
rect 15867 32064 15931 32068
rect 15947 32124 16011 32128
rect 15947 32068 15951 32124
rect 15951 32068 16007 32124
rect 16007 32068 16011 32124
rect 15947 32064 16011 32068
rect 16027 32124 16091 32128
rect 16027 32068 16031 32124
rect 16031 32068 16087 32124
rect 16087 32068 16091 32124
rect 16027 32064 16091 32068
rect 21721 32124 21785 32128
rect 21721 32068 21725 32124
rect 21725 32068 21781 32124
rect 21781 32068 21785 32124
rect 21721 32064 21785 32068
rect 21801 32124 21865 32128
rect 21801 32068 21805 32124
rect 21805 32068 21861 32124
rect 21861 32068 21865 32124
rect 21801 32064 21865 32068
rect 21881 32124 21945 32128
rect 21881 32068 21885 32124
rect 21885 32068 21941 32124
rect 21941 32068 21945 32124
rect 21881 32064 21945 32068
rect 21961 32124 22025 32128
rect 21961 32068 21965 32124
rect 21965 32068 22021 32124
rect 22021 32068 22025 32124
rect 21961 32064 22025 32068
rect 12020 31724 12084 31788
rect 6886 31580 6950 31584
rect 6886 31524 6890 31580
rect 6890 31524 6946 31580
rect 6946 31524 6950 31580
rect 6886 31520 6950 31524
rect 6966 31580 7030 31584
rect 6966 31524 6970 31580
rect 6970 31524 7026 31580
rect 7026 31524 7030 31580
rect 6966 31520 7030 31524
rect 7046 31580 7110 31584
rect 7046 31524 7050 31580
rect 7050 31524 7106 31580
rect 7106 31524 7110 31580
rect 7046 31520 7110 31524
rect 7126 31580 7190 31584
rect 7126 31524 7130 31580
rect 7130 31524 7186 31580
rect 7186 31524 7190 31580
rect 7126 31520 7190 31524
rect 12820 31580 12884 31584
rect 12820 31524 12824 31580
rect 12824 31524 12880 31580
rect 12880 31524 12884 31580
rect 12820 31520 12884 31524
rect 12900 31580 12964 31584
rect 12900 31524 12904 31580
rect 12904 31524 12960 31580
rect 12960 31524 12964 31580
rect 12900 31520 12964 31524
rect 12980 31580 13044 31584
rect 12980 31524 12984 31580
rect 12984 31524 13040 31580
rect 13040 31524 13044 31580
rect 12980 31520 13044 31524
rect 13060 31580 13124 31584
rect 13060 31524 13064 31580
rect 13064 31524 13120 31580
rect 13120 31524 13124 31580
rect 13060 31520 13124 31524
rect 18754 31580 18818 31584
rect 18754 31524 18758 31580
rect 18758 31524 18814 31580
rect 18814 31524 18818 31580
rect 18754 31520 18818 31524
rect 18834 31580 18898 31584
rect 18834 31524 18838 31580
rect 18838 31524 18894 31580
rect 18894 31524 18898 31580
rect 18834 31520 18898 31524
rect 18914 31580 18978 31584
rect 18914 31524 18918 31580
rect 18918 31524 18974 31580
rect 18974 31524 18978 31580
rect 18914 31520 18978 31524
rect 18994 31580 19058 31584
rect 18994 31524 18998 31580
rect 18998 31524 19054 31580
rect 19054 31524 19058 31580
rect 18994 31520 19058 31524
rect 24688 31580 24752 31584
rect 24688 31524 24692 31580
rect 24692 31524 24748 31580
rect 24748 31524 24752 31580
rect 24688 31520 24752 31524
rect 24768 31580 24832 31584
rect 24768 31524 24772 31580
rect 24772 31524 24828 31580
rect 24828 31524 24832 31580
rect 24768 31520 24832 31524
rect 24848 31580 24912 31584
rect 24848 31524 24852 31580
rect 24852 31524 24908 31580
rect 24908 31524 24912 31580
rect 24848 31520 24912 31524
rect 24928 31580 24992 31584
rect 24928 31524 24932 31580
rect 24932 31524 24988 31580
rect 24988 31524 24992 31580
rect 24928 31520 24992 31524
rect 4660 31316 4724 31380
rect 7420 31316 7484 31380
rect 7604 31180 7668 31244
rect 21036 31180 21100 31244
rect 3919 31036 3983 31040
rect 3919 30980 3923 31036
rect 3923 30980 3979 31036
rect 3979 30980 3983 31036
rect 3919 30976 3983 30980
rect 3999 31036 4063 31040
rect 3999 30980 4003 31036
rect 4003 30980 4059 31036
rect 4059 30980 4063 31036
rect 3999 30976 4063 30980
rect 4079 31036 4143 31040
rect 4079 30980 4083 31036
rect 4083 30980 4139 31036
rect 4139 30980 4143 31036
rect 4079 30976 4143 30980
rect 4159 31036 4223 31040
rect 4159 30980 4163 31036
rect 4163 30980 4219 31036
rect 4219 30980 4223 31036
rect 4159 30976 4223 30980
rect 9853 31036 9917 31040
rect 9853 30980 9857 31036
rect 9857 30980 9913 31036
rect 9913 30980 9917 31036
rect 9853 30976 9917 30980
rect 9933 31036 9997 31040
rect 9933 30980 9937 31036
rect 9937 30980 9993 31036
rect 9993 30980 9997 31036
rect 9933 30976 9997 30980
rect 10013 31036 10077 31040
rect 10013 30980 10017 31036
rect 10017 30980 10073 31036
rect 10073 30980 10077 31036
rect 10013 30976 10077 30980
rect 10093 31036 10157 31040
rect 10093 30980 10097 31036
rect 10097 30980 10153 31036
rect 10153 30980 10157 31036
rect 10093 30976 10157 30980
rect 15787 31036 15851 31040
rect 15787 30980 15791 31036
rect 15791 30980 15847 31036
rect 15847 30980 15851 31036
rect 15787 30976 15851 30980
rect 15867 31036 15931 31040
rect 15867 30980 15871 31036
rect 15871 30980 15927 31036
rect 15927 30980 15931 31036
rect 15867 30976 15931 30980
rect 15947 31036 16011 31040
rect 15947 30980 15951 31036
rect 15951 30980 16007 31036
rect 16007 30980 16011 31036
rect 15947 30976 16011 30980
rect 16027 31036 16091 31040
rect 16027 30980 16031 31036
rect 16031 30980 16087 31036
rect 16087 30980 16091 31036
rect 16027 30976 16091 30980
rect 21721 31036 21785 31040
rect 21721 30980 21725 31036
rect 21725 30980 21781 31036
rect 21781 30980 21785 31036
rect 21721 30976 21785 30980
rect 21801 31036 21865 31040
rect 21801 30980 21805 31036
rect 21805 30980 21861 31036
rect 21861 30980 21865 31036
rect 21801 30976 21865 30980
rect 21881 31036 21945 31040
rect 21881 30980 21885 31036
rect 21885 30980 21941 31036
rect 21941 30980 21945 31036
rect 21881 30976 21945 30980
rect 21961 31036 22025 31040
rect 21961 30980 21965 31036
rect 21965 30980 22021 31036
rect 22021 30980 22025 31036
rect 21961 30976 22025 30980
rect 2268 30636 2332 30700
rect 11468 30636 11532 30700
rect 6886 30492 6950 30496
rect 6886 30436 6890 30492
rect 6890 30436 6946 30492
rect 6946 30436 6950 30492
rect 6886 30432 6950 30436
rect 6966 30492 7030 30496
rect 6966 30436 6970 30492
rect 6970 30436 7026 30492
rect 7026 30436 7030 30492
rect 6966 30432 7030 30436
rect 7046 30492 7110 30496
rect 7046 30436 7050 30492
rect 7050 30436 7106 30492
rect 7106 30436 7110 30492
rect 7046 30432 7110 30436
rect 7126 30492 7190 30496
rect 7126 30436 7130 30492
rect 7130 30436 7186 30492
rect 7186 30436 7190 30492
rect 7126 30432 7190 30436
rect 12820 30492 12884 30496
rect 12820 30436 12824 30492
rect 12824 30436 12880 30492
rect 12880 30436 12884 30492
rect 12820 30432 12884 30436
rect 12900 30492 12964 30496
rect 12900 30436 12904 30492
rect 12904 30436 12960 30492
rect 12960 30436 12964 30492
rect 12900 30432 12964 30436
rect 12980 30492 13044 30496
rect 12980 30436 12984 30492
rect 12984 30436 13040 30492
rect 13040 30436 13044 30492
rect 12980 30432 13044 30436
rect 13060 30492 13124 30496
rect 13060 30436 13064 30492
rect 13064 30436 13120 30492
rect 13120 30436 13124 30492
rect 13060 30432 13124 30436
rect 18754 30492 18818 30496
rect 18754 30436 18758 30492
rect 18758 30436 18814 30492
rect 18814 30436 18818 30492
rect 18754 30432 18818 30436
rect 18834 30492 18898 30496
rect 18834 30436 18838 30492
rect 18838 30436 18894 30492
rect 18894 30436 18898 30492
rect 18834 30432 18898 30436
rect 18914 30492 18978 30496
rect 18914 30436 18918 30492
rect 18918 30436 18974 30492
rect 18974 30436 18978 30492
rect 18914 30432 18978 30436
rect 18994 30492 19058 30496
rect 18994 30436 18998 30492
rect 18998 30436 19054 30492
rect 19054 30436 19058 30492
rect 18994 30432 19058 30436
rect 24688 30492 24752 30496
rect 24688 30436 24692 30492
rect 24692 30436 24748 30492
rect 24748 30436 24752 30492
rect 24688 30432 24752 30436
rect 24768 30492 24832 30496
rect 24768 30436 24772 30492
rect 24772 30436 24828 30492
rect 24828 30436 24832 30492
rect 24768 30432 24832 30436
rect 24848 30492 24912 30496
rect 24848 30436 24852 30492
rect 24852 30436 24908 30492
rect 24908 30436 24912 30492
rect 24848 30432 24912 30436
rect 24928 30492 24992 30496
rect 24928 30436 24932 30492
rect 24932 30436 24988 30492
rect 24988 30436 24992 30492
rect 24928 30432 24992 30436
rect 3372 30364 3436 30428
rect 4844 30424 4908 30428
rect 4844 30368 4894 30424
rect 4894 30368 4908 30424
rect 4844 30364 4908 30368
rect 4476 30228 4540 30292
rect 21588 30364 21652 30428
rect 3919 29948 3983 29952
rect 3919 29892 3923 29948
rect 3923 29892 3979 29948
rect 3979 29892 3983 29948
rect 3919 29888 3983 29892
rect 3999 29948 4063 29952
rect 3999 29892 4003 29948
rect 4003 29892 4059 29948
rect 4059 29892 4063 29948
rect 3999 29888 4063 29892
rect 4079 29948 4143 29952
rect 4079 29892 4083 29948
rect 4083 29892 4139 29948
rect 4139 29892 4143 29948
rect 4079 29888 4143 29892
rect 4159 29948 4223 29952
rect 4159 29892 4163 29948
rect 4163 29892 4219 29948
rect 4219 29892 4223 29948
rect 4159 29888 4223 29892
rect 9853 29948 9917 29952
rect 9853 29892 9857 29948
rect 9857 29892 9913 29948
rect 9913 29892 9917 29948
rect 9853 29888 9917 29892
rect 9933 29948 9997 29952
rect 9933 29892 9937 29948
rect 9937 29892 9993 29948
rect 9993 29892 9997 29948
rect 9933 29888 9997 29892
rect 10013 29948 10077 29952
rect 10013 29892 10017 29948
rect 10017 29892 10073 29948
rect 10073 29892 10077 29948
rect 10013 29888 10077 29892
rect 10093 29948 10157 29952
rect 10093 29892 10097 29948
rect 10097 29892 10153 29948
rect 10153 29892 10157 29948
rect 10093 29888 10157 29892
rect 15787 29948 15851 29952
rect 15787 29892 15791 29948
rect 15791 29892 15847 29948
rect 15847 29892 15851 29948
rect 15787 29888 15851 29892
rect 15867 29948 15931 29952
rect 15867 29892 15871 29948
rect 15871 29892 15927 29948
rect 15927 29892 15931 29948
rect 15867 29888 15931 29892
rect 15947 29948 16011 29952
rect 15947 29892 15951 29948
rect 15951 29892 16007 29948
rect 16007 29892 16011 29948
rect 15947 29888 16011 29892
rect 16027 29948 16091 29952
rect 16027 29892 16031 29948
rect 16031 29892 16087 29948
rect 16087 29892 16091 29948
rect 16027 29888 16091 29892
rect 21721 29948 21785 29952
rect 21721 29892 21725 29948
rect 21725 29892 21781 29948
rect 21781 29892 21785 29948
rect 21721 29888 21785 29892
rect 21801 29948 21865 29952
rect 21801 29892 21805 29948
rect 21805 29892 21861 29948
rect 21861 29892 21865 29948
rect 21801 29888 21865 29892
rect 21881 29948 21945 29952
rect 21881 29892 21885 29948
rect 21885 29892 21941 29948
rect 21941 29892 21945 29948
rect 21881 29888 21945 29892
rect 21961 29948 22025 29952
rect 21961 29892 21965 29948
rect 21965 29892 22021 29948
rect 22021 29892 22025 29948
rect 21961 29888 22025 29892
rect 2820 29684 2884 29748
rect 5396 29684 5460 29748
rect 13492 29548 13556 29612
rect 6886 29404 6950 29408
rect 6886 29348 6890 29404
rect 6890 29348 6946 29404
rect 6946 29348 6950 29404
rect 6886 29344 6950 29348
rect 6966 29404 7030 29408
rect 6966 29348 6970 29404
rect 6970 29348 7026 29404
rect 7026 29348 7030 29404
rect 6966 29344 7030 29348
rect 7046 29404 7110 29408
rect 7046 29348 7050 29404
rect 7050 29348 7106 29404
rect 7106 29348 7110 29404
rect 7046 29344 7110 29348
rect 7126 29404 7190 29408
rect 7126 29348 7130 29404
rect 7130 29348 7186 29404
rect 7186 29348 7190 29404
rect 7126 29344 7190 29348
rect 12820 29404 12884 29408
rect 12820 29348 12824 29404
rect 12824 29348 12880 29404
rect 12880 29348 12884 29404
rect 12820 29344 12884 29348
rect 12900 29404 12964 29408
rect 12900 29348 12904 29404
rect 12904 29348 12960 29404
rect 12960 29348 12964 29404
rect 12900 29344 12964 29348
rect 12980 29404 13044 29408
rect 12980 29348 12984 29404
rect 12984 29348 13040 29404
rect 13040 29348 13044 29404
rect 12980 29344 13044 29348
rect 13060 29404 13124 29408
rect 13060 29348 13064 29404
rect 13064 29348 13120 29404
rect 13120 29348 13124 29404
rect 13060 29344 13124 29348
rect 18754 29404 18818 29408
rect 18754 29348 18758 29404
rect 18758 29348 18814 29404
rect 18814 29348 18818 29404
rect 18754 29344 18818 29348
rect 18834 29404 18898 29408
rect 18834 29348 18838 29404
rect 18838 29348 18894 29404
rect 18894 29348 18898 29404
rect 18834 29344 18898 29348
rect 18914 29404 18978 29408
rect 18914 29348 18918 29404
rect 18918 29348 18974 29404
rect 18974 29348 18978 29404
rect 18914 29344 18978 29348
rect 18994 29404 19058 29408
rect 18994 29348 18998 29404
rect 18998 29348 19054 29404
rect 19054 29348 19058 29404
rect 18994 29344 19058 29348
rect 24688 29404 24752 29408
rect 24688 29348 24692 29404
rect 24692 29348 24748 29404
rect 24748 29348 24752 29404
rect 24688 29344 24752 29348
rect 24768 29404 24832 29408
rect 24768 29348 24772 29404
rect 24772 29348 24828 29404
rect 24828 29348 24832 29404
rect 24768 29344 24832 29348
rect 24848 29404 24912 29408
rect 24848 29348 24852 29404
rect 24852 29348 24908 29404
rect 24908 29348 24912 29404
rect 24848 29344 24912 29348
rect 24928 29404 24992 29408
rect 24928 29348 24932 29404
rect 24932 29348 24988 29404
rect 24988 29348 24992 29404
rect 24928 29344 24992 29348
rect 2084 29004 2148 29068
rect 10548 29276 10612 29340
rect 16620 29140 16684 29204
rect 5396 29004 5460 29068
rect 16252 29004 16316 29068
rect 3919 28860 3983 28864
rect 3919 28804 3923 28860
rect 3923 28804 3979 28860
rect 3979 28804 3983 28860
rect 3919 28800 3983 28804
rect 3999 28860 4063 28864
rect 3999 28804 4003 28860
rect 4003 28804 4059 28860
rect 4059 28804 4063 28860
rect 3999 28800 4063 28804
rect 4079 28860 4143 28864
rect 4079 28804 4083 28860
rect 4083 28804 4139 28860
rect 4139 28804 4143 28860
rect 4079 28800 4143 28804
rect 4159 28860 4223 28864
rect 4159 28804 4163 28860
rect 4163 28804 4219 28860
rect 4219 28804 4223 28860
rect 4159 28800 4223 28804
rect 9853 28860 9917 28864
rect 9853 28804 9857 28860
rect 9857 28804 9913 28860
rect 9913 28804 9917 28860
rect 9853 28800 9917 28804
rect 9933 28860 9997 28864
rect 9933 28804 9937 28860
rect 9937 28804 9993 28860
rect 9993 28804 9997 28860
rect 9933 28800 9997 28804
rect 10013 28860 10077 28864
rect 10013 28804 10017 28860
rect 10017 28804 10073 28860
rect 10073 28804 10077 28860
rect 10013 28800 10077 28804
rect 10093 28860 10157 28864
rect 10093 28804 10097 28860
rect 10097 28804 10153 28860
rect 10153 28804 10157 28860
rect 10093 28800 10157 28804
rect 15787 28860 15851 28864
rect 15787 28804 15791 28860
rect 15791 28804 15847 28860
rect 15847 28804 15851 28860
rect 15787 28800 15851 28804
rect 15867 28860 15931 28864
rect 15867 28804 15871 28860
rect 15871 28804 15927 28860
rect 15927 28804 15931 28860
rect 15867 28800 15931 28804
rect 15947 28860 16011 28864
rect 15947 28804 15951 28860
rect 15951 28804 16007 28860
rect 16007 28804 16011 28860
rect 15947 28800 16011 28804
rect 16027 28860 16091 28864
rect 16027 28804 16031 28860
rect 16031 28804 16087 28860
rect 16087 28804 16091 28860
rect 16027 28800 16091 28804
rect 21721 28860 21785 28864
rect 21721 28804 21725 28860
rect 21725 28804 21781 28860
rect 21781 28804 21785 28860
rect 21721 28800 21785 28804
rect 21801 28860 21865 28864
rect 21801 28804 21805 28860
rect 21805 28804 21861 28860
rect 21861 28804 21865 28860
rect 21801 28800 21865 28804
rect 21881 28860 21945 28864
rect 21881 28804 21885 28860
rect 21885 28804 21941 28860
rect 21941 28804 21945 28860
rect 21881 28800 21945 28804
rect 21961 28860 22025 28864
rect 21961 28804 21965 28860
rect 21965 28804 22021 28860
rect 22021 28804 22025 28860
rect 21961 28800 22025 28804
rect 10364 28732 10428 28796
rect 16804 28732 16868 28796
rect 1900 28656 1964 28660
rect 1900 28600 1950 28656
rect 1950 28600 1964 28656
rect 1900 28596 1964 28600
rect 17172 28596 17236 28660
rect 2636 28520 2700 28524
rect 2636 28464 2650 28520
rect 2650 28464 2700 28520
rect 2636 28460 2700 28464
rect 5028 28520 5092 28524
rect 5028 28464 5042 28520
rect 5042 28464 5092 28520
rect 5028 28460 5092 28464
rect 1716 28324 1780 28388
rect 13676 28460 13740 28524
rect 6886 28316 6950 28320
rect 6886 28260 6890 28316
rect 6890 28260 6946 28316
rect 6946 28260 6950 28316
rect 6886 28256 6950 28260
rect 6966 28316 7030 28320
rect 6966 28260 6970 28316
rect 6970 28260 7026 28316
rect 7026 28260 7030 28316
rect 6966 28256 7030 28260
rect 7046 28316 7110 28320
rect 7046 28260 7050 28316
rect 7050 28260 7106 28316
rect 7106 28260 7110 28316
rect 7046 28256 7110 28260
rect 7126 28316 7190 28320
rect 7126 28260 7130 28316
rect 7130 28260 7186 28316
rect 7186 28260 7190 28316
rect 7126 28256 7190 28260
rect 12820 28316 12884 28320
rect 12820 28260 12824 28316
rect 12824 28260 12880 28316
rect 12880 28260 12884 28316
rect 12820 28256 12884 28260
rect 12900 28316 12964 28320
rect 12900 28260 12904 28316
rect 12904 28260 12960 28316
rect 12960 28260 12964 28316
rect 12900 28256 12964 28260
rect 12980 28316 13044 28320
rect 12980 28260 12984 28316
rect 12984 28260 13040 28316
rect 13040 28260 13044 28316
rect 12980 28256 13044 28260
rect 13060 28316 13124 28320
rect 13060 28260 13064 28316
rect 13064 28260 13120 28316
rect 13120 28260 13124 28316
rect 13060 28256 13124 28260
rect 18754 28316 18818 28320
rect 18754 28260 18758 28316
rect 18758 28260 18814 28316
rect 18814 28260 18818 28316
rect 18754 28256 18818 28260
rect 18834 28316 18898 28320
rect 18834 28260 18838 28316
rect 18838 28260 18894 28316
rect 18894 28260 18898 28316
rect 18834 28256 18898 28260
rect 18914 28316 18978 28320
rect 18914 28260 18918 28316
rect 18918 28260 18974 28316
rect 18974 28260 18978 28316
rect 18914 28256 18978 28260
rect 18994 28316 19058 28320
rect 18994 28260 18998 28316
rect 18998 28260 19054 28316
rect 19054 28260 19058 28316
rect 18994 28256 19058 28260
rect 24688 28316 24752 28320
rect 24688 28260 24692 28316
rect 24692 28260 24748 28316
rect 24748 28260 24752 28316
rect 24688 28256 24752 28260
rect 24768 28316 24832 28320
rect 24768 28260 24772 28316
rect 24772 28260 24828 28316
rect 24828 28260 24832 28316
rect 24768 28256 24832 28260
rect 24848 28316 24912 28320
rect 24848 28260 24852 28316
rect 24852 28260 24908 28316
rect 24908 28260 24912 28316
rect 24848 28256 24912 28260
rect 24928 28316 24992 28320
rect 24928 28260 24932 28316
rect 24932 28260 24988 28316
rect 24988 28260 24992 28316
rect 24928 28256 24992 28260
rect 612 28188 676 28252
rect 20668 27916 20732 27980
rect 16252 27780 16316 27844
rect 3919 27772 3983 27776
rect 3919 27716 3923 27772
rect 3923 27716 3979 27772
rect 3979 27716 3983 27772
rect 3919 27712 3983 27716
rect 3999 27772 4063 27776
rect 3999 27716 4003 27772
rect 4003 27716 4059 27772
rect 4059 27716 4063 27772
rect 3999 27712 4063 27716
rect 4079 27772 4143 27776
rect 4079 27716 4083 27772
rect 4083 27716 4139 27772
rect 4139 27716 4143 27772
rect 4079 27712 4143 27716
rect 4159 27772 4223 27776
rect 4159 27716 4163 27772
rect 4163 27716 4219 27772
rect 4219 27716 4223 27772
rect 4159 27712 4223 27716
rect 9853 27772 9917 27776
rect 9853 27716 9857 27772
rect 9857 27716 9913 27772
rect 9913 27716 9917 27772
rect 9853 27712 9917 27716
rect 9933 27772 9997 27776
rect 9933 27716 9937 27772
rect 9937 27716 9993 27772
rect 9993 27716 9997 27772
rect 9933 27712 9997 27716
rect 10013 27772 10077 27776
rect 10013 27716 10017 27772
rect 10017 27716 10073 27772
rect 10073 27716 10077 27772
rect 10013 27712 10077 27716
rect 10093 27772 10157 27776
rect 10093 27716 10097 27772
rect 10097 27716 10153 27772
rect 10153 27716 10157 27772
rect 10093 27712 10157 27716
rect 15787 27772 15851 27776
rect 15787 27716 15791 27772
rect 15791 27716 15847 27772
rect 15847 27716 15851 27772
rect 15787 27712 15851 27716
rect 15867 27772 15931 27776
rect 15867 27716 15871 27772
rect 15871 27716 15927 27772
rect 15927 27716 15931 27772
rect 15867 27712 15931 27716
rect 15947 27772 16011 27776
rect 15947 27716 15951 27772
rect 15951 27716 16007 27772
rect 16007 27716 16011 27772
rect 15947 27712 16011 27716
rect 16027 27772 16091 27776
rect 16027 27716 16031 27772
rect 16031 27716 16087 27772
rect 16087 27716 16091 27772
rect 16027 27712 16091 27716
rect 21721 27772 21785 27776
rect 21721 27716 21725 27772
rect 21725 27716 21781 27772
rect 21781 27716 21785 27772
rect 21721 27712 21785 27716
rect 21801 27772 21865 27776
rect 21801 27716 21805 27772
rect 21805 27716 21861 27772
rect 21861 27716 21865 27772
rect 21801 27712 21865 27716
rect 21881 27772 21945 27776
rect 21881 27716 21885 27772
rect 21885 27716 21941 27772
rect 21941 27716 21945 27772
rect 21881 27712 21945 27716
rect 21961 27772 22025 27776
rect 21961 27716 21965 27772
rect 21965 27716 22021 27772
rect 22021 27716 22025 27772
rect 21961 27712 22025 27716
rect 17540 27644 17604 27708
rect 20852 27644 20916 27708
rect 3004 27432 3068 27436
rect 3004 27376 3018 27432
rect 3018 27376 3068 27432
rect 3004 27372 3068 27376
rect 5948 27372 6012 27436
rect 6886 27228 6950 27232
rect 6886 27172 6890 27228
rect 6890 27172 6946 27228
rect 6946 27172 6950 27228
rect 6886 27168 6950 27172
rect 6966 27228 7030 27232
rect 6966 27172 6970 27228
rect 6970 27172 7026 27228
rect 7026 27172 7030 27228
rect 6966 27168 7030 27172
rect 7046 27228 7110 27232
rect 7046 27172 7050 27228
rect 7050 27172 7106 27228
rect 7106 27172 7110 27228
rect 7046 27168 7110 27172
rect 7126 27228 7190 27232
rect 7126 27172 7130 27228
rect 7130 27172 7186 27228
rect 7186 27172 7190 27228
rect 7126 27168 7190 27172
rect 12820 27228 12884 27232
rect 12820 27172 12824 27228
rect 12824 27172 12880 27228
rect 12880 27172 12884 27228
rect 12820 27168 12884 27172
rect 12900 27228 12964 27232
rect 12900 27172 12904 27228
rect 12904 27172 12960 27228
rect 12960 27172 12964 27228
rect 12900 27168 12964 27172
rect 12980 27228 13044 27232
rect 12980 27172 12984 27228
rect 12984 27172 13040 27228
rect 13040 27172 13044 27228
rect 12980 27168 13044 27172
rect 13060 27228 13124 27232
rect 13060 27172 13064 27228
rect 13064 27172 13120 27228
rect 13120 27172 13124 27228
rect 13060 27168 13124 27172
rect 18754 27228 18818 27232
rect 18754 27172 18758 27228
rect 18758 27172 18814 27228
rect 18814 27172 18818 27228
rect 18754 27168 18818 27172
rect 18834 27228 18898 27232
rect 18834 27172 18838 27228
rect 18838 27172 18894 27228
rect 18894 27172 18898 27228
rect 18834 27168 18898 27172
rect 18914 27228 18978 27232
rect 18914 27172 18918 27228
rect 18918 27172 18974 27228
rect 18974 27172 18978 27228
rect 18914 27168 18978 27172
rect 18994 27228 19058 27232
rect 18994 27172 18998 27228
rect 18998 27172 19054 27228
rect 19054 27172 19058 27228
rect 18994 27168 19058 27172
rect 24688 27228 24752 27232
rect 24688 27172 24692 27228
rect 24692 27172 24748 27228
rect 24748 27172 24752 27228
rect 24688 27168 24752 27172
rect 24768 27228 24832 27232
rect 24768 27172 24772 27228
rect 24772 27172 24828 27228
rect 24828 27172 24832 27228
rect 24768 27168 24832 27172
rect 24848 27228 24912 27232
rect 24848 27172 24852 27228
rect 24852 27172 24908 27228
rect 24908 27172 24912 27228
rect 24848 27168 24912 27172
rect 24928 27228 24992 27232
rect 24928 27172 24932 27228
rect 24932 27172 24988 27228
rect 24988 27172 24992 27228
rect 24928 27168 24992 27172
rect 1348 26828 1412 26892
rect 2084 26828 2148 26892
rect 20852 26888 20916 26892
rect 20852 26832 20866 26888
rect 20866 26832 20916 26888
rect 20852 26828 20916 26832
rect 2452 26692 2516 26756
rect 11284 26692 11348 26756
rect 3919 26684 3983 26688
rect 3919 26628 3923 26684
rect 3923 26628 3979 26684
rect 3979 26628 3983 26684
rect 3919 26624 3983 26628
rect 3999 26684 4063 26688
rect 3999 26628 4003 26684
rect 4003 26628 4059 26684
rect 4059 26628 4063 26684
rect 3999 26624 4063 26628
rect 4079 26684 4143 26688
rect 4079 26628 4083 26684
rect 4083 26628 4139 26684
rect 4139 26628 4143 26684
rect 4079 26624 4143 26628
rect 4159 26684 4223 26688
rect 4159 26628 4163 26684
rect 4163 26628 4219 26684
rect 4219 26628 4223 26684
rect 4159 26624 4223 26628
rect 9853 26684 9917 26688
rect 9853 26628 9857 26684
rect 9857 26628 9913 26684
rect 9913 26628 9917 26684
rect 9853 26624 9917 26628
rect 9933 26684 9997 26688
rect 9933 26628 9937 26684
rect 9937 26628 9993 26684
rect 9993 26628 9997 26684
rect 9933 26624 9997 26628
rect 10013 26684 10077 26688
rect 10013 26628 10017 26684
rect 10017 26628 10073 26684
rect 10073 26628 10077 26684
rect 10013 26624 10077 26628
rect 10093 26684 10157 26688
rect 10093 26628 10097 26684
rect 10097 26628 10153 26684
rect 10153 26628 10157 26684
rect 10093 26624 10157 26628
rect 15787 26684 15851 26688
rect 15787 26628 15791 26684
rect 15791 26628 15847 26684
rect 15847 26628 15851 26684
rect 15787 26624 15851 26628
rect 15867 26684 15931 26688
rect 15867 26628 15871 26684
rect 15871 26628 15927 26684
rect 15927 26628 15931 26684
rect 15867 26624 15931 26628
rect 15947 26684 16011 26688
rect 15947 26628 15951 26684
rect 15951 26628 16007 26684
rect 16007 26628 16011 26684
rect 15947 26624 16011 26628
rect 16027 26684 16091 26688
rect 16027 26628 16031 26684
rect 16031 26628 16087 26684
rect 16087 26628 16091 26684
rect 16027 26624 16091 26628
rect 21721 26684 21785 26688
rect 21721 26628 21725 26684
rect 21725 26628 21781 26684
rect 21781 26628 21785 26684
rect 21721 26624 21785 26628
rect 21801 26684 21865 26688
rect 21801 26628 21805 26684
rect 21805 26628 21861 26684
rect 21861 26628 21865 26684
rect 21801 26624 21865 26628
rect 21881 26684 21945 26688
rect 21881 26628 21885 26684
rect 21885 26628 21941 26684
rect 21941 26628 21945 26684
rect 21881 26624 21945 26628
rect 21961 26684 22025 26688
rect 21961 26628 21965 26684
rect 21965 26628 22021 26684
rect 22021 26628 22025 26684
rect 21961 26624 22025 26628
rect 9260 26420 9324 26484
rect 6132 26148 6196 26212
rect 6886 26140 6950 26144
rect 6886 26084 6890 26140
rect 6890 26084 6946 26140
rect 6946 26084 6950 26140
rect 6886 26080 6950 26084
rect 6966 26140 7030 26144
rect 6966 26084 6970 26140
rect 6970 26084 7026 26140
rect 7026 26084 7030 26140
rect 6966 26080 7030 26084
rect 7046 26140 7110 26144
rect 7046 26084 7050 26140
rect 7050 26084 7106 26140
rect 7106 26084 7110 26140
rect 7046 26080 7110 26084
rect 7126 26140 7190 26144
rect 7126 26084 7130 26140
rect 7130 26084 7186 26140
rect 7186 26084 7190 26140
rect 7126 26080 7190 26084
rect 12820 26140 12884 26144
rect 12820 26084 12824 26140
rect 12824 26084 12880 26140
rect 12880 26084 12884 26140
rect 12820 26080 12884 26084
rect 12900 26140 12964 26144
rect 12900 26084 12904 26140
rect 12904 26084 12960 26140
rect 12960 26084 12964 26140
rect 12900 26080 12964 26084
rect 12980 26140 13044 26144
rect 12980 26084 12984 26140
rect 12984 26084 13040 26140
rect 13040 26084 13044 26140
rect 12980 26080 13044 26084
rect 13060 26140 13124 26144
rect 13060 26084 13064 26140
rect 13064 26084 13120 26140
rect 13120 26084 13124 26140
rect 13060 26080 13124 26084
rect 18754 26140 18818 26144
rect 18754 26084 18758 26140
rect 18758 26084 18814 26140
rect 18814 26084 18818 26140
rect 18754 26080 18818 26084
rect 18834 26140 18898 26144
rect 18834 26084 18838 26140
rect 18838 26084 18894 26140
rect 18894 26084 18898 26140
rect 18834 26080 18898 26084
rect 18914 26140 18978 26144
rect 18914 26084 18918 26140
rect 18918 26084 18974 26140
rect 18974 26084 18978 26140
rect 18914 26080 18978 26084
rect 18994 26140 19058 26144
rect 18994 26084 18998 26140
rect 18998 26084 19054 26140
rect 19054 26084 19058 26140
rect 18994 26080 19058 26084
rect 24688 26140 24752 26144
rect 24688 26084 24692 26140
rect 24692 26084 24748 26140
rect 24748 26084 24752 26140
rect 24688 26080 24752 26084
rect 24768 26140 24832 26144
rect 24768 26084 24772 26140
rect 24772 26084 24828 26140
rect 24828 26084 24832 26140
rect 24768 26080 24832 26084
rect 24848 26140 24912 26144
rect 24848 26084 24852 26140
rect 24852 26084 24908 26140
rect 24908 26084 24912 26140
rect 24848 26080 24912 26084
rect 24928 26140 24992 26144
rect 24928 26084 24932 26140
rect 24932 26084 24988 26140
rect 24988 26084 24992 26140
rect 24928 26080 24992 26084
rect 2268 26012 2332 26076
rect 2452 26012 2516 26076
rect 4660 25876 4724 25940
rect 6500 25876 6564 25940
rect 6132 25604 6196 25668
rect 3919 25596 3983 25600
rect 3919 25540 3923 25596
rect 3923 25540 3979 25596
rect 3979 25540 3983 25596
rect 3919 25536 3983 25540
rect 3999 25596 4063 25600
rect 3999 25540 4003 25596
rect 4003 25540 4059 25596
rect 4059 25540 4063 25596
rect 3999 25536 4063 25540
rect 4079 25596 4143 25600
rect 4079 25540 4083 25596
rect 4083 25540 4139 25596
rect 4139 25540 4143 25596
rect 4079 25536 4143 25540
rect 4159 25596 4223 25600
rect 4159 25540 4163 25596
rect 4163 25540 4219 25596
rect 4219 25540 4223 25596
rect 4159 25536 4223 25540
rect 10732 25740 10796 25804
rect 9853 25596 9917 25600
rect 9853 25540 9857 25596
rect 9857 25540 9913 25596
rect 9913 25540 9917 25596
rect 9853 25536 9917 25540
rect 9933 25596 9997 25600
rect 9933 25540 9937 25596
rect 9937 25540 9993 25596
rect 9993 25540 9997 25596
rect 9933 25536 9997 25540
rect 10013 25596 10077 25600
rect 10013 25540 10017 25596
rect 10017 25540 10073 25596
rect 10073 25540 10077 25596
rect 10013 25536 10077 25540
rect 10093 25596 10157 25600
rect 10093 25540 10097 25596
rect 10097 25540 10153 25596
rect 10153 25540 10157 25596
rect 10093 25536 10157 25540
rect 15787 25596 15851 25600
rect 15787 25540 15791 25596
rect 15791 25540 15847 25596
rect 15847 25540 15851 25596
rect 15787 25536 15851 25540
rect 15867 25596 15931 25600
rect 15867 25540 15871 25596
rect 15871 25540 15927 25596
rect 15927 25540 15931 25596
rect 15867 25536 15931 25540
rect 15947 25596 16011 25600
rect 15947 25540 15951 25596
rect 15951 25540 16007 25596
rect 16007 25540 16011 25596
rect 15947 25536 16011 25540
rect 16027 25596 16091 25600
rect 16027 25540 16031 25596
rect 16031 25540 16087 25596
rect 16087 25540 16091 25596
rect 16027 25536 16091 25540
rect 21721 25596 21785 25600
rect 21721 25540 21725 25596
rect 21725 25540 21781 25596
rect 21781 25540 21785 25596
rect 21721 25536 21785 25540
rect 21801 25596 21865 25600
rect 21801 25540 21805 25596
rect 21805 25540 21861 25596
rect 21861 25540 21865 25596
rect 21801 25536 21865 25540
rect 21881 25596 21945 25600
rect 21881 25540 21885 25596
rect 21885 25540 21941 25596
rect 21941 25540 21945 25596
rect 21881 25536 21945 25540
rect 21961 25596 22025 25600
rect 21961 25540 21965 25596
rect 21965 25540 22021 25596
rect 22021 25540 22025 25596
rect 21961 25536 22025 25540
rect 10364 25392 10428 25396
rect 10364 25336 10378 25392
rect 10378 25336 10428 25392
rect 10364 25332 10428 25336
rect 16620 25196 16684 25260
rect 21588 25196 21652 25260
rect 6886 25052 6950 25056
rect 6886 24996 6890 25052
rect 6890 24996 6946 25052
rect 6946 24996 6950 25052
rect 6886 24992 6950 24996
rect 6966 25052 7030 25056
rect 6966 24996 6970 25052
rect 6970 24996 7026 25052
rect 7026 24996 7030 25052
rect 6966 24992 7030 24996
rect 7046 25052 7110 25056
rect 7046 24996 7050 25052
rect 7050 24996 7106 25052
rect 7106 24996 7110 25052
rect 7046 24992 7110 24996
rect 7126 25052 7190 25056
rect 7126 24996 7130 25052
rect 7130 24996 7186 25052
rect 7186 24996 7190 25052
rect 7126 24992 7190 24996
rect 12820 25052 12884 25056
rect 12820 24996 12824 25052
rect 12824 24996 12880 25052
rect 12880 24996 12884 25052
rect 12820 24992 12884 24996
rect 12900 25052 12964 25056
rect 12900 24996 12904 25052
rect 12904 24996 12960 25052
rect 12960 24996 12964 25052
rect 12900 24992 12964 24996
rect 12980 25052 13044 25056
rect 12980 24996 12984 25052
rect 12984 24996 13040 25052
rect 13040 24996 13044 25052
rect 12980 24992 13044 24996
rect 13060 25052 13124 25056
rect 13060 24996 13064 25052
rect 13064 24996 13120 25052
rect 13120 24996 13124 25052
rect 13060 24992 13124 24996
rect 18754 25052 18818 25056
rect 18754 24996 18758 25052
rect 18758 24996 18814 25052
rect 18814 24996 18818 25052
rect 18754 24992 18818 24996
rect 18834 25052 18898 25056
rect 18834 24996 18838 25052
rect 18838 24996 18894 25052
rect 18894 24996 18898 25052
rect 18834 24992 18898 24996
rect 18914 25052 18978 25056
rect 18914 24996 18918 25052
rect 18918 24996 18974 25052
rect 18974 24996 18978 25052
rect 18914 24992 18978 24996
rect 18994 25052 19058 25056
rect 18994 24996 18998 25052
rect 18998 24996 19054 25052
rect 19054 24996 19058 25052
rect 18994 24992 19058 24996
rect 24688 25052 24752 25056
rect 24688 24996 24692 25052
rect 24692 24996 24748 25052
rect 24748 24996 24752 25052
rect 24688 24992 24752 24996
rect 24768 25052 24832 25056
rect 24768 24996 24772 25052
rect 24772 24996 24828 25052
rect 24828 24996 24832 25052
rect 24768 24992 24832 24996
rect 24848 25052 24912 25056
rect 24848 24996 24852 25052
rect 24852 24996 24908 25052
rect 24908 24996 24912 25052
rect 24848 24992 24912 24996
rect 24928 25052 24992 25056
rect 24928 24996 24932 25052
rect 24932 24996 24988 25052
rect 24988 24996 24992 25052
rect 24928 24992 24992 24996
rect 5580 24788 5644 24852
rect 3919 24508 3983 24512
rect 3919 24452 3923 24508
rect 3923 24452 3979 24508
rect 3979 24452 3983 24508
rect 3919 24448 3983 24452
rect 3999 24508 4063 24512
rect 3999 24452 4003 24508
rect 4003 24452 4059 24508
rect 4059 24452 4063 24508
rect 3999 24448 4063 24452
rect 4079 24508 4143 24512
rect 4079 24452 4083 24508
rect 4083 24452 4139 24508
rect 4139 24452 4143 24508
rect 4079 24448 4143 24452
rect 4159 24508 4223 24512
rect 4159 24452 4163 24508
rect 4163 24452 4219 24508
rect 4219 24452 4223 24508
rect 4159 24448 4223 24452
rect 12204 24652 12268 24716
rect 9853 24508 9917 24512
rect 9853 24452 9857 24508
rect 9857 24452 9913 24508
rect 9913 24452 9917 24508
rect 9853 24448 9917 24452
rect 9933 24508 9997 24512
rect 9933 24452 9937 24508
rect 9937 24452 9993 24508
rect 9993 24452 9997 24508
rect 9933 24448 9997 24452
rect 10013 24508 10077 24512
rect 10013 24452 10017 24508
rect 10017 24452 10073 24508
rect 10073 24452 10077 24508
rect 10013 24448 10077 24452
rect 10093 24508 10157 24512
rect 10093 24452 10097 24508
rect 10097 24452 10153 24508
rect 10153 24452 10157 24508
rect 10093 24448 10157 24452
rect 15787 24508 15851 24512
rect 15787 24452 15791 24508
rect 15791 24452 15847 24508
rect 15847 24452 15851 24508
rect 15787 24448 15851 24452
rect 15867 24508 15931 24512
rect 15867 24452 15871 24508
rect 15871 24452 15927 24508
rect 15927 24452 15931 24508
rect 15867 24448 15931 24452
rect 15947 24508 16011 24512
rect 15947 24452 15951 24508
rect 15951 24452 16007 24508
rect 16007 24452 16011 24508
rect 15947 24448 16011 24452
rect 16027 24508 16091 24512
rect 16027 24452 16031 24508
rect 16031 24452 16087 24508
rect 16087 24452 16091 24508
rect 16027 24448 16091 24452
rect 21721 24508 21785 24512
rect 21721 24452 21725 24508
rect 21725 24452 21781 24508
rect 21781 24452 21785 24508
rect 21721 24448 21785 24452
rect 21801 24508 21865 24512
rect 21801 24452 21805 24508
rect 21805 24452 21861 24508
rect 21861 24452 21865 24508
rect 21801 24448 21865 24452
rect 21881 24508 21945 24512
rect 21881 24452 21885 24508
rect 21885 24452 21941 24508
rect 21941 24452 21945 24508
rect 21881 24448 21945 24452
rect 21961 24508 22025 24512
rect 21961 24452 21965 24508
rect 21965 24452 22021 24508
rect 22021 24452 22025 24508
rect 21961 24448 22025 24452
rect 3004 24244 3068 24308
rect 10916 24304 10980 24308
rect 10916 24248 10930 24304
rect 10930 24248 10980 24304
rect 10916 24244 10980 24248
rect 6886 23964 6950 23968
rect 6886 23908 6890 23964
rect 6890 23908 6946 23964
rect 6946 23908 6950 23964
rect 6886 23904 6950 23908
rect 6966 23964 7030 23968
rect 6966 23908 6970 23964
rect 6970 23908 7026 23964
rect 7026 23908 7030 23964
rect 6966 23904 7030 23908
rect 7046 23964 7110 23968
rect 7046 23908 7050 23964
rect 7050 23908 7106 23964
rect 7106 23908 7110 23964
rect 7046 23904 7110 23908
rect 7126 23964 7190 23968
rect 7126 23908 7130 23964
rect 7130 23908 7186 23964
rect 7186 23908 7190 23964
rect 7126 23904 7190 23908
rect 12820 23964 12884 23968
rect 12820 23908 12824 23964
rect 12824 23908 12880 23964
rect 12880 23908 12884 23964
rect 12820 23904 12884 23908
rect 12900 23964 12964 23968
rect 12900 23908 12904 23964
rect 12904 23908 12960 23964
rect 12960 23908 12964 23964
rect 12900 23904 12964 23908
rect 12980 23964 13044 23968
rect 12980 23908 12984 23964
rect 12984 23908 13040 23964
rect 13040 23908 13044 23964
rect 12980 23904 13044 23908
rect 13060 23964 13124 23968
rect 13060 23908 13064 23964
rect 13064 23908 13120 23964
rect 13120 23908 13124 23964
rect 13060 23904 13124 23908
rect 18754 23964 18818 23968
rect 18754 23908 18758 23964
rect 18758 23908 18814 23964
rect 18814 23908 18818 23964
rect 18754 23904 18818 23908
rect 18834 23964 18898 23968
rect 18834 23908 18838 23964
rect 18838 23908 18894 23964
rect 18894 23908 18898 23964
rect 18834 23904 18898 23908
rect 18914 23964 18978 23968
rect 18914 23908 18918 23964
rect 18918 23908 18974 23964
rect 18974 23908 18978 23964
rect 18914 23904 18978 23908
rect 18994 23964 19058 23968
rect 18994 23908 18998 23964
rect 18998 23908 19054 23964
rect 19054 23908 19058 23964
rect 18994 23904 19058 23908
rect 24688 23964 24752 23968
rect 24688 23908 24692 23964
rect 24692 23908 24748 23964
rect 24748 23908 24752 23964
rect 24688 23904 24752 23908
rect 24768 23964 24832 23968
rect 24768 23908 24772 23964
rect 24772 23908 24828 23964
rect 24828 23908 24832 23964
rect 24768 23904 24832 23908
rect 24848 23964 24912 23968
rect 24848 23908 24852 23964
rect 24852 23908 24908 23964
rect 24908 23908 24912 23964
rect 24848 23904 24912 23908
rect 24928 23964 24992 23968
rect 24928 23908 24932 23964
rect 24932 23908 24988 23964
rect 24988 23908 24992 23964
rect 24928 23904 24992 23908
rect 2820 23896 2884 23900
rect 2820 23840 2834 23896
rect 2834 23840 2884 23896
rect 2820 23836 2884 23840
rect 21404 23564 21468 23628
rect 1716 23428 1780 23492
rect 4844 23428 4908 23492
rect 3919 23420 3983 23424
rect 3919 23364 3923 23420
rect 3923 23364 3979 23420
rect 3979 23364 3983 23420
rect 3919 23360 3983 23364
rect 3999 23420 4063 23424
rect 3999 23364 4003 23420
rect 4003 23364 4059 23420
rect 4059 23364 4063 23420
rect 3999 23360 4063 23364
rect 4079 23420 4143 23424
rect 4079 23364 4083 23420
rect 4083 23364 4139 23420
rect 4139 23364 4143 23420
rect 4079 23360 4143 23364
rect 4159 23420 4223 23424
rect 4159 23364 4163 23420
rect 4163 23364 4219 23420
rect 4219 23364 4223 23420
rect 4159 23360 4223 23364
rect 5948 23428 6012 23492
rect 6500 23428 6564 23492
rect 13492 23428 13556 23492
rect 9853 23420 9917 23424
rect 9853 23364 9857 23420
rect 9857 23364 9913 23420
rect 9913 23364 9917 23420
rect 9853 23360 9917 23364
rect 9933 23420 9997 23424
rect 9933 23364 9937 23420
rect 9937 23364 9993 23420
rect 9993 23364 9997 23420
rect 9933 23360 9997 23364
rect 10013 23420 10077 23424
rect 10013 23364 10017 23420
rect 10017 23364 10073 23420
rect 10073 23364 10077 23420
rect 10013 23360 10077 23364
rect 10093 23420 10157 23424
rect 10093 23364 10097 23420
rect 10097 23364 10153 23420
rect 10153 23364 10157 23420
rect 10093 23360 10157 23364
rect 15787 23420 15851 23424
rect 15787 23364 15791 23420
rect 15791 23364 15847 23420
rect 15847 23364 15851 23420
rect 15787 23360 15851 23364
rect 15867 23420 15931 23424
rect 15867 23364 15871 23420
rect 15871 23364 15927 23420
rect 15927 23364 15931 23420
rect 15867 23360 15931 23364
rect 15947 23420 16011 23424
rect 15947 23364 15951 23420
rect 15951 23364 16007 23420
rect 16007 23364 16011 23420
rect 15947 23360 16011 23364
rect 16027 23420 16091 23424
rect 16027 23364 16031 23420
rect 16031 23364 16087 23420
rect 16087 23364 16091 23420
rect 16027 23360 16091 23364
rect 21721 23420 21785 23424
rect 21721 23364 21725 23420
rect 21725 23364 21781 23420
rect 21781 23364 21785 23420
rect 21721 23360 21785 23364
rect 21801 23420 21865 23424
rect 21801 23364 21805 23420
rect 21805 23364 21861 23420
rect 21861 23364 21865 23420
rect 21801 23360 21865 23364
rect 21881 23420 21945 23424
rect 21881 23364 21885 23420
rect 21885 23364 21941 23420
rect 21941 23364 21945 23420
rect 21881 23360 21945 23364
rect 21961 23420 22025 23424
rect 21961 23364 21965 23420
rect 21965 23364 22021 23420
rect 22021 23364 22025 23420
rect 21961 23360 22025 23364
rect 13676 23352 13740 23356
rect 13676 23296 13726 23352
rect 13726 23296 13740 23352
rect 13676 23292 13740 23296
rect 11652 23156 11716 23220
rect 2268 22612 2332 22676
rect 17540 23020 17604 23084
rect 12020 22884 12084 22948
rect 13676 22884 13740 22948
rect 6886 22876 6950 22880
rect 6886 22820 6890 22876
rect 6890 22820 6946 22876
rect 6946 22820 6950 22876
rect 6886 22816 6950 22820
rect 6966 22876 7030 22880
rect 6966 22820 6970 22876
rect 6970 22820 7026 22876
rect 7026 22820 7030 22876
rect 6966 22816 7030 22820
rect 7046 22876 7110 22880
rect 7046 22820 7050 22876
rect 7050 22820 7106 22876
rect 7106 22820 7110 22876
rect 7046 22816 7110 22820
rect 7126 22876 7190 22880
rect 7126 22820 7130 22876
rect 7130 22820 7186 22876
rect 7186 22820 7190 22876
rect 7126 22816 7190 22820
rect 12820 22876 12884 22880
rect 12820 22820 12824 22876
rect 12824 22820 12880 22876
rect 12880 22820 12884 22876
rect 12820 22816 12884 22820
rect 12900 22876 12964 22880
rect 12900 22820 12904 22876
rect 12904 22820 12960 22876
rect 12960 22820 12964 22876
rect 12900 22816 12964 22820
rect 12980 22876 13044 22880
rect 12980 22820 12984 22876
rect 12984 22820 13040 22876
rect 13040 22820 13044 22876
rect 12980 22816 13044 22820
rect 13060 22876 13124 22880
rect 13060 22820 13064 22876
rect 13064 22820 13120 22876
rect 13120 22820 13124 22876
rect 13060 22816 13124 22820
rect 18754 22876 18818 22880
rect 18754 22820 18758 22876
rect 18758 22820 18814 22876
rect 18814 22820 18818 22876
rect 18754 22816 18818 22820
rect 18834 22876 18898 22880
rect 18834 22820 18838 22876
rect 18838 22820 18894 22876
rect 18894 22820 18898 22876
rect 18834 22816 18898 22820
rect 18914 22876 18978 22880
rect 18914 22820 18918 22876
rect 18918 22820 18974 22876
rect 18974 22820 18978 22876
rect 18914 22816 18978 22820
rect 18994 22876 19058 22880
rect 18994 22820 18998 22876
rect 18998 22820 19054 22876
rect 19054 22820 19058 22876
rect 18994 22816 19058 22820
rect 24688 22876 24752 22880
rect 24688 22820 24692 22876
rect 24692 22820 24748 22876
rect 24748 22820 24752 22876
rect 24688 22816 24752 22820
rect 24768 22876 24832 22880
rect 24768 22820 24772 22876
rect 24772 22820 24828 22876
rect 24828 22820 24832 22876
rect 24768 22816 24832 22820
rect 24848 22876 24912 22880
rect 24848 22820 24852 22876
rect 24852 22820 24908 22876
rect 24908 22820 24912 22876
rect 24848 22816 24912 22820
rect 24928 22876 24992 22880
rect 24928 22820 24932 22876
rect 24932 22820 24988 22876
rect 24988 22820 24992 22876
rect 24928 22816 24992 22820
rect 4660 22808 4724 22812
rect 4660 22752 4674 22808
rect 4674 22752 4724 22808
rect 4660 22748 4724 22752
rect 1900 21932 1964 21996
rect 11100 22476 11164 22540
rect 11468 22476 11532 22540
rect 3919 22332 3983 22336
rect 3919 22276 3923 22332
rect 3923 22276 3979 22332
rect 3979 22276 3983 22332
rect 3919 22272 3983 22276
rect 3999 22332 4063 22336
rect 3999 22276 4003 22332
rect 4003 22276 4059 22332
rect 4059 22276 4063 22332
rect 3999 22272 4063 22276
rect 4079 22332 4143 22336
rect 4079 22276 4083 22332
rect 4083 22276 4139 22332
rect 4139 22276 4143 22332
rect 4079 22272 4143 22276
rect 4159 22332 4223 22336
rect 4159 22276 4163 22332
rect 4163 22276 4219 22332
rect 4219 22276 4223 22332
rect 4159 22272 4223 22276
rect 9853 22332 9917 22336
rect 9853 22276 9857 22332
rect 9857 22276 9913 22332
rect 9913 22276 9917 22332
rect 9853 22272 9917 22276
rect 9933 22332 9997 22336
rect 9933 22276 9937 22332
rect 9937 22276 9993 22332
rect 9993 22276 9997 22332
rect 9933 22272 9997 22276
rect 10013 22332 10077 22336
rect 10013 22276 10017 22332
rect 10017 22276 10073 22332
rect 10073 22276 10077 22332
rect 10013 22272 10077 22276
rect 10093 22332 10157 22336
rect 10093 22276 10097 22332
rect 10097 22276 10153 22332
rect 10153 22276 10157 22332
rect 10093 22272 10157 22276
rect 15787 22332 15851 22336
rect 15787 22276 15791 22332
rect 15791 22276 15847 22332
rect 15847 22276 15851 22332
rect 15787 22272 15851 22276
rect 15867 22332 15931 22336
rect 15867 22276 15871 22332
rect 15871 22276 15927 22332
rect 15927 22276 15931 22332
rect 15867 22272 15931 22276
rect 15947 22332 16011 22336
rect 15947 22276 15951 22332
rect 15951 22276 16007 22332
rect 16007 22276 16011 22332
rect 15947 22272 16011 22276
rect 16027 22332 16091 22336
rect 16027 22276 16031 22332
rect 16031 22276 16087 22332
rect 16087 22276 16091 22332
rect 16027 22272 16091 22276
rect 21721 22332 21785 22336
rect 21721 22276 21725 22332
rect 21725 22276 21781 22332
rect 21781 22276 21785 22332
rect 21721 22272 21785 22276
rect 21801 22332 21865 22336
rect 21801 22276 21805 22332
rect 21805 22276 21861 22332
rect 21861 22276 21865 22332
rect 21801 22272 21865 22276
rect 21881 22332 21945 22336
rect 21881 22276 21885 22332
rect 21885 22276 21941 22332
rect 21941 22276 21945 22332
rect 21881 22272 21945 22276
rect 21961 22332 22025 22336
rect 21961 22276 21965 22332
rect 21965 22276 22021 22332
rect 22021 22276 22025 22332
rect 21961 22272 22025 22276
rect 5396 21932 5460 21996
rect 6132 21856 6196 21860
rect 6132 21800 6182 21856
rect 6182 21800 6196 21856
rect 6132 21796 6196 21800
rect 9260 21796 9324 21860
rect 6886 21788 6950 21792
rect 6886 21732 6890 21788
rect 6890 21732 6946 21788
rect 6946 21732 6950 21788
rect 6886 21728 6950 21732
rect 6966 21788 7030 21792
rect 6966 21732 6970 21788
rect 6970 21732 7026 21788
rect 7026 21732 7030 21788
rect 6966 21728 7030 21732
rect 7046 21788 7110 21792
rect 7046 21732 7050 21788
rect 7050 21732 7106 21788
rect 7106 21732 7110 21788
rect 7046 21728 7110 21732
rect 7126 21788 7190 21792
rect 7126 21732 7130 21788
rect 7130 21732 7186 21788
rect 7186 21732 7190 21788
rect 7126 21728 7190 21732
rect 12820 21788 12884 21792
rect 12820 21732 12824 21788
rect 12824 21732 12880 21788
rect 12880 21732 12884 21788
rect 12820 21728 12884 21732
rect 12900 21788 12964 21792
rect 12900 21732 12904 21788
rect 12904 21732 12960 21788
rect 12960 21732 12964 21788
rect 12900 21728 12964 21732
rect 12980 21788 13044 21792
rect 12980 21732 12984 21788
rect 12984 21732 13040 21788
rect 13040 21732 13044 21788
rect 12980 21728 13044 21732
rect 13060 21788 13124 21792
rect 13060 21732 13064 21788
rect 13064 21732 13120 21788
rect 13120 21732 13124 21788
rect 13060 21728 13124 21732
rect 18754 21788 18818 21792
rect 18754 21732 18758 21788
rect 18758 21732 18814 21788
rect 18814 21732 18818 21788
rect 18754 21728 18818 21732
rect 18834 21788 18898 21792
rect 18834 21732 18838 21788
rect 18838 21732 18894 21788
rect 18894 21732 18898 21788
rect 18834 21728 18898 21732
rect 18914 21788 18978 21792
rect 18914 21732 18918 21788
rect 18918 21732 18974 21788
rect 18974 21732 18978 21788
rect 18914 21728 18978 21732
rect 18994 21788 19058 21792
rect 18994 21732 18998 21788
rect 18998 21732 19054 21788
rect 19054 21732 19058 21788
rect 18994 21728 19058 21732
rect 24688 21788 24752 21792
rect 24688 21732 24692 21788
rect 24692 21732 24748 21788
rect 24748 21732 24752 21788
rect 24688 21728 24752 21732
rect 24768 21788 24832 21792
rect 24768 21732 24772 21788
rect 24772 21732 24828 21788
rect 24828 21732 24832 21788
rect 24768 21728 24832 21732
rect 24848 21788 24912 21792
rect 24848 21732 24852 21788
rect 24852 21732 24908 21788
rect 24908 21732 24912 21788
rect 24848 21728 24912 21732
rect 24928 21788 24992 21792
rect 24928 21732 24932 21788
rect 24932 21732 24988 21788
rect 24988 21732 24992 21788
rect 24928 21728 24992 21732
rect 16804 21720 16868 21724
rect 16804 21664 16818 21720
rect 16818 21664 16868 21720
rect 16804 21660 16868 21664
rect 3919 21244 3983 21248
rect 3919 21188 3923 21244
rect 3923 21188 3979 21244
rect 3979 21188 3983 21244
rect 3919 21184 3983 21188
rect 3999 21244 4063 21248
rect 3999 21188 4003 21244
rect 4003 21188 4059 21244
rect 4059 21188 4063 21244
rect 3999 21184 4063 21188
rect 4079 21244 4143 21248
rect 4079 21188 4083 21244
rect 4083 21188 4139 21244
rect 4139 21188 4143 21244
rect 4079 21184 4143 21188
rect 4159 21244 4223 21248
rect 4159 21188 4163 21244
rect 4163 21188 4219 21244
rect 4219 21188 4223 21244
rect 4159 21184 4223 21188
rect 9853 21244 9917 21248
rect 9853 21188 9857 21244
rect 9857 21188 9913 21244
rect 9913 21188 9917 21244
rect 9853 21184 9917 21188
rect 9933 21244 9997 21248
rect 9933 21188 9937 21244
rect 9937 21188 9993 21244
rect 9993 21188 9997 21244
rect 9933 21184 9997 21188
rect 10013 21244 10077 21248
rect 10013 21188 10017 21244
rect 10017 21188 10073 21244
rect 10073 21188 10077 21244
rect 10013 21184 10077 21188
rect 10093 21244 10157 21248
rect 10093 21188 10097 21244
rect 10097 21188 10153 21244
rect 10153 21188 10157 21244
rect 10093 21184 10157 21188
rect 15787 21244 15851 21248
rect 15787 21188 15791 21244
rect 15791 21188 15847 21244
rect 15847 21188 15851 21244
rect 15787 21184 15851 21188
rect 15867 21244 15931 21248
rect 15867 21188 15871 21244
rect 15871 21188 15927 21244
rect 15927 21188 15931 21244
rect 15867 21184 15931 21188
rect 15947 21244 16011 21248
rect 15947 21188 15951 21244
rect 15951 21188 16007 21244
rect 16007 21188 16011 21244
rect 15947 21184 16011 21188
rect 16027 21244 16091 21248
rect 16027 21188 16031 21244
rect 16031 21188 16087 21244
rect 16087 21188 16091 21244
rect 16027 21184 16091 21188
rect 21721 21244 21785 21248
rect 21721 21188 21725 21244
rect 21725 21188 21781 21244
rect 21781 21188 21785 21244
rect 21721 21184 21785 21188
rect 21801 21244 21865 21248
rect 21801 21188 21805 21244
rect 21805 21188 21861 21244
rect 21861 21188 21865 21244
rect 21801 21184 21865 21188
rect 21881 21244 21945 21248
rect 21881 21188 21885 21244
rect 21885 21188 21941 21244
rect 21941 21188 21945 21244
rect 21881 21184 21945 21188
rect 21961 21244 22025 21248
rect 21961 21188 21965 21244
rect 21965 21188 22021 21244
rect 22021 21188 22025 21244
rect 21961 21184 22025 21188
rect 4476 20980 4540 21044
rect 1348 20844 1412 20908
rect 5396 20844 5460 20908
rect 6886 20700 6950 20704
rect 6886 20644 6890 20700
rect 6890 20644 6946 20700
rect 6946 20644 6950 20700
rect 6886 20640 6950 20644
rect 6966 20700 7030 20704
rect 6966 20644 6970 20700
rect 6970 20644 7026 20700
rect 7026 20644 7030 20700
rect 6966 20640 7030 20644
rect 7046 20700 7110 20704
rect 7046 20644 7050 20700
rect 7050 20644 7106 20700
rect 7106 20644 7110 20700
rect 7046 20640 7110 20644
rect 7126 20700 7190 20704
rect 7126 20644 7130 20700
rect 7130 20644 7186 20700
rect 7186 20644 7190 20700
rect 7126 20640 7190 20644
rect 12820 20700 12884 20704
rect 12820 20644 12824 20700
rect 12824 20644 12880 20700
rect 12880 20644 12884 20700
rect 12820 20640 12884 20644
rect 12900 20700 12964 20704
rect 12900 20644 12904 20700
rect 12904 20644 12960 20700
rect 12960 20644 12964 20700
rect 12900 20640 12964 20644
rect 12980 20700 13044 20704
rect 12980 20644 12984 20700
rect 12984 20644 13040 20700
rect 13040 20644 13044 20700
rect 12980 20640 13044 20644
rect 13060 20700 13124 20704
rect 13060 20644 13064 20700
rect 13064 20644 13120 20700
rect 13120 20644 13124 20700
rect 13060 20640 13124 20644
rect 18754 20700 18818 20704
rect 18754 20644 18758 20700
rect 18758 20644 18814 20700
rect 18814 20644 18818 20700
rect 18754 20640 18818 20644
rect 18834 20700 18898 20704
rect 18834 20644 18838 20700
rect 18838 20644 18894 20700
rect 18894 20644 18898 20700
rect 18834 20640 18898 20644
rect 18914 20700 18978 20704
rect 18914 20644 18918 20700
rect 18918 20644 18974 20700
rect 18974 20644 18978 20700
rect 18914 20640 18978 20644
rect 18994 20700 19058 20704
rect 18994 20644 18998 20700
rect 18998 20644 19054 20700
rect 19054 20644 19058 20700
rect 18994 20640 19058 20644
rect 24688 20700 24752 20704
rect 24688 20644 24692 20700
rect 24692 20644 24748 20700
rect 24748 20644 24752 20700
rect 24688 20640 24752 20644
rect 24768 20700 24832 20704
rect 24768 20644 24772 20700
rect 24772 20644 24828 20700
rect 24828 20644 24832 20700
rect 24768 20640 24832 20644
rect 24848 20700 24912 20704
rect 24848 20644 24852 20700
rect 24852 20644 24908 20700
rect 24908 20644 24912 20700
rect 24848 20640 24912 20644
rect 24928 20700 24992 20704
rect 24928 20644 24932 20700
rect 24932 20644 24988 20700
rect 24988 20644 24992 20700
rect 24928 20640 24992 20644
rect 3004 20224 3068 20228
rect 3004 20168 3018 20224
rect 3018 20168 3068 20224
rect 3004 20164 3068 20168
rect 9260 20300 9324 20364
rect 3919 20156 3983 20160
rect 3919 20100 3923 20156
rect 3923 20100 3979 20156
rect 3979 20100 3983 20156
rect 3919 20096 3983 20100
rect 3999 20156 4063 20160
rect 3999 20100 4003 20156
rect 4003 20100 4059 20156
rect 4059 20100 4063 20156
rect 3999 20096 4063 20100
rect 4079 20156 4143 20160
rect 4079 20100 4083 20156
rect 4083 20100 4139 20156
rect 4139 20100 4143 20156
rect 4079 20096 4143 20100
rect 4159 20156 4223 20160
rect 4159 20100 4163 20156
rect 4163 20100 4219 20156
rect 4219 20100 4223 20156
rect 4159 20096 4223 20100
rect 9853 20156 9917 20160
rect 9853 20100 9857 20156
rect 9857 20100 9913 20156
rect 9913 20100 9917 20156
rect 9853 20096 9917 20100
rect 9933 20156 9997 20160
rect 9933 20100 9937 20156
rect 9937 20100 9993 20156
rect 9993 20100 9997 20156
rect 9933 20096 9997 20100
rect 10013 20156 10077 20160
rect 10013 20100 10017 20156
rect 10017 20100 10073 20156
rect 10073 20100 10077 20156
rect 10013 20096 10077 20100
rect 10093 20156 10157 20160
rect 10093 20100 10097 20156
rect 10097 20100 10153 20156
rect 10153 20100 10157 20156
rect 10093 20096 10157 20100
rect 15787 20156 15851 20160
rect 15787 20100 15791 20156
rect 15791 20100 15847 20156
rect 15847 20100 15851 20156
rect 15787 20096 15851 20100
rect 15867 20156 15931 20160
rect 15867 20100 15871 20156
rect 15871 20100 15927 20156
rect 15927 20100 15931 20156
rect 15867 20096 15931 20100
rect 15947 20156 16011 20160
rect 15947 20100 15951 20156
rect 15951 20100 16007 20156
rect 16007 20100 16011 20156
rect 15947 20096 16011 20100
rect 16027 20156 16091 20160
rect 16027 20100 16031 20156
rect 16031 20100 16087 20156
rect 16087 20100 16091 20156
rect 16027 20096 16091 20100
rect 21721 20156 21785 20160
rect 21721 20100 21725 20156
rect 21725 20100 21781 20156
rect 21781 20100 21785 20156
rect 21721 20096 21785 20100
rect 21801 20156 21865 20160
rect 21801 20100 21805 20156
rect 21805 20100 21861 20156
rect 21861 20100 21865 20156
rect 21801 20096 21865 20100
rect 21881 20156 21945 20160
rect 21881 20100 21885 20156
rect 21885 20100 21941 20156
rect 21941 20100 21945 20156
rect 21881 20096 21945 20100
rect 21961 20156 22025 20160
rect 21961 20100 21965 20156
rect 21965 20100 22021 20156
rect 22021 20100 22025 20156
rect 21961 20096 22025 20100
rect 22508 19892 22572 19956
rect 22692 19816 22756 19820
rect 22692 19760 22742 19816
rect 22742 19760 22756 19816
rect 22692 19756 22756 19760
rect 10364 19620 10428 19684
rect 6886 19612 6950 19616
rect 6886 19556 6890 19612
rect 6890 19556 6946 19612
rect 6946 19556 6950 19612
rect 6886 19552 6950 19556
rect 6966 19612 7030 19616
rect 6966 19556 6970 19612
rect 6970 19556 7026 19612
rect 7026 19556 7030 19612
rect 6966 19552 7030 19556
rect 7046 19612 7110 19616
rect 7046 19556 7050 19612
rect 7050 19556 7106 19612
rect 7106 19556 7110 19612
rect 7046 19552 7110 19556
rect 7126 19612 7190 19616
rect 7126 19556 7130 19612
rect 7130 19556 7186 19612
rect 7186 19556 7190 19612
rect 7126 19552 7190 19556
rect 12820 19612 12884 19616
rect 12820 19556 12824 19612
rect 12824 19556 12880 19612
rect 12880 19556 12884 19612
rect 12820 19552 12884 19556
rect 12900 19612 12964 19616
rect 12900 19556 12904 19612
rect 12904 19556 12960 19612
rect 12960 19556 12964 19612
rect 12900 19552 12964 19556
rect 12980 19612 13044 19616
rect 12980 19556 12984 19612
rect 12984 19556 13040 19612
rect 13040 19556 13044 19612
rect 12980 19552 13044 19556
rect 13060 19612 13124 19616
rect 13060 19556 13064 19612
rect 13064 19556 13120 19612
rect 13120 19556 13124 19612
rect 13060 19552 13124 19556
rect 18754 19612 18818 19616
rect 18754 19556 18758 19612
rect 18758 19556 18814 19612
rect 18814 19556 18818 19612
rect 18754 19552 18818 19556
rect 18834 19612 18898 19616
rect 18834 19556 18838 19612
rect 18838 19556 18894 19612
rect 18894 19556 18898 19612
rect 18834 19552 18898 19556
rect 18914 19612 18978 19616
rect 18914 19556 18918 19612
rect 18918 19556 18974 19612
rect 18974 19556 18978 19612
rect 18914 19552 18978 19556
rect 18994 19612 19058 19616
rect 18994 19556 18998 19612
rect 18998 19556 19054 19612
rect 19054 19556 19058 19612
rect 18994 19552 19058 19556
rect 24688 19612 24752 19616
rect 24688 19556 24692 19612
rect 24692 19556 24748 19612
rect 24748 19556 24752 19612
rect 24688 19552 24752 19556
rect 24768 19612 24832 19616
rect 24768 19556 24772 19612
rect 24772 19556 24828 19612
rect 24828 19556 24832 19612
rect 24768 19552 24832 19556
rect 24848 19612 24912 19616
rect 24848 19556 24852 19612
rect 24852 19556 24908 19612
rect 24908 19556 24912 19612
rect 24848 19552 24912 19556
rect 24928 19612 24992 19616
rect 24928 19556 24932 19612
rect 24932 19556 24988 19612
rect 24988 19556 24992 19612
rect 24928 19552 24992 19556
rect 3919 19068 3983 19072
rect 3919 19012 3923 19068
rect 3923 19012 3979 19068
rect 3979 19012 3983 19068
rect 3919 19008 3983 19012
rect 3999 19068 4063 19072
rect 3999 19012 4003 19068
rect 4003 19012 4059 19068
rect 4059 19012 4063 19068
rect 3999 19008 4063 19012
rect 4079 19068 4143 19072
rect 4079 19012 4083 19068
rect 4083 19012 4139 19068
rect 4139 19012 4143 19068
rect 4079 19008 4143 19012
rect 4159 19068 4223 19072
rect 4159 19012 4163 19068
rect 4163 19012 4219 19068
rect 4219 19012 4223 19068
rect 4159 19008 4223 19012
rect 2452 18804 2516 18868
rect 9853 19068 9917 19072
rect 9853 19012 9857 19068
rect 9857 19012 9913 19068
rect 9913 19012 9917 19068
rect 9853 19008 9917 19012
rect 9933 19068 9997 19072
rect 9933 19012 9937 19068
rect 9937 19012 9993 19068
rect 9993 19012 9997 19068
rect 9933 19008 9997 19012
rect 10013 19068 10077 19072
rect 10013 19012 10017 19068
rect 10017 19012 10073 19068
rect 10073 19012 10077 19068
rect 10013 19008 10077 19012
rect 10093 19068 10157 19072
rect 10093 19012 10097 19068
rect 10097 19012 10153 19068
rect 10153 19012 10157 19068
rect 10093 19008 10157 19012
rect 15787 19068 15851 19072
rect 15787 19012 15791 19068
rect 15791 19012 15847 19068
rect 15847 19012 15851 19068
rect 15787 19008 15851 19012
rect 15867 19068 15931 19072
rect 15867 19012 15871 19068
rect 15871 19012 15927 19068
rect 15927 19012 15931 19068
rect 15867 19008 15931 19012
rect 15947 19068 16011 19072
rect 15947 19012 15951 19068
rect 15951 19012 16007 19068
rect 16007 19012 16011 19068
rect 15947 19008 16011 19012
rect 16027 19068 16091 19072
rect 16027 19012 16031 19068
rect 16031 19012 16087 19068
rect 16087 19012 16091 19068
rect 16027 19008 16091 19012
rect 21721 19068 21785 19072
rect 21721 19012 21725 19068
rect 21725 19012 21781 19068
rect 21781 19012 21785 19068
rect 21721 19008 21785 19012
rect 21801 19068 21865 19072
rect 21801 19012 21805 19068
rect 21805 19012 21861 19068
rect 21861 19012 21865 19068
rect 21801 19008 21865 19012
rect 21881 19068 21945 19072
rect 21881 19012 21885 19068
rect 21885 19012 21941 19068
rect 21941 19012 21945 19068
rect 21881 19008 21945 19012
rect 21961 19068 22025 19072
rect 21961 19012 21965 19068
rect 21965 19012 22021 19068
rect 22021 19012 22025 19068
rect 21961 19008 22025 19012
rect 11652 19000 11716 19004
rect 11652 18944 11666 19000
rect 11666 18944 11716 19000
rect 11652 18940 11716 18944
rect 17172 19000 17236 19004
rect 17172 18944 17186 19000
rect 17186 18944 17236 19000
rect 17172 18940 17236 18944
rect 13676 18728 13740 18732
rect 13676 18672 13690 18728
rect 13690 18672 13740 18728
rect 13676 18668 13740 18672
rect 6886 18524 6950 18528
rect 6886 18468 6890 18524
rect 6890 18468 6946 18524
rect 6946 18468 6950 18524
rect 6886 18464 6950 18468
rect 6966 18524 7030 18528
rect 6966 18468 6970 18524
rect 6970 18468 7026 18524
rect 7026 18468 7030 18524
rect 6966 18464 7030 18468
rect 7046 18524 7110 18528
rect 7046 18468 7050 18524
rect 7050 18468 7106 18524
rect 7106 18468 7110 18524
rect 7046 18464 7110 18468
rect 7126 18524 7190 18528
rect 7126 18468 7130 18524
rect 7130 18468 7186 18524
rect 7186 18468 7190 18524
rect 7126 18464 7190 18468
rect 12820 18524 12884 18528
rect 12820 18468 12824 18524
rect 12824 18468 12880 18524
rect 12880 18468 12884 18524
rect 12820 18464 12884 18468
rect 12900 18524 12964 18528
rect 12900 18468 12904 18524
rect 12904 18468 12960 18524
rect 12960 18468 12964 18524
rect 12900 18464 12964 18468
rect 12980 18524 13044 18528
rect 12980 18468 12984 18524
rect 12984 18468 13040 18524
rect 13040 18468 13044 18524
rect 12980 18464 13044 18468
rect 13060 18524 13124 18528
rect 13060 18468 13064 18524
rect 13064 18468 13120 18524
rect 13120 18468 13124 18524
rect 13060 18464 13124 18468
rect 18754 18524 18818 18528
rect 18754 18468 18758 18524
rect 18758 18468 18814 18524
rect 18814 18468 18818 18524
rect 18754 18464 18818 18468
rect 18834 18524 18898 18528
rect 18834 18468 18838 18524
rect 18838 18468 18894 18524
rect 18894 18468 18898 18524
rect 18834 18464 18898 18468
rect 18914 18524 18978 18528
rect 18914 18468 18918 18524
rect 18918 18468 18974 18524
rect 18974 18468 18978 18524
rect 18914 18464 18978 18468
rect 18994 18524 19058 18528
rect 18994 18468 18998 18524
rect 18998 18468 19054 18524
rect 19054 18468 19058 18524
rect 18994 18464 19058 18468
rect 24688 18524 24752 18528
rect 24688 18468 24692 18524
rect 24692 18468 24748 18524
rect 24748 18468 24752 18524
rect 24688 18464 24752 18468
rect 24768 18524 24832 18528
rect 24768 18468 24772 18524
rect 24772 18468 24828 18524
rect 24828 18468 24832 18524
rect 24768 18464 24832 18468
rect 24848 18524 24912 18528
rect 24848 18468 24852 18524
rect 24852 18468 24908 18524
rect 24908 18468 24912 18524
rect 24848 18464 24912 18468
rect 24928 18524 24992 18528
rect 24928 18468 24932 18524
rect 24932 18468 24988 18524
rect 24988 18468 24992 18524
rect 24928 18464 24992 18468
rect 2636 18456 2700 18460
rect 2636 18400 2650 18456
rect 2650 18400 2700 18456
rect 2636 18396 2700 18400
rect 5396 18456 5460 18460
rect 5396 18400 5410 18456
rect 5410 18400 5460 18456
rect 5396 18396 5460 18400
rect 4844 18124 4908 18188
rect 16988 18124 17052 18188
rect 20852 18124 20916 18188
rect 14596 17988 14660 18052
rect 15516 17988 15580 18052
rect 20852 17988 20916 18052
rect 3919 17980 3983 17984
rect 3919 17924 3923 17980
rect 3923 17924 3979 17980
rect 3979 17924 3983 17980
rect 3919 17920 3983 17924
rect 3999 17980 4063 17984
rect 3999 17924 4003 17980
rect 4003 17924 4059 17980
rect 4059 17924 4063 17980
rect 3999 17920 4063 17924
rect 4079 17980 4143 17984
rect 4079 17924 4083 17980
rect 4083 17924 4139 17980
rect 4139 17924 4143 17980
rect 4079 17920 4143 17924
rect 4159 17980 4223 17984
rect 4159 17924 4163 17980
rect 4163 17924 4219 17980
rect 4219 17924 4223 17980
rect 4159 17920 4223 17924
rect 9853 17980 9917 17984
rect 9853 17924 9857 17980
rect 9857 17924 9913 17980
rect 9913 17924 9917 17980
rect 9853 17920 9917 17924
rect 9933 17980 9997 17984
rect 9933 17924 9937 17980
rect 9937 17924 9993 17980
rect 9993 17924 9997 17980
rect 9933 17920 9997 17924
rect 10013 17980 10077 17984
rect 10013 17924 10017 17980
rect 10017 17924 10073 17980
rect 10073 17924 10077 17980
rect 10013 17920 10077 17924
rect 10093 17980 10157 17984
rect 10093 17924 10097 17980
rect 10097 17924 10153 17980
rect 10153 17924 10157 17980
rect 10093 17920 10157 17924
rect 15787 17980 15851 17984
rect 15787 17924 15791 17980
rect 15791 17924 15847 17980
rect 15847 17924 15851 17980
rect 15787 17920 15851 17924
rect 15867 17980 15931 17984
rect 15867 17924 15871 17980
rect 15871 17924 15927 17980
rect 15927 17924 15931 17980
rect 15867 17920 15931 17924
rect 15947 17980 16011 17984
rect 15947 17924 15951 17980
rect 15951 17924 16007 17980
rect 16007 17924 16011 17980
rect 15947 17920 16011 17924
rect 16027 17980 16091 17984
rect 16027 17924 16031 17980
rect 16031 17924 16087 17980
rect 16087 17924 16091 17980
rect 16027 17920 16091 17924
rect 21721 17980 21785 17984
rect 21721 17924 21725 17980
rect 21725 17924 21781 17980
rect 21781 17924 21785 17980
rect 21721 17920 21785 17924
rect 21801 17980 21865 17984
rect 21801 17924 21805 17980
rect 21805 17924 21861 17980
rect 21861 17924 21865 17980
rect 21801 17920 21865 17924
rect 21881 17980 21945 17984
rect 21881 17924 21885 17980
rect 21885 17924 21941 17980
rect 21941 17924 21945 17980
rect 21881 17920 21945 17924
rect 21961 17980 22025 17984
rect 21961 17924 21965 17980
rect 21965 17924 22021 17980
rect 22021 17924 22025 17980
rect 21961 17920 22025 17924
rect 10732 17852 10796 17916
rect 12020 17852 12084 17916
rect 2084 17308 2148 17372
rect 19748 17852 19812 17916
rect 17724 17716 17788 17780
rect 21220 17444 21284 17508
rect 6886 17436 6950 17440
rect 6886 17380 6890 17436
rect 6890 17380 6946 17436
rect 6946 17380 6950 17436
rect 6886 17376 6950 17380
rect 6966 17436 7030 17440
rect 6966 17380 6970 17436
rect 6970 17380 7026 17436
rect 7026 17380 7030 17436
rect 6966 17376 7030 17380
rect 7046 17436 7110 17440
rect 7046 17380 7050 17436
rect 7050 17380 7106 17436
rect 7106 17380 7110 17436
rect 7046 17376 7110 17380
rect 7126 17436 7190 17440
rect 7126 17380 7130 17436
rect 7130 17380 7186 17436
rect 7186 17380 7190 17436
rect 7126 17376 7190 17380
rect 12820 17436 12884 17440
rect 12820 17380 12824 17436
rect 12824 17380 12880 17436
rect 12880 17380 12884 17436
rect 12820 17376 12884 17380
rect 12900 17436 12964 17440
rect 12900 17380 12904 17436
rect 12904 17380 12960 17436
rect 12960 17380 12964 17436
rect 12900 17376 12964 17380
rect 12980 17436 13044 17440
rect 12980 17380 12984 17436
rect 12984 17380 13040 17436
rect 13040 17380 13044 17436
rect 12980 17376 13044 17380
rect 13060 17436 13124 17440
rect 13060 17380 13064 17436
rect 13064 17380 13120 17436
rect 13120 17380 13124 17436
rect 13060 17376 13124 17380
rect 18754 17436 18818 17440
rect 18754 17380 18758 17436
rect 18758 17380 18814 17436
rect 18814 17380 18818 17436
rect 18754 17376 18818 17380
rect 18834 17436 18898 17440
rect 18834 17380 18838 17436
rect 18838 17380 18894 17436
rect 18894 17380 18898 17436
rect 18834 17376 18898 17380
rect 18914 17436 18978 17440
rect 18914 17380 18918 17436
rect 18918 17380 18974 17436
rect 18974 17380 18978 17436
rect 18914 17376 18978 17380
rect 18994 17436 19058 17440
rect 18994 17380 18998 17436
rect 18998 17380 19054 17436
rect 19054 17380 19058 17436
rect 18994 17376 19058 17380
rect 24688 17436 24752 17440
rect 24688 17380 24692 17436
rect 24692 17380 24748 17436
rect 24748 17380 24752 17436
rect 24688 17376 24752 17380
rect 24768 17436 24832 17440
rect 24768 17380 24772 17436
rect 24772 17380 24828 17436
rect 24828 17380 24832 17436
rect 24768 17376 24832 17380
rect 24848 17436 24912 17440
rect 24848 17380 24852 17436
rect 24852 17380 24908 17436
rect 24908 17380 24912 17436
rect 24848 17376 24912 17380
rect 24928 17436 24992 17440
rect 24928 17380 24932 17436
rect 24932 17380 24988 17436
rect 24988 17380 24992 17436
rect 24928 17376 24992 17380
rect 3919 16892 3983 16896
rect 3919 16836 3923 16892
rect 3923 16836 3979 16892
rect 3979 16836 3983 16892
rect 3919 16832 3983 16836
rect 3999 16892 4063 16896
rect 3999 16836 4003 16892
rect 4003 16836 4059 16892
rect 4059 16836 4063 16892
rect 3999 16832 4063 16836
rect 4079 16892 4143 16896
rect 4079 16836 4083 16892
rect 4083 16836 4139 16892
rect 4139 16836 4143 16892
rect 4079 16832 4143 16836
rect 4159 16892 4223 16896
rect 4159 16836 4163 16892
rect 4163 16836 4219 16892
rect 4219 16836 4223 16892
rect 4159 16832 4223 16836
rect 9853 16892 9917 16896
rect 9853 16836 9857 16892
rect 9857 16836 9913 16892
rect 9913 16836 9917 16892
rect 9853 16832 9917 16836
rect 9933 16892 9997 16896
rect 9933 16836 9937 16892
rect 9937 16836 9993 16892
rect 9993 16836 9997 16892
rect 9933 16832 9997 16836
rect 10013 16892 10077 16896
rect 10013 16836 10017 16892
rect 10017 16836 10073 16892
rect 10073 16836 10077 16892
rect 10013 16832 10077 16836
rect 10093 16892 10157 16896
rect 10093 16836 10097 16892
rect 10097 16836 10153 16892
rect 10153 16836 10157 16892
rect 10093 16832 10157 16836
rect 15787 16892 15851 16896
rect 15787 16836 15791 16892
rect 15791 16836 15847 16892
rect 15847 16836 15851 16892
rect 15787 16832 15851 16836
rect 15867 16892 15931 16896
rect 15867 16836 15871 16892
rect 15871 16836 15927 16892
rect 15927 16836 15931 16892
rect 15867 16832 15931 16836
rect 15947 16892 16011 16896
rect 15947 16836 15951 16892
rect 15951 16836 16007 16892
rect 16007 16836 16011 16892
rect 15947 16832 16011 16836
rect 16027 16892 16091 16896
rect 16027 16836 16031 16892
rect 16031 16836 16087 16892
rect 16087 16836 16091 16892
rect 16027 16832 16091 16836
rect 21721 16892 21785 16896
rect 21721 16836 21725 16892
rect 21725 16836 21781 16892
rect 21781 16836 21785 16892
rect 21721 16832 21785 16836
rect 21801 16892 21865 16896
rect 21801 16836 21805 16892
rect 21805 16836 21861 16892
rect 21861 16836 21865 16892
rect 21801 16832 21865 16836
rect 21881 16892 21945 16896
rect 21881 16836 21885 16892
rect 21885 16836 21941 16892
rect 21941 16836 21945 16892
rect 21881 16832 21945 16836
rect 21961 16892 22025 16896
rect 21961 16836 21965 16892
rect 21965 16836 22021 16892
rect 22021 16836 22025 16892
rect 21961 16832 22025 16836
rect 1900 16824 1964 16828
rect 1900 16768 1914 16824
rect 1914 16768 1964 16824
rect 1900 16764 1964 16768
rect 7972 16492 8036 16556
rect 20300 16356 20364 16420
rect 6886 16348 6950 16352
rect 6886 16292 6890 16348
rect 6890 16292 6946 16348
rect 6946 16292 6950 16348
rect 6886 16288 6950 16292
rect 6966 16348 7030 16352
rect 6966 16292 6970 16348
rect 6970 16292 7026 16348
rect 7026 16292 7030 16348
rect 6966 16288 7030 16292
rect 7046 16348 7110 16352
rect 7046 16292 7050 16348
rect 7050 16292 7106 16348
rect 7106 16292 7110 16348
rect 7046 16288 7110 16292
rect 7126 16348 7190 16352
rect 7126 16292 7130 16348
rect 7130 16292 7186 16348
rect 7186 16292 7190 16348
rect 7126 16288 7190 16292
rect 12820 16348 12884 16352
rect 12820 16292 12824 16348
rect 12824 16292 12880 16348
rect 12880 16292 12884 16348
rect 12820 16288 12884 16292
rect 12900 16348 12964 16352
rect 12900 16292 12904 16348
rect 12904 16292 12960 16348
rect 12960 16292 12964 16348
rect 12900 16288 12964 16292
rect 12980 16348 13044 16352
rect 12980 16292 12984 16348
rect 12984 16292 13040 16348
rect 13040 16292 13044 16348
rect 12980 16288 13044 16292
rect 13060 16348 13124 16352
rect 13060 16292 13064 16348
rect 13064 16292 13120 16348
rect 13120 16292 13124 16348
rect 13060 16288 13124 16292
rect 18754 16348 18818 16352
rect 18754 16292 18758 16348
rect 18758 16292 18814 16348
rect 18814 16292 18818 16348
rect 18754 16288 18818 16292
rect 18834 16348 18898 16352
rect 18834 16292 18838 16348
rect 18838 16292 18894 16348
rect 18894 16292 18898 16348
rect 18834 16288 18898 16292
rect 18914 16348 18978 16352
rect 18914 16292 18918 16348
rect 18918 16292 18974 16348
rect 18974 16292 18978 16348
rect 18914 16288 18978 16292
rect 18994 16348 19058 16352
rect 18994 16292 18998 16348
rect 18998 16292 19054 16348
rect 19054 16292 19058 16348
rect 18994 16288 19058 16292
rect 24688 16348 24752 16352
rect 24688 16292 24692 16348
rect 24692 16292 24748 16348
rect 24748 16292 24752 16348
rect 24688 16288 24752 16292
rect 24768 16348 24832 16352
rect 24768 16292 24772 16348
rect 24772 16292 24828 16348
rect 24828 16292 24832 16348
rect 24768 16288 24832 16292
rect 24848 16348 24912 16352
rect 24848 16292 24852 16348
rect 24852 16292 24908 16348
rect 24908 16292 24912 16348
rect 24848 16288 24912 16292
rect 24928 16348 24992 16352
rect 24928 16292 24932 16348
rect 24932 16292 24988 16348
rect 24988 16292 24992 16348
rect 24928 16288 24992 16292
rect 3556 16220 3620 16284
rect 15516 15948 15580 16012
rect 3919 15804 3983 15808
rect 3919 15748 3923 15804
rect 3923 15748 3979 15804
rect 3979 15748 3983 15804
rect 3919 15744 3983 15748
rect 3999 15804 4063 15808
rect 3999 15748 4003 15804
rect 4003 15748 4059 15804
rect 4059 15748 4063 15804
rect 3999 15744 4063 15748
rect 4079 15804 4143 15808
rect 4079 15748 4083 15804
rect 4083 15748 4139 15804
rect 4139 15748 4143 15804
rect 4079 15744 4143 15748
rect 4159 15804 4223 15808
rect 4159 15748 4163 15804
rect 4163 15748 4219 15804
rect 4219 15748 4223 15804
rect 4159 15744 4223 15748
rect 9853 15804 9917 15808
rect 9853 15748 9857 15804
rect 9857 15748 9913 15804
rect 9913 15748 9917 15804
rect 9853 15744 9917 15748
rect 9933 15804 9997 15808
rect 9933 15748 9937 15804
rect 9937 15748 9993 15804
rect 9993 15748 9997 15804
rect 9933 15744 9997 15748
rect 10013 15804 10077 15808
rect 10013 15748 10017 15804
rect 10017 15748 10073 15804
rect 10073 15748 10077 15804
rect 10013 15744 10077 15748
rect 10093 15804 10157 15808
rect 10093 15748 10097 15804
rect 10097 15748 10153 15804
rect 10153 15748 10157 15804
rect 10093 15744 10157 15748
rect 15787 15804 15851 15808
rect 15787 15748 15791 15804
rect 15791 15748 15847 15804
rect 15847 15748 15851 15804
rect 15787 15744 15851 15748
rect 15867 15804 15931 15808
rect 15867 15748 15871 15804
rect 15871 15748 15927 15804
rect 15927 15748 15931 15804
rect 15867 15744 15931 15748
rect 15947 15804 16011 15808
rect 15947 15748 15951 15804
rect 15951 15748 16007 15804
rect 16007 15748 16011 15804
rect 15947 15744 16011 15748
rect 16027 15804 16091 15808
rect 16027 15748 16031 15804
rect 16031 15748 16087 15804
rect 16087 15748 16091 15804
rect 16027 15744 16091 15748
rect 21721 15804 21785 15808
rect 21721 15748 21725 15804
rect 21725 15748 21781 15804
rect 21781 15748 21785 15804
rect 21721 15744 21785 15748
rect 21801 15804 21865 15808
rect 21801 15748 21805 15804
rect 21805 15748 21861 15804
rect 21861 15748 21865 15804
rect 21801 15744 21865 15748
rect 21881 15804 21945 15808
rect 21881 15748 21885 15804
rect 21885 15748 21941 15804
rect 21941 15748 21945 15804
rect 21881 15744 21945 15748
rect 21961 15804 22025 15808
rect 21961 15748 21965 15804
rect 21965 15748 22021 15804
rect 22021 15748 22025 15804
rect 21961 15744 22025 15748
rect 3372 15540 3436 15604
rect 14412 15404 14476 15468
rect 6886 15260 6950 15264
rect 6886 15204 6890 15260
rect 6890 15204 6946 15260
rect 6946 15204 6950 15260
rect 6886 15200 6950 15204
rect 6966 15260 7030 15264
rect 6966 15204 6970 15260
rect 6970 15204 7026 15260
rect 7026 15204 7030 15260
rect 6966 15200 7030 15204
rect 7046 15260 7110 15264
rect 7046 15204 7050 15260
rect 7050 15204 7106 15260
rect 7106 15204 7110 15260
rect 7046 15200 7110 15204
rect 7126 15260 7190 15264
rect 7126 15204 7130 15260
rect 7130 15204 7186 15260
rect 7186 15204 7190 15260
rect 7126 15200 7190 15204
rect 12820 15260 12884 15264
rect 12820 15204 12824 15260
rect 12824 15204 12880 15260
rect 12880 15204 12884 15260
rect 12820 15200 12884 15204
rect 12900 15260 12964 15264
rect 12900 15204 12904 15260
rect 12904 15204 12960 15260
rect 12960 15204 12964 15260
rect 12900 15200 12964 15204
rect 12980 15260 13044 15264
rect 12980 15204 12984 15260
rect 12984 15204 13040 15260
rect 13040 15204 13044 15260
rect 12980 15200 13044 15204
rect 13060 15260 13124 15264
rect 13060 15204 13064 15260
rect 13064 15204 13120 15260
rect 13120 15204 13124 15260
rect 13060 15200 13124 15204
rect 18754 15260 18818 15264
rect 18754 15204 18758 15260
rect 18758 15204 18814 15260
rect 18814 15204 18818 15260
rect 18754 15200 18818 15204
rect 18834 15260 18898 15264
rect 18834 15204 18838 15260
rect 18838 15204 18894 15260
rect 18894 15204 18898 15260
rect 18834 15200 18898 15204
rect 18914 15260 18978 15264
rect 18914 15204 18918 15260
rect 18918 15204 18974 15260
rect 18974 15204 18978 15260
rect 18914 15200 18978 15204
rect 18994 15260 19058 15264
rect 18994 15204 18998 15260
rect 18998 15204 19054 15260
rect 19054 15204 19058 15260
rect 18994 15200 19058 15204
rect 24688 15260 24752 15264
rect 24688 15204 24692 15260
rect 24692 15204 24748 15260
rect 24748 15204 24752 15260
rect 24688 15200 24752 15204
rect 24768 15260 24832 15264
rect 24768 15204 24772 15260
rect 24772 15204 24828 15260
rect 24828 15204 24832 15260
rect 24768 15200 24832 15204
rect 24848 15260 24912 15264
rect 24848 15204 24852 15260
rect 24852 15204 24908 15260
rect 24908 15204 24912 15260
rect 24848 15200 24912 15204
rect 24928 15260 24992 15264
rect 24928 15204 24932 15260
rect 24932 15204 24988 15260
rect 24988 15204 24992 15260
rect 24928 15200 24992 15204
rect 4660 15192 4724 15196
rect 4660 15136 4674 15192
rect 4674 15136 4724 15192
rect 4660 15132 4724 15136
rect 11652 15132 11716 15196
rect 16252 15192 16316 15196
rect 16252 15136 16266 15192
rect 16266 15136 16316 15192
rect 16252 15132 16316 15136
rect 5948 14724 6012 14788
rect 3919 14716 3983 14720
rect 3919 14660 3923 14716
rect 3923 14660 3979 14716
rect 3979 14660 3983 14716
rect 3919 14656 3983 14660
rect 3999 14716 4063 14720
rect 3999 14660 4003 14716
rect 4003 14660 4059 14716
rect 4059 14660 4063 14716
rect 3999 14656 4063 14660
rect 4079 14716 4143 14720
rect 4079 14660 4083 14716
rect 4083 14660 4139 14716
rect 4139 14660 4143 14716
rect 4079 14656 4143 14660
rect 4159 14716 4223 14720
rect 4159 14660 4163 14716
rect 4163 14660 4219 14716
rect 4219 14660 4223 14716
rect 4159 14656 4223 14660
rect 9853 14716 9917 14720
rect 9853 14660 9857 14716
rect 9857 14660 9913 14716
rect 9913 14660 9917 14716
rect 9853 14656 9917 14660
rect 9933 14716 9997 14720
rect 9933 14660 9937 14716
rect 9937 14660 9993 14716
rect 9993 14660 9997 14716
rect 9933 14656 9997 14660
rect 10013 14716 10077 14720
rect 10013 14660 10017 14716
rect 10017 14660 10073 14716
rect 10073 14660 10077 14716
rect 10013 14656 10077 14660
rect 10093 14716 10157 14720
rect 10093 14660 10097 14716
rect 10097 14660 10153 14716
rect 10153 14660 10157 14716
rect 10093 14656 10157 14660
rect 15787 14716 15851 14720
rect 15787 14660 15791 14716
rect 15791 14660 15847 14716
rect 15847 14660 15851 14716
rect 15787 14656 15851 14660
rect 15867 14716 15931 14720
rect 15867 14660 15871 14716
rect 15871 14660 15927 14716
rect 15927 14660 15931 14716
rect 15867 14656 15931 14660
rect 15947 14716 16011 14720
rect 15947 14660 15951 14716
rect 15951 14660 16007 14716
rect 16007 14660 16011 14716
rect 15947 14656 16011 14660
rect 16027 14716 16091 14720
rect 16027 14660 16031 14716
rect 16031 14660 16087 14716
rect 16087 14660 16091 14716
rect 16027 14656 16091 14660
rect 21721 14716 21785 14720
rect 21721 14660 21725 14716
rect 21725 14660 21781 14716
rect 21781 14660 21785 14716
rect 21721 14656 21785 14660
rect 21801 14716 21865 14720
rect 21801 14660 21805 14716
rect 21805 14660 21861 14716
rect 21861 14660 21865 14716
rect 21801 14656 21865 14660
rect 21881 14716 21945 14720
rect 21881 14660 21885 14716
rect 21885 14660 21941 14716
rect 21941 14660 21945 14716
rect 21881 14656 21945 14660
rect 21961 14716 22025 14720
rect 21961 14660 21965 14716
rect 21965 14660 22021 14716
rect 22021 14660 22025 14716
rect 21961 14656 22025 14660
rect 6132 14588 6196 14652
rect 6886 14172 6950 14176
rect 6886 14116 6890 14172
rect 6890 14116 6946 14172
rect 6946 14116 6950 14172
rect 6886 14112 6950 14116
rect 6966 14172 7030 14176
rect 6966 14116 6970 14172
rect 6970 14116 7026 14172
rect 7026 14116 7030 14172
rect 6966 14112 7030 14116
rect 7046 14172 7110 14176
rect 7046 14116 7050 14172
rect 7050 14116 7106 14172
rect 7106 14116 7110 14172
rect 7046 14112 7110 14116
rect 7126 14172 7190 14176
rect 7126 14116 7130 14172
rect 7130 14116 7186 14172
rect 7186 14116 7190 14172
rect 7126 14112 7190 14116
rect 12820 14172 12884 14176
rect 12820 14116 12824 14172
rect 12824 14116 12880 14172
rect 12880 14116 12884 14172
rect 12820 14112 12884 14116
rect 12900 14172 12964 14176
rect 12900 14116 12904 14172
rect 12904 14116 12960 14172
rect 12960 14116 12964 14172
rect 12900 14112 12964 14116
rect 12980 14172 13044 14176
rect 12980 14116 12984 14172
rect 12984 14116 13040 14172
rect 13040 14116 13044 14172
rect 12980 14112 13044 14116
rect 13060 14172 13124 14176
rect 13060 14116 13064 14172
rect 13064 14116 13120 14172
rect 13120 14116 13124 14172
rect 13060 14112 13124 14116
rect 18754 14172 18818 14176
rect 18754 14116 18758 14172
rect 18758 14116 18814 14172
rect 18814 14116 18818 14172
rect 18754 14112 18818 14116
rect 18834 14172 18898 14176
rect 18834 14116 18838 14172
rect 18838 14116 18894 14172
rect 18894 14116 18898 14172
rect 18834 14112 18898 14116
rect 18914 14172 18978 14176
rect 18914 14116 18918 14172
rect 18918 14116 18974 14172
rect 18974 14116 18978 14172
rect 18914 14112 18978 14116
rect 18994 14172 19058 14176
rect 18994 14116 18998 14172
rect 18998 14116 19054 14172
rect 19054 14116 19058 14172
rect 18994 14112 19058 14116
rect 24688 14172 24752 14176
rect 24688 14116 24692 14172
rect 24692 14116 24748 14172
rect 24748 14116 24752 14172
rect 24688 14112 24752 14116
rect 24768 14172 24832 14176
rect 24768 14116 24772 14172
rect 24772 14116 24828 14172
rect 24828 14116 24832 14172
rect 24768 14112 24832 14116
rect 24848 14172 24912 14176
rect 24848 14116 24852 14172
rect 24852 14116 24908 14172
rect 24908 14116 24912 14172
rect 24848 14112 24912 14116
rect 24928 14172 24992 14176
rect 24928 14116 24932 14172
rect 24932 14116 24988 14172
rect 24988 14116 24992 14172
rect 24928 14112 24992 14116
rect 5396 13908 5460 13972
rect 10916 13636 10980 13700
rect 22324 13636 22388 13700
rect 3919 13628 3983 13632
rect 3919 13572 3923 13628
rect 3923 13572 3979 13628
rect 3979 13572 3983 13628
rect 3919 13568 3983 13572
rect 3999 13628 4063 13632
rect 3999 13572 4003 13628
rect 4003 13572 4059 13628
rect 4059 13572 4063 13628
rect 3999 13568 4063 13572
rect 4079 13628 4143 13632
rect 4079 13572 4083 13628
rect 4083 13572 4139 13628
rect 4139 13572 4143 13628
rect 4079 13568 4143 13572
rect 4159 13628 4223 13632
rect 4159 13572 4163 13628
rect 4163 13572 4219 13628
rect 4219 13572 4223 13628
rect 4159 13568 4223 13572
rect 9853 13628 9917 13632
rect 9853 13572 9857 13628
rect 9857 13572 9913 13628
rect 9913 13572 9917 13628
rect 9853 13568 9917 13572
rect 9933 13628 9997 13632
rect 9933 13572 9937 13628
rect 9937 13572 9993 13628
rect 9993 13572 9997 13628
rect 9933 13568 9997 13572
rect 10013 13628 10077 13632
rect 10013 13572 10017 13628
rect 10017 13572 10073 13628
rect 10073 13572 10077 13628
rect 10013 13568 10077 13572
rect 10093 13628 10157 13632
rect 10093 13572 10097 13628
rect 10097 13572 10153 13628
rect 10153 13572 10157 13628
rect 10093 13568 10157 13572
rect 15787 13628 15851 13632
rect 15787 13572 15791 13628
rect 15791 13572 15847 13628
rect 15847 13572 15851 13628
rect 15787 13568 15851 13572
rect 15867 13628 15931 13632
rect 15867 13572 15871 13628
rect 15871 13572 15927 13628
rect 15927 13572 15931 13628
rect 15867 13568 15931 13572
rect 15947 13628 16011 13632
rect 15947 13572 15951 13628
rect 15951 13572 16007 13628
rect 16007 13572 16011 13628
rect 15947 13568 16011 13572
rect 16027 13628 16091 13632
rect 16027 13572 16031 13628
rect 16031 13572 16087 13628
rect 16087 13572 16091 13628
rect 16027 13568 16091 13572
rect 21721 13628 21785 13632
rect 21721 13572 21725 13628
rect 21725 13572 21781 13628
rect 21781 13572 21785 13628
rect 21721 13568 21785 13572
rect 21801 13628 21865 13632
rect 21801 13572 21805 13628
rect 21805 13572 21861 13628
rect 21861 13572 21865 13628
rect 21801 13568 21865 13572
rect 21881 13628 21945 13632
rect 21881 13572 21885 13628
rect 21885 13572 21941 13628
rect 21941 13572 21945 13628
rect 21881 13568 21945 13572
rect 21961 13628 22025 13632
rect 21961 13572 21965 13628
rect 21965 13572 22021 13628
rect 22021 13572 22025 13628
rect 21961 13568 22025 13572
rect 5948 13560 6012 13564
rect 5948 13504 5962 13560
rect 5962 13504 6012 13560
rect 5948 13500 6012 13504
rect 3556 13228 3620 13292
rect 12388 13288 12452 13292
rect 12388 13232 12438 13288
rect 12438 13232 12452 13288
rect 12388 13228 12452 13232
rect 6886 13084 6950 13088
rect 6886 13028 6890 13084
rect 6890 13028 6946 13084
rect 6946 13028 6950 13084
rect 6886 13024 6950 13028
rect 6966 13084 7030 13088
rect 6966 13028 6970 13084
rect 6970 13028 7026 13084
rect 7026 13028 7030 13084
rect 6966 13024 7030 13028
rect 7046 13084 7110 13088
rect 7046 13028 7050 13084
rect 7050 13028 7106 13084
rect 7106 13028 7110 13084
rect 7046 13024 7110 13028
rect 7126 13084 7190 13088
rect 7126 13028 7130 13084
rect 7130 13028 7186 13084
rect 7186 13028 7190 13084
rect 7126 13024 7190 13028
rect 12820 13084 12884 13088
rect 12820 13028 12824 13084
rect 12824 13028 12880 13084
rect 12880 13028 12884 13084
rect 12820 13024 12884 13028
rect 12900 13084 12964 13088
rect 12900 13028 12904 13084
rect 12904 13028 12960 13084
rect 12960 13028 12964 13084
rect 12900 13024 12964 13028
rect 12980 13084 13044 13088
rect 12980 13028 12984 13084
rect 12984 13028 13040 13084
rect 13040 13028 13044 13084
rect 12980 13024 13044 13028
rect 13060 13084 13124 13088
rect 13060 13028 13064 13084
rect 13064 13028 13120 13084
rect 13120 13028 13124 13084
rect 13060 13024 13124 13028
rect 18754 13084 18818 13088
rect 18754 13028 18758 13084
rect 18758 13028 18814 13084
rect 18814 13028 18818 13084
rect 18754 13024 18818 13028
rect 18834 13084 18898 13088
rect 18834 13028 18838 13084
rect 18838 13028 18894 13084
rect 18894 13028 18898 13084
rect 18834 13024 18898 13028
rect 18914 13084 18978 13088
rect 18914 13028 18918 13084
rect 18918 13028 18974 13084
rect 18974 13028 18978 13084
rect 18914 13024 18978 13028
rect 18994 13084 19058 13088
rect 18994 13028 18998 13084
rect 18998 13028 19054 13084
rect 19054 13028 19058 13084
rect 18994 13024 19058 13028
rect 24688 13084 24752 13088
rect 24688 13028 24692 13084
rect 24692 13028 24748 13084
rect 24748 13028 24752 13084
rect 24688 13024 24752 13028
rect 24768 13084 24832 13088
rect 24768 13028 24772 13084
rect 24772 13028 24828 13084
rect 24828 13028 24832 13084
rect 24768 13024 24832 13028
rect 24848 13084 24912 13088
rect 24848 13028 24852 13084
rect 24852 13028 24908 13084
rect 24908 13028 24912 13084
rect 24848 13024 24912 13028
rect 24928 13084 24992 13088
rect 24928 13028 24932 13084
rect 24932 13028 24988 13084
rect 24988 13028 24992 13084
rect 24928 13024 24992 13028
rect 3919 12540 3983 12544
rect 3919 12484 3923 12540
rect 3923 12484 3979 12540
rect 3979 12484 3983 12540
rect 3919 12480 3983 12484
rect 3999 12540 4063 12544
rect 3999 12484 4003 12540
rect 4003 12484 4059 12540
rect 4059 12484 4063 12540
rect 3999 12480 4063 12484
rect 4079 12540 4143 12544
rect 4079 12484 4083 12540
rect 4083 12484 4139 12540
rect 4139 12484 4143 12540
rect 4079 12480 4143 12484
rect 4159 12540 4223 12544
rect 4159 12484 4163 12540
rect 4163 12484 4219 12540
rect 4219 12484 4223 12540
rect 4159 12480 4223 12484
rect 10548 12684 10612 12748
rect 11652 12684 11716 12748
rect 9853 12540 9917 12544
rect 9853 12484 9857 12540
rect 9857 12484 9913 12540
rect 9913 12484 9917 12540
rect 9853 12480 9917 12484
rect 9933 12540 9997 12544
rect 9933 12484 9937 12540
rect 9937 12484 9993 12540
rect 9993 12484 9997 12540
rect 9933 12480 9997 12484
rect 10013 12540 10077 12544
rect 10013 12484 10017 12540
rect 10017 12484 10073 12540
rect 10073 12484 10077 12540
rect 10013 12480 10077 12484
rect 10093 12540 10157 12544
rect 10093 12484 10097 12540
rect 10097 12484 10153 12540
rect 10153 12484 10157 12540
rect 10093 12480 10157 12484
rect 15787 12540 15851 12544
rect 15787 12484 15791 12540
rect 15791 12484 15847 12540
rect 15847 12484 15851 12540
rect 15787 12480 15851 12484
rect 15867 12540 15931 12544
rect 15867 12484 15871 12540
rect 15871 12484 15927 12540
rect 15927 12484 15931 12540
rect 15867 12480 15931 12484
rect 15947 12540 16011 12544
rect 15947 12484 15951 12540
rect 15951 12484 16007 12540
rect 16007 12484 16011 12540
rect 15947 12480 16011 12484
rect 16027 12540 16091 12544
rect 16027 12484 16031 12540
rect 16031 12484 16087 12540
rect 16087 12484 16091 12540
rect 16027 12480 16091 12484
rect 21721 12540 21785 12544
rect 21721 12484 21725 12540
rect 21725 12484 21781 12540
rect 21781 12484 21785 12540
rect 21721 12480 21785 12484
rect 21801 12540 21865 12544
rect 21801 12484 21805 12540
rect 21805 12484 21861 12540
rect 21861 12484 21865 12540
rect 21801 12480 21865 12484
rect 21881 12540 21945 12544
rect 21881 12484 21885 12540
rect 21885 12484 21941 12540
rect 21941 12484 21945 12540
rect 21881 12480 21945 12484
rect 21961 12540 22025 12544
rect 21961 12484 21965 12540
rect 21965 12484 22021 12540
rect 22021 12484 22025 12540
rect 21961 12480 22025 12484
rect 21220 12336 21284 12340
rect 21220 12280 21234 12336
rect 21234 12280 21284 12336
rect 21220 12276 21284 12280
rect 3372 12140 3436 12204
rect 6886 11996 6950 12000
rect 6886 11940 6890 11996
rect 6890 11940 6946 11996
rect 6946 11940 6950 11996
rect 6886 11936 6950 11940
rect 6966 11996 7030 12000
rect 6966 11940 6970 11996
rect 6970 11940 7026 11996
rect 7026 11940 7030 11996
rect 6966 11936 7030 11940
rect 7046 11996 7110 12000
rect 7046 11940 7050 11996
rect 7050 11940 7106 11996
rect 7106 11940 7110 11996
rect 7046 11936 7110 11940
rect 7126 11996 7190 12000
rect 7126 11940 7130 11996
rect 7130 11940 7186 11996
rect 7186 11940 7190 11996
rect 7126 11936 7190 11940
rect 12820 11996 12884 12000
rect 12820 11940 12824 11996
rect 12824 11940 12880 11996
rect 12880 11940 12884 11996
rect 12820 11936 12884 11940
rect 12900 11996 12964 12000
rect 12900 11940 12904 11996
rect 12904 11940 12960 11996
rect 12960 11940 12964 11996
rect 12900 11936 12964 11940
rect 12980 11996 13044 12000
rect 12980 11940 12984 11996
rect 12984 11940 13040 11996
rect 13040 11940 13044 11996
rect 12980 11936 13044 11940
rect 13060 11996 13124 12000
rect 13060 11940 13064 11996
rect 13064 11940 13120 11996
rect 13120 11940 13124 11996
rect 13060 11936 13124 11940
rect 18754 11996 18818 12000
rect 18754 11940 18758 11996
rect 18758 11940 18814 11996
rect 18814 11940 18818 11996
rect 18754 11936 18818 11940
rect 18834 11996 18898 12000
rect 18834 11940 18838 11996
rect 18838 11940 18894 11996
rect 18894 11940 18898 11996
rect 18834 11936 18898 11940
rect 18914 11996 18978 12000
rect 18914 11940 18918 11996
rect 18918 11940 18974 11996
rect 18974 11940 18978 11996
rect 18914 11936 18978 11940
rect 18994 11996 19058 12000
rect 18994 11940 18998 11996
rect 18998 11940 19054 11996
rect 19054 11940 19058 11996
rect 18994 11936 19058 11940
rect 24688 11996 24752 12000
rect 24688 11940 24692 11996
rect 24692 11940 24748 11996
rect 24748 11940 24752 11996
rect 24688 11936 24752 11940
rect 24768 11996 24832 12000
rect 24768 11940 24772 11996
rect 24772 11940 24828 11996
rect 24828 11940 24832 11996
rect 24768 11936 24832 11940
rect 24848 11996 24912 12000
rect 24848 11940 24852 11996
rect 24852 11940 24908 11996
rect 24908 11940 24912 11996
rect 24848 11936 24912 11940
rect 24928 11996 24992 12000
rect 24928 11940 24932 11996
rect 24932 11940 24988 11996
rect 24988 11940 24992 11996
rect 24928 11936 24992 11940
rect 5028 11732 5092 11796
rect 3919 11452 3983 11456
rect 3919 11396 3923 11452
rect 3923 11396 3979 11452
rect 3979 11396 3983 11452
rect 3919 11392 3983 11396
rect 3999 11452 4063 11456
rect 3999 11396 4003 11452
rect 4003 11396 4059 11452
rect 4059 11396 4063 11452
rect 3999 11392 4063 11396
rect 4079 11452 4143 11456
rect 4079 11396 4083 11452
rect 4083 11396 4139 11452
rect 4139 11396 4143 11452
rect 4079 11392 4143 11396
rect 4159 11452 4223 11456
rect 4159 11396 4163 11452
rect 4163 11396 4219 11452
rect 4219 11396 4223 11452
rect 4159 11392 4223 11396
rect 9853 11452 9917 11456
rect 9853 11396 9857 11452
rect 9857 11396 9913 11452
rect 9913 11396 9917 11452
rect 9853 11392 9917 11396
rect 9933 11452 9997 11456
rect 9933 11396 9937 11452
rect 9937 11396 9993 11452
rect 9993 11396 9997 11452
rect 9933 11392 9997 11396
rect 10013 11452 10077 11456
rect 10013 11396 10017 11452
rect 10017 11396 10073 11452
rect 10073 11396 10077 11452
rect 10013 11392 10077 11396
rect 10093 11452 10157 11456
rect 10093 11396 10097 11452
rect 10097 11396 10153 11452
rect 10153 11396 10157 11452
rect 10093 11392 10157 11396
rect 15787 11452 15851 11456
rect 15787 11396 15791 11452
rect 15791 11396 15847 11452
rect 15847 11396 15851 11452
rect 15787 11392 15851 11396
rect 15867 11452 15931 11456
rect 15867 11396 15871 11452
rect 15871 11396 15927 11452
rect 15927 11396 15931 11452
rect 15867 11392 15931 11396
rect 15947 11452 16011 11456
rect 15947 11396 15951 11452
rect 15951 11396 16007 11452
rect 16007 11396 16011 11452
rect 15947 11392 16011 11396
rect 16027 11452 16091 11456
rect 16027 11396 16031 11452
rect 16031 11396 16087 11452
rect 16087 11396 16091 11452
rect 16027 11392 16091 11396
rect 21721 11452 21785 11456
rect 21721 11396 21725 11452
rect 21725 11396 21781 11452
rect 21781 11396 21785 11452
rect 21721 11392 21785 11396
rect 21801 11452 21865 11456
rect 21801 11396 21805 11452
rect 21805 11396 21861 11452
rect 21861 11396 21865 11452
rect 21801 11392 21865 11396
rect 21881 11452 21945 11456
rect 21881 11396 21885 11452
rect 21885 11396 21941 11452
rect 21941 11396 21945 11452
rect 21881 11392 21945 11396
rect 21961 11452 22025 11456
rect 21961 11396 21965 11452
rect 21965 11396 22021 11452
rect 22021 11396 22025 11452
rect 21961 11392 22025 11396
rect 20852 11324 20916 11388
rect 7420 11052 7484 11116
rect 10916 11052 10980 11116
rect 11836 11052 11900 11116
rect 19380 11052 19444 11116
rect 16252 10916 16316 10980
rect 6886 10908 6950 10912
rect 6886 10852 6890 10908
rect 6890 10852 6946 10908
rect 6946 10852 6950 10908
rect 6886 10848 6950 10852
rect 6966 10908 7030 10912
rect 6966 10852 6970 10908
rect 6970 10852 7026 10908
rect 7026 10852 7030 10908
rect 6966 10848 7030 10852
rect 7046 10908 7110 10912
rect 7046 10852 7050 10908
rect 7050 10852 7106 10908
rect 7106 10852 7110 10908
rect 7046 10848 7110 10852
rect 7126 10908 7190 10912
rect 7126 10852 7130 10908
rect 7130 10852 7186 10908
rect 7186 10852 7190 10908
rect 7126 10848 7190 10852
rect 12820 10908 12884 10912
rect 12820 10852 12824 10908
rect 12824 10852 12880 10908
rect 12880 10852 12884 10908
rect 12820 10848 12884 10852
rect 12900 10908 12964 10912
rect 12900 10852 12904 10908
rect 12904 10852 12960 10908
rect 12960 10852 12964 10908
rect 12900 10848 12964 10852
rect 12980 10908 13044 10912
rect 12980 10852 12984 10908
rect 12984 10852 13040 10908
rect 13040 10852 13044 10908
rect 12980 10848 13044 10852
rect 13060 10908 13124 10912
rect 13060 10852 13064 10908
rect 13064 10852 13120 10908
rect 13120 10852 13124 10908
rect 13060 10848 13124 10852
rect 18754 10908 18818 10912
rect 18754 10852 18758 10908
rect 18758 10852 18814 10908
rect 18814 10852 18818 10908
rect 18754 10848 18818 10852
rect 18834 10908 18898 10912
rect 18834 10852 18838 10908
rect 18838 10852 18894 10908
rect 18894 10852 18898 10908
rect 18834 10848 18898 10852
rect 18914 10908 18978 10912
rect 18914 10852 18918 10908
rect 18918 10852 18974 10908
rect 18974 10852 18978 10908
rect 18914 10848 18978 10852
rect 18994 10908 19058 10912
rect 18994 10852 18998 10908
rect 18998 10852 19054 10908
rect 19054 10852 19058 10908
rect 18994 10848 19058 10852
rect 24688 10908 24752 10912
rect 24688 10852 24692 10908
rect 24692 10852 24748 10908
rect 24748 10852 24752 10908
rect 24688 10848 24752 10852
rect 24768 10908 24832 10912
rect 24768 10852 24772 10908
rect 24772 10852 24828 10908
rect 24828 10852 24832 10908
rect 24768 10848 24832 10852
rect 24848 10908 24912 10912
rect 24848 10852 24852 10908
rect 24852 10852 24908 10908
rect 24908 10852 24912 10908
rect 24848 10848 24912 10852
rect 24928 10908 24992 10912
rect 24928 10852 24932 10908
rect 24932 10852 24988 10908
rect 24988 10852 24992 10908
rect 24928 10848 24992 10852
rect 15516 10840 15580 10844
rect 15516 10784 15530 10840
rect 15530 10784 15580 10840
rect 15516 10780 15580 10784
rect 11468 10644 11532 10708
rect 12572 10508 12636 10572
rect 3919 10364 3983 10368
rect 3919 10308 3923 10364
rect 3923 10308 3979 10364
rect 3979 10308 3983 10364
rect 3919 10304 3983 10308
rect 3999 10364 4063 10368
rect 3999 10308 4003 10364
rect 4003 10308 4059 10364
rect 4059 10308 4063 10364
rect 3999 10304 4063 10308
rect 4079 10364 4143 10368
rect 4079 10308 4083 10364
rect 4083 10308 4139 10364
rect 4139 10308 4143 10364
rect 4079 10304 4143 10308
rect 4159 10364 4223 10368
rect 4159 10308 4163 10364
rect 4163 10308 4219 10364
rect 4219 10308 4223 10364
rect 4159 10304 4223 10308
rect 9853 10364 9917 10368
rect 9853 10308 9857 10364
rect 9857 10308 9913 10364
rect 9913 10308 9917 10364
rect 9853 10304 9917 10308
rect 9933 10364 9997 10368
rect 9933 10308 9937 10364
rect 9937 10308 9993 10364
rect 9993 10308 9997 10364
rect 9933 10304 9997 10308
rect 10013 10364 10077 10368
rect 10013 10308 10017 10364
rect 10017 10308 10073 10364
rect 10073 10308 10077 10364
rect 10013 10304 10077 10308
rect 10093 10364 10157 10368
rect 10093 10308 10097 10364
rect 10097 10308 10153 10364
rect 10153 10308 10157 10364
rect 10093 10304 10157 10308
rect 15787 10364 15851 10368
rect 15787 10308 15791 10364
rect 15791 10308 15847 10364
rect 15847 10308 15851 10364
rect 15787 10304 15851 10308
rect 15867 10364 15931 10368
rect 15867 10308 15871 10364
rect 15871 10308 15927 10364
rect 15927 10308 15931 10364
rect 15867 10304 15931 10308
rect 15947 10364 16011 10368
rect 15947 10308 15951 10364
rect 15951 10308 16007 10364
rect 16007 10308 16011 10364
rect 15947 10304 16011 10308
rect 16027 10364 16091 10368
rect 16027 10308 16031 10364
rect 16031 10308 16087 10364
rect 16087 10308 16091 10364
rect 16027 10304 16091 10308
rect 21721 10364 21785 10368
rect 21721 10308 21725 10364
rect 21725 10308 21781 10364
rect 21781 10308 21785 10364
rect 21721 10304 21785 10308
rect 21801 10364 21865 10368
rect 21801 10308 21805 10364
rect 21805 10308 21861 10364
rect 21861 10308 21865 10364
rect 21801 10304 21865 10308
rect 21881 10364 21945 10368
rect 21881 10308 21885 10364
rect 21885 10308 21941 10364
rect 21941 10308 21945 10364
rect 21881 10304 21945 10308
rect 21961 10364 22025 10368
rect 21961 10308 21965 10364
rect 21965 10308 22021 10364
rect 22021 10308 22025 10364
rect 21961 10304 22025 10308
rect 1900 9964 1964 10028
rect 6316 9964 6380 10028
rect 20300 9828 20364 9892
rect 6886 9820 6950 9824
rect 6886 9764 6890 9820
rect 6890 9764 6946 9820
rect 6946 9764 6950 9820
rect 6886 9760 6950 9764
rect 6966 9820 7030 9824
rect 6966 9764 6970 9820
rect 6970 9764 7026 9820
rect 7026 9764 7030 9820
rect 6966 9760 7030 9764
rect 7046 9820 7110 9824
rect 7046 9764 7050 9820
rect 7050 9764 7106 9820
rect 7106 9764 7110 9820
rect 7046 9760 7110 9764
rect 7126 9820 7190 9824
rect 7126 9764 7130 9820
rect 7130 9764 7186 9820
rect 7186 9764 7190 9820
rect 7126 9760 7190 9764
rect 12820 9820 12884 9824
rect 12820 9764 12824 9820
rect 12824 9764 12880 9820
rect 12880 9764 12884 9820
rect 12820 9760 12884 9764
rect 12900 9820 12964 9824
rect 12900 9764 12904 9820
rect 12904 9764 12960 9820
rect 12960 9764 12964 9820
rect 12900 9760 12964 9764
rect 12980 9820 13044 9824
rect 12980 9764 12984 9820
rect 12984 9764 13040 9820
rect 13040 9764 13044 9820
rect 12980 9760 13044 9764
rect 13060 9820 13124 9824
rect 13060 9764 13064 9820
rect 13064 9764 13120 9820
rect 13120 9764 13124 9820
rect 13060 9760 13124 9764
rect 18754 9820 18818 9824
rect 18754 9764 18758 9820
rect 18758 9764 18814 9820
rect 18814 9764 18818 9820
rect 18754 9760 18818 9764
rect 18834 9820 18898 9824
rect 18834 9764 18838 9820
rect 18838 9764 18894 9820
rect 18894 9764 18898 9820
rect 18834 9760 18898 9764
rect 18914 9820 18978 9824
rect 18914 9764 18918 9820
rect 18918 9764 18974 9820
rect 18974 9764 18978 9820
rect 18914 9760 18978 9764
rect 18994 9820 19058 9824
rect 18994 9764 18998 9820
rect 18998 9764 19054 9820
rect 19054 9764 19058 9820
rect 18994 9760 19058 9764
rect 24688 9820 24752 9824
rect 24688 9764 24692 9820
rect 24692 9764 24748 9820
rect 24748 9764 24752 9820
rect 24688 9760 24752 9764
rect 24768 9820 24832 9824
rect 24768 9764 24772 9820
rect 24772 9764 24828 9820
rect 24828 9764 24832 9820
rect 24768 9760 24832 9764
rect 24848 9820 24912 9824
rect 24848 9764 24852 9820
rect 24852 9764 24908 9820
rect 24908 9764 24912 9820
rect 24848 9760 24912 9764
rect 24928 9820 24992 9824
rect 24928 9764 24932 9820
rect 24932 9764 24988 9820
rect 24988 9764 24992 9820
rect 24928 9760 24992 9764
rect 12204 9752 12268 9756
rect 12204 9696 12254 9752
rect 12254 9696 12268 9752
rect 12204 9692 12268 9696
rect 16252 9752 16316 9756
rect 16252 9696 16266 9752
rect 16266 9696 16316 9752
rect 16252 9692 16316 9696
rect 3004 9556 3068 9620
rect 3919 9276 3983 9280
rect 3919 9220 3923 9276
rect 3923 9220 3979 9276
rect 3979 9220 3983 9276
rect 3919 9216 3983 9220
rect 3999 9276 4063 9280
rect 3999 9220 4003 9276
rect 4003 9220 4059 9276
rect 4059 9220 4063 9276
rect 3999 9216 4063 9220
rect 4079 9276 4143 9280
rect 4079 9220 4083 9276
rect 4083 9220 4139 9276
rect 4139 9220 4143 9276
rect 4079 9216 4143 9220
rect 4159 9276 4223 9280
rect 4159 9220 4163 9276
rect 4163 9220 4219 9276
rect 4219 9220 4223 9276
rect 4159 9216 4223 9220
rect 9853 9276 9917 9280
rect 9853 9220 9857 9276
rect 9857 9220 9913 9276
rect 9913 9220 9917 9276
rect 9853 9216 9917 9220
rect 9933 9276 9997 9280
rect 9933 9220 9937 9276
rect 9937 9220 9993 9276
rect 9993 9220 9997 9276
rect 9933 9216 9997 9220
rect 10013 9276 10077 9280
rect 10013 9220 10017 9276
rect 10017 9220 10073 9276
rect 10073 9220 10077 9276
rect 10013 9216 10077 9220
rect 10093 9276 10157 9280
rect 10093 9220 10097 9276
rect 10097 9220 10153 9276
rect 10153 9220 10157 9276
rect 10093 9216 10157 9220
rect 15787 9276 15851 9280
rect 15787 9220 15791 9276
rect 15791 9220 15847 9276
rect 15847 9220 15851 9276
rect 15787 9216 15851 9220
rect 15867 9276 15931 9280
rect 15867 9220 15871 9276
rect 15871 9220 15927 9276
rect 15927 9220 15931 9276
rect 15867 9216 15931 9220
rect 15947 9276 16011 9280
rect 15947 9220 15951 9276
rect 15951 9220 16007 9276
rect 16007 9220 16011 9276
rect 15947 9216 16011 9220
rect 16027 9276 16091 9280
rect 16027 9220 16031 9276
rect 16031 9220 16087 9276
rect 16087 9220 16091 9276
rect 16027 9216 16091 9220
rect 21721 9276 21785 9280
rect 21721 9220 21725 9276
rect 21725 9220 21781 9276
rect 21781 9220 21785 9276
rect 21721 9216 21785 9220
rect 21801 9276 21865 9280
rect 21801 9220 21805 9276
rect 21805 9220 21861 9276
rect 21861 9220 21865 9276
rect 21801 9216 21865 9220
rect 21881 9276 21945 9280
rect 21881 9220 21885 9276
rect 21885 9220 21941 9276
rect 21941 9220 21945 9276
rect 21881 9216 21945 9220
rect 21961 9276 22025 9280
rect 21961 9220 21965 9276
rect 21965 9220 22021 9276
rect 22021 9220 22025 9276
rect 21961 9216 22025 9220
rect 6886 8732 6950 8736
rect 6886 8676 6890 8732
rect 6890 8676 6946 8732
rect 6946 8676 6950 8732
rect 6886 8672 6950 8676
rect 6966 8732 7030 8736
rect 6966 8676 6970 8732
rect 6970 8676 7026 8732
rect 7026 8676 7030 8732
rect 6966 8672 7030 8676
rect 7046 8732 7110 8736
rect 7046 8676 7050 8732
rect 7050 8676 7106 8732
rect 7106 8676 7110 8732
rect 7046 8672 7110 8676
rect 7126 8732 7190 8736
rect 7126 8676 7130 8732
rect 7130 8676 7186 8732
rect 7186 8676 7190 8732
rect 7126 8672 7190 8676
rect 12820 8732 12884 8736
rect 12820 8676 12824 8732
rect 12824 8676 12880 8732
rect 12880 8676 12884 8732
rect 12820 8672 12884 8676
rect 12900 8732 12964 8736
rect 12900 8676 12904 8732
rect 12904 8676 12960 8732
rect 12960 8676 12964 8732
rect 12900 8672 12964 8676
rect 12980 8732 13044 8736
rect 12980 8676 12984 8732
rect 12984 8676 13040 8732
rect 13040 8676 13044 8732
rect 12980 8672 13044 8676
rect 13060 8732 13124 8736
rect 13060 8676 13064 8732
rect 13064 8676 13120 8732
rect 13120 8676 13124 8732
rect 13060 8672 13124 8676
rect 18754 8732 18818 8736
rect 18754 8676 18758 8732
rect 18758 8676 18814 8732
rect 18814 8676 18818 8732
rect 18754 8672 18818 8676
rect 18834 8732 18898 8736
rect 18834 8676 18838 8732
rect 18838 8676 18894 8732
rect 18894 8676 18898 8732
rect 18834 8672 18898 8676
rect 18914 8732 18978 8736
rect 18914 8676 18918 8732
rect 18918 8676 18974 8732
rect 18974 8676 18978 8732
rect 18914 8672 18978 8676
rect 18994 8732 19058 8736
rect 18994 8676 18998 8732
rect 18998 8676 19054 8732
rect 19054 8676 19058 8732
rect 18994 8672 19058 8676
rect 24688 8732 24752 8736
rect 24688 8676 24692 8732
rect 24692 8676 24748 8732
rect 24748 8676 24752 8732
rect 24688 8672 24752 8676
rect 24768 8732 24832 8736
rect 24768 8676 24772 8732
rect 24772 8676 24828 8732
rect 24828 8676 24832 8732
rect 24768 8672 24832 8676
rect 24848 8732 24912 8736
rect 24848 8676 24852 8732
rect 24852 8676 24908 8732
rect 24908 8676 24912 8732
rect 24848 8672 24912 8676
rect 24928 8732 24992 8736
rect 24928 8676 24932 8732
rect 24932 8676 24988 8732
rect 24988 8676 24992 8732
rect 24928 8672 24992 8676
rect 13860 8196 13924 8260
rect 3919 8188 3983 8192
rect 3919 8132 3923 8188
rect 3923 8132 3979 8188
rect 3979 8132 3983 8188
rect 3919 8128 3983 8132
rect 3999 8188 4063 8192
rect 3999 8132 4003 8188
rect 4003 8132 4059 8188
rect 4059 8132 4063 8188
rect 3999 8128 4063 8132
rect 4079 8188 4143 8192
rect 4079 8132 4083 8188
rect 4083 8132 4139 8188
rect 4139 8132 4143 8188
rect 4079 8128 4143 8132
rect 4159 8188 4223 8192
rect 4159 8132 4163 8188
rect 4163 8132 4219 8188
rect 4219 8132 4223 8188
rect 4159 8128 4223 8132
rect 9853 8188 9917 8192
rect 9853 8132 9857 8188
rect 9857 8132 9913 8188
rect 9913 8132 9917 8188
rect 9853 8128 9917 8132
rect 9933 8188 9997 8192
rect 9933 8132 9937 8188
rect 9937 8132 9993 8188
rect 9993 8132 9997 8188
rect 9933 8128 9997 8132
rect 10013 8188 10077 8192
rect 10013 8132 10017 8188
rect 10017 8132 10073 8188
rect 10073 8132 10077 8188
rect 10013 8128 10077 8132
rect 10093 8188 10157 8192
rect 10093 8132 10097 8188
rect 10097 8132 10153 8188
rect 10153 8132 10157 8188
rect 10093 8128 10157 8132
rect 15787 8188 15851 8192
rect 15787 8132 15791 8188
rect 15791 8132 15847 8188
rect 15847 8132 15851 8188
rect 15787 8128 15851 8132
rect 15867 8188 15931 8192
rect 15867 8132 15871 8188
rect 15871 8132 15927 8188
rect 15927 8132 15931 8188
rect 15867 8128 15931 8132
rect 15947 8188 16011 8192
rect 15947 8132 15951 8188
rect 15951 8132 16007 8188
rect 16007 8132 16011 8188
rect 15947 8128 16011 8132
rect 16027 8188 16091 8192
rect 16027 8132 16031 8188
rect 16031 8132 16087 8188
rect 16087 8132 16091 8188
rect 16027 8128 16091 8132
rect 21721 8188 21785 8192
rect 21721 8132 21725 8188
rect 21725 8132 21781 8188
rect 21781 8132 21785 8188
rect 21721 8128 21785 8132
rect 21801 8188 21865 8192
rect 21801 8132 21805 8188
rect 21805 8132 21861 8188
rect 21861 8132 21865 8188
rect 21801 8128 21865 8132
rect 21881 8188 21945 8192
rect 21881 8132 21885 8188
rect 21885 8132 21941 8188
rect 21941 8132 21945 8188
rect 21881 8128 21945 8132
rect 21961 8188 22025 8192
rect 21961 8132 21965 8188
rect 21965 8132 22021 8188
rect 22021 8132 22025 8188
rect 21961 8128 22025 8132
rect 6886 7644 6950 7648
rect 6886 7588 6890 7644
rect 6890 7588 6946 7644
rect 6946 7588 6950 7644
rect 6886 7584 6950 7588
rect 6966 7644 7030 7648
rect 6966 7588 6970 7644
rect 6970 7588 7026 7644
rect 7026 7588 7030 7644
rect 6966 7584 7030 7588
rect 7046 7644 7110 7648
rect 7046 7588 7050 7644
rect 7050 7588 7106 7644
rect 7106 7588 7110 7644
rect 7046 7584 7110 7588
rect 7126 7644 7190 7648
rect 7126 7588 7130 7644
rect 7130 7588 7186 7644
rect 7186 7588 7190 7644
rect 7126 7584 7190 7588
rect 12820 7644 12884 7648
rect 12820 7588 12824 7644
rect 12824 7588 12880 7644
rect 12880 7588 12884 7644
rect 12820 7584 12884 7588
rect 12900 7644 12964 7648
rect 12900 7588 12904 7644
rect 12904 7588 12960 7644
rect 12960 7588 12964 7644
rect 12900 7584 12964 7588
rect 12980 7644 13044 7648
rect 12980 7588 12984 7644
rect 12984 7588 13040 7644
rect 13040 7588 13044 7644
rect 12980 7584 13044 7588
rect 13060 7644 13124 7648
rect 13060 7588 13064 7644
rect 13064 7588 13120 7644
rect 13120 7588 13124 7644
rect 13060 7584 13124 7588
rect 18754 7644 18818 7648
rect 18754 7588 18758 7644
rect 18758 7588 18814 7644
rect 18814 7588 18818 7644
rect 18754 7584 18818 7588
rect 18834 7644 18898 7648
rect 18834 7588 18838 7644
rect 18838 7588 18894 7644
rect 18894 7588 18898 7644
rect 18834 7584 18898 7588
rect 18914 7644 18978 7648
rect 18914 7588 18918 7644
rect 18918 7588 18974 7644
rect 18974 7588 18978 7644
rect 18914 7584 18978 7588
rect 18994 7644 19058 7648
rect 18994 7588 18998 7644
rect 18998 7588 19054 7644
rect 19054 7588 19058 7644
rect 18994 7584 19058 7588
rect 24688 7644 24752 7648
rect 24688 7588 24692 7644
rect 24692 7588 24748 7644
rect 24748 7588 24752 7644
rect 24688 7584 24752 7588
rect 24768 7644 24832 7648
rect 24768 7588 24772 7644
rect 24772 7588 24828 7644
rect 24828 7588 24832 7644
rect 24768 7584 24832 7588
rect 24848 7644 24912 7648
rect 24848 7588 24852 7644
rect 24852 7588 24908 7644
rect 24908 7588 24912 7644
rect 24848 7584 24912 7588
rect 24928 7644 24992 7648
rect 24928 7588 24932 7644
rect 24932 7588 24988 7644
rect 24988 7588 24992 7644
rect 24928 7584 24992 7588
rect 17908 7516 17972 7580
rect 14964 7244 15028 7308
rect 3919 7100 3983 7104
rect 3919 7044 3923 7100
rect 3923 7044 3979 7100
rect 3979 7044 3983 7100
rect 3919 7040 3983 7044
rect 3999 7100 4063 7104
rect 3999 7044 4003 7100
rect 4003 7044 4059 7100
rect 4059 7044 4063 7100
rect 3999 7040 4063 7044
rect 4079 7100 4143 7104
rect 4079 7044 4083 7100
rect 4083 7044 4139 7100
rect 4139 7044 4143 7100
rect 4079 7040 4143 7044
rect 4159 7100 4223 7104
rect 4159 7044 4163 7100
rect 4163 7044 4219 7100
rect 4219 7044 4223 7100
rect 4159 7040 4223 7044
rect 9853 7100 9917 7104
rect 9853 7044 9857 7100
rect 9857 7044 9913 7100
rect 9913 7044 9917 7100
rect 9853 7040 9917 7044
rect 9933 7100 9997 7104
rect 9933 7044 9937 7100
rect 9937 7044 9993 7100
rect 9993 7044 9997 7100
rect 9933 7040 9997 7044
rect 10013 7100 10077 7104
rect 10013 7044 10017 7100
rect 10017 7044 10073 7100
rect 10073 7044 10077 7100
rect 10013 7040 10077 7044
rect 10093 7100 10157 7104
rect 10093 7044 10097 7100
rect 10097 7044 10153 7100
rect 10153 7044 10157 7100
rect 10093 7040 10157 7044
rect 15787 7100 15851 7104
rect 15787 7044 15791 7100
rect 15791 7044 15847 7100
rect 15847 7044 15851 7100
rect 15787 7040 15851 7044
rect 15867 7100 15931 7104
rect 15867 7044 15871 7100
rect 15871 7044 15927 7100
rect 15927 7044 15931 7100
rect 15867 7040 15931 7044
rect 15947 7100 16011 7104
rect 15947 7044 15951 7100
rect 15951 7044 16007 7100
rect 16007 7044 16011 7100
rect 15947 7040 16011 7044
rect 16027 7100 16091 7104
rect 16027 7044 16031 7100
rect 16031 7044 16087 7100
rect 16087 7044 16091 7100
rect 16027 7040 16091 7044
rect 21721 7100 21785 7104
rect 21721 7044 21725 7100
rect 21725 7044 21781 7100
rect 21781 7044 21785 7100
rect 21721 7040 21785 7044
rect 21801 7100 21865 7104
rect 21801 7044 21805 7100
rect 21805 7044 21861 7100
rect 21861 7044 21865 7100
rect 21801 7040 21865 7044
rect 21881 7100 21945 7104
rect 21881 7044 21885 7100
rect 21885 7044 21941 7100
rect 21941 7044 21945 7100
rect 21881 7040 21945 7044
rect 21961 7100 22025 7104
rect 21961 7044 21965 7100
rect 21965 7044 22021 7100
rect 22021 7044 22025 7100
rect 21961 7040 22025 7044
rect 4660 6836 4724 6900
rect 22140 6700 22204 6764
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 21404 6216 21468 6220
rect 21404 6160 21418 6216
rect 21418 6160 21468 6216
rect 21404 6156 21468 6160
rect 10548 6020 10612 6084
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 3556 5748 3620 5812
rect 11652 5884 11716 5948
rect 22692 5536 22756 5540
rect 22692 5480 22742 5536
rect 22742 5480 22756 5536
rect 22692 5476 22756 5480
rect 22876 5476 22940 5540
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 16988 5068 17052 5132
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 980 3980 1044 4044
rect 12204 4040 12268 4044
rect 12204 3984 12254 4040
rect 12254 3984 12268 4040
rect 12204 3980 12268 3984
rect 14596 3980 14660 4044
rect 18276 4040 18340 4044
rect 18276 3984 18326 4040
rect 18326 3984 18340 4040
rect 18276 3980 18340 3984
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 17540 3708 17604 3772
rect 19196 3768 19260 3772
rect 19196 3712 19210 3768
rect 19210 3712 19260 3768
rect 19196 3708 19260 3712
rect 796 3300 860 3364
rect 10916 3300 10980 3364
rect 12572 3360 12636 3364
rect 12572 3304 12622 3360
rect 12622 3304 12636 3360
rect 12572 3300 12636 3304
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 22140 3164 22204 3228
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 2084 2680 2148 2684
rect 2084 2624 2134 2680
rect 2134 2624 2148 2680
rect 2084 2620 2148 2624
rect 9444 2680 9508 2684
rect 9444 2624 9494 2680
rect 9494 2624 9508 2680
rect 9444 2620 9508 2624
rect 13308 2620 13372 2684
rect 17356 2620 17420 2684
rect 18460 2680 18524 2684
rect 18460 2624 18510 2680
rect 18510 2624 18524 2680
rect 18460 2620 18524 2624
rect 19196 2620 19260 2684
rect 19564 2620 19628 2684
rect 19932 2620 19996 2684
rect 2636 2484 2700 2548
rect 1164 2348 1228 2412
rect 10548 2348 10612 2412
rect 12020 2348 12084 2412
rect 17724 2348 17788 2412
rect 7788 2272 7852 2276
rect 7788 2216 7802 2272
rect 7802 2216 7852 2272
rect 7788 2212 7852 2216
rect 8156 2272 8220 2276
rect 8156 2216 8170 2272
rect 8170 2216 8220 2272
rect 8156 2212 8220 2216
rect 8524 2212 8588 2276
rect 8892 2272 8956 2276
rect 8892 2216 8906 2272
rect 8906 2216 8956 2272
rect 8892 2212 8956 2216
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 20668 1940 20732 2004
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 4844 1260 4908 1324
rect 5580 1320 5644 1324
rect 5580 1264 5594 1320
rect 5594 1264 5644 1320
rect 5580 1260 5644 1264
rect 6500 1320 6564 1324
rect 6500 1264 6550 1320
rect 6550 1264 6564 1320
rect 6500 1260 6564 1264
rect 7972 1320 8036 1324
rect 7972 1264 7986 1320
rect 7986 1264 8036 1320
rect 7972 1260 8036 1264
rect 8708 1320 8772 1324
rect 8708 1264 8722 1320
rect 8722 1264 8772 1320
rect 8708 1260 8772 1264
rect 16436 1320 16500 1324
rect 16436 1264 16486 1320
rect 16486 1264 16500 1320
rect 16436 1260 16500 1264
rect 612 1124 676 1188
rect 6132 1124 6196 1188
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
<< metal4 >>
rect 3911 43008 4231 43568
rect 3911 42944 3919 43008
rect 3983 42944 3999 43008
rect 4063 42944 4079 43008
rect 4143 42944 4159 43008
rect 4223 42944 4231 43008
rect 3911 41920 4231 42944
rect 3911 41856 3919 41920
rect 3983 41856 3999 41920
rect 4063 41856 4079 41920
rect 4143 41856 4159 41920
rect 4223 41856 4231 41920
rect 1163 41716 1229 41717
rect 1163 41652 1164 41716
rect 1228 41652 1229 41716
rect 1163 41651 1229 41652
rect 795 41580 861 41581
rect 795 41516 796 41580
rect 860 41516 861 41580
rect 795 41515 861 41516
rect 611 28252 677 28253
rect 611 28188 612 28252
rect 676 28188 677 28252
rect 611 28187 677 28188
rect 614 1189 674 28187
rect 798 3365 858 41515
rect 979 41444 1045 41445
rect 979 41380 980 41444
rect 1044 41380 1045 41444
rect 979 41379 1045 41380
rect 982 4045 1042 41379
rect 979 4044 1045 4045
rect 979 3980 980 4044
rect 1044 3980 1045 4044
rect 979 3979 1045 3980
rect 795 3364 861 3365
rect 795 3300 796 3364
rect 860 3300 861 3364
rect 795 3299 861 3300
rect 1166 2413 1226 41651
rect 3911 40832 4231 41856
rect 6878 43552 7198 43568
rect 6878 43488 6886 43552
rect 6950 43488 6966 43552
rect 7030 43488 7046 43552
rect 7110 43488 7126 43552
rect 7190 43488 7198 43552
rect 6878 42464 7198 43488
rect 6878 42400 6886 42464
rect 6950 42400 6966 42464
rect 7030 42400 7046 42464
rect 7110 42400 7126 42464
rect 7190 42400 7198 42464
rect 6315 41852 6381 41853
rect 6315 41788 6316 41852
rect 6380 41788 6381 41852
rect 6315 41787 6381 41788
rect 4659 41580 4725 41581
rect 4659 41516 4660 41580
rect 4724 41516 4725 41580
rect 4659 41515 4725 41516
rect 6131 41580 6197 41581
rect 6131 41516 6132 41580
rect 6196 41516 6197 41580
rect 6131 41515 6197 41516
rect 3911 40768 3919 40832
rect 3983 40768 3999 40832
rect 4063 40768 4079 40832
rect 4143 40768 4159 40832
rect 4223 40768 4231 40832
rect 3911 39744 4231 40768
rect 3911 39680 3919 39744
rect 3983 39680 3999 39744
rect 4063 39680 4079 39744
rect 4143 39680 4159 39744
rect 4223 39680 4231 39744
rect 2635 39132 2701 39133
rect 2635 39068 2636 39132
rect 2700 39068 2701 39132
rect 2635 39067 2701 39068
rect 2451 36140 2517 36141
rect 2451 36076 2452 36140
rect 2516 36076 2517 36140
rect 2451 36075 2517 36076
rect 2083 34644 2149 34645
rect 2083 34580 2084 34644
rect 2148 34580 2149 34644
rect 2083 34579 2149 34580
rect 2086 30970 2146 34579
rect 2454 33421 2514 36075
rect 2451 33420 2517 33421
rect 2451 33356 2452 33420
rect 2516 33356 2517 33420
rect 2451 33355 2517 33356
rect 2086 30910 2330 30970
rect 2270 30701 2330 30910
rect 2267 30700 2333 30701
rect 2267 30636 2268 30700
rect 2332 30636 2333 30700
rect 2267 30635 2333 30636
rect 2083 29068 2149 29069
rect 2083 29004 2084 29068
rect 2148 29004 2149 29068
rect 2083 29003 2149 29004
rect 1899 28660 1965 28661
rect 1899 28596 1900 28660
rect 1964 28596 1965 28660
rect 1899 28595 1965 28596
rect 1715 28388 1781 28389
rect 1715 28324 1716 28388
rect 1780 28324 1781 28388
rect 1715 28323 1781 28324
rect 1347 26892 1413 26893
rect 1347 26828 1348 26892
rect 1412 26828 1413 26892
rect 1347 26827 1413 26828
rect 1350 20909 1410 26827
rect 1718 23493 1778 28323
rect 1715 23492 1781 23493
rect 1715 23428 1716 23492
rect 1780 23428 1781 23492
rect 1715 23427 1781 23428
rect 1902 21997 1962 28595
rect 2086 26893 2146 29003
rect 2083 26892 2149 26893
rect 2083 26828 2084 26892
rect 2148 26828 2149 26892
rect 2083 26827 2149 26828
rect 2270 26077 2330 30635
rect 2638 28930 2698 39067
rect 3911 38656 4231 39680
rect 3911 38592 3919 38656
rect 3983 38592 3999 38656
rect 4063 38592 4079 38656
rect 4143 38592 4159 38656
rect 4223 38592 4231 38656
rect 2819 38180 2885 38181
rect 2819 38116 2820 38180
rect 2884 38116 2885 38180
rect 2819 38115 2885 38116
rect 2822 29749 2882 38115
rect 3911 37568 4231 38592
rect 3911 37504 3919 37568
rect 3983 37504 3999 37568
rect 4063 37504 4079 37568
rect 4143 37504 4159 37568
rect 4223 37504 4231 37568
rect 3003 37500 3069 37501
rect 3003 37436 3004 37500
rect 3068 37436 3069 37500
rect 3003 37435 3069 37436
rect 3006 36141 3066 37435
rect 3911 36480 4231 37504
rect 3911 36416 3919 36480
rect 3983 36416 3999 36480
rect 4063 36416 4079 36480
rect 4143 36416 4159 36480
rect 4223 36416 4231 36480
rect 3003 36140 3069 36141
rect 3003 36076 3004 36140
rect 3068 36076 3069 36140
rect 3003 36075 3069 36076
rect 3006 33829 3066 36075
rect 3739 36004 3805 36005
rect 3739 35940 3740 36004
rect 3804 35940 3805 36004
rect 3739 35939 3805 35940
rect 3003 33828 3069 33829
rect 3003 33764 3004 33828
rect 3068 33764 3069 33828
rect 3003 33763 3069 33764
rect 3742 33693 3802 35939
rect 3911 35392 4231 36416
rect 3911 35328 3919 35392
rect 3983 35328 3999 35392
rect 4063 35328 4079 35392
rect 4143 35328 4159 35392
rect 4223 35328 4231 35392
rect 3911 34304 4231 35328
rect 4475 34644 4541 34645
rect 4475 34580 4476 34644
rect 4540 34580 4541 34644
rect 4475 34579 4541 34580
rect 3911 34240 3919 34304
rect 3983 34240 3999 34304
rect 4063 34240 4079 34304
rect 4143 34240 4159 34304
rect 4223 34240 4231 34304
rect 3739 33692 3805 33693
rect 3739 33628 3740 33692
rect 3804 33628 3805 33692
rect 3739 33627 3805 33628
rect 3911 33216 4231 34240
rect 3911 33152 3919 33216
rect 3983 33152 3999 33216
rect 4063 33152 4079 33216
rect 4143 33152 4159 33216
rect 4223 33152 4231 33216
rect 3555 32332 3621 32333
rect 3555 32268 3556 32332
rect 3620 32268 3621 32332
rect 3555 32267 3621 32268
rect 3371 30428 3437 30429
rect 3371 30364 3372 30428
rect 3436 30364 3437 30428
rect 3371 30363 3437 30364
rect 2819 29748 2885 29749
rect 2819 29684 2820 29748
rect 2884 29684 2885 29748
rect 2819 29683 2885 29684
rect 2454 28870 2698 28930
rect 2454 26757 2514 28870
rect 2635 28524 2701 28525
rect 2635 28460 2636 28524
rect 2700 28460 2701 28524
rect 2635 28459 2701 28460
rect 2451 26756 2517 26757
rect 2451 26692 2452 26756
rect 2516 26692 2517 26756
rect 2451 26691 2517 26692
rect 2267 26076 2333 26077
rect 2267 26012 2268 26076
rect 2332 26012 2333 26076
rect 2267 26011 2333 26012
rect 2451 26076 2517 26077
rect 2451 26012 2452 26076
rect 2516 26012 2517 26076
rect 2451 26011 2517 26012
rect 2267 22676 2333 22677
rect 2267 22612 2268 22676
rect 2332 22612 2333 22676
rect 2267 22611 2333 22612
rect 1899 21996 1965 21997
rect 1899 21932 1900 21996
rect 1964 21932 1965 21996
rect 1899 21931 1965 21932
rect 1347 20908 1413 20909
rect 1347 20844 1348 20908
rect 1412 20844 1413 20908
rect 1347 20843 1413 20844
rect 2083 17372 2149 17373
rect 2083 17308 2084 17372
rect 2148 17308 2149 17372
rect 2083 17307 2149 17308
rect 1899 16828 1965 16829
rect 1899 16764 1900 16828
rect 1964 16764 1965 16828
rect 1899 16763 1965 16764
rect 1902 10029 1962 16763
rect 1899 10028 1965 10029
rect 1899 9964 1900 10028
rect 1964 9964 1965 10028
rect 1899 9963 1965 9964
rect 2086 2685 2146 17307
rect 2270 12450 2330 22611
rect 2454 18869 2514 26011
rect 2451 18868 2517 18869
rect 2451 18804 2452 18868
rect 2516 18804 2517 18868
rect 2451 18803 2517 18804
rect 2638 18461 2698 28459
rect 2822 23901 2882 29683
rect 3003 27436 3069 27437
rect 3003 27372 3004 27436
rect 3068 27372 3069 27436
rect 3003 27371 3069 27372
rect 3006 24309 3066 27371
rect 3003 24308 3069 24309
rect 3003 24244 3004 24308
rect 3068 24244 3069 24308
rect 3003 24243 3069 24244
rect 2819 23900 2885 23901
rect 2819 23836 2820 23900
rect 2884 23836 2885 23900
rect 2819 23835 2885 23836
rect 3006 20229 3066 24243
rect 3003 20228 3069 20229
rect 3003 20164 3004 20228
rect 3068 20164 3069 20228
rect 3003 20163 3069 20164
rect 2635 18460 2701 18461
rect 2635 18396 2636 18460
rect 2700 18396 2701 18460
rect 2635 18395 2701 18396
rect 2270 12390 2698 12450
rect 2083 2684 2149 2685
rect 2083 2620 2084 2684
rect 2148 2620 2149 2684
rect 2083 2619 2149 2620
rect 2638 2549 2698 12390
rect 3006 9621 3066 20163
rect 3374 15605 3434 30363
rect 3558 16285 3618 32267
rect 3911 32128 4231 33152
rect 3911 32064 3919 32128
rect 3983 32064 3999 32128
rect 4063 32064 4079 32128
rect 4143 32064 4159 32128
rect 4223 32064 4231 32128
rect 3911 31040 4231 32064
rect 3911 30976 3919 31040
rect 3983 30976 3999 31040
rect 4063 30976 4079 31040
rect 4143 30976 4159 31040
rect 4223 30976 4231 31040
rect 3911 29952 4231 30976
rect 4478 30293 4538 34579
rect 4662 34101 4722 41515
rect 5579 35188 5645 35189
rect 5579 35124 5580 35188
rect 5644 35124 5645 35188
rect 5579 35123 5645 35124
rect 5395 34508 5461 34509
rect 5395 34444 5396 34508
rect 5460 34444 5461 34508
rect 5395 34443 5461 34444
rect 4659 34100 4725 34101
rect 4659 34036 4660 34100
rect 4724 34036 4725 34100
rect 4659 34035 4725 34036
rect 4659 31380 4725 31381
rect 4659 31316 4660 31380
rect 4724 31316 4725 31380
rect 4659 31315 4725 31316
rect 4475 30292 4541 30293
rect 4475 30228 4476 30292
rect 4540 30228 4541 30292
rect 4475 30227 4541 30228
rect 3911 29888 3919 29952
rect 3983 29888 3999 29952
rect 4063 29888 4079 29952
rect 4143 29888 4159 29952
rect 4223 29888 4231 29952
rect 3911 28864 4231 29888
rect 3911 28800 3919 28864
rect 3983 28800 3999 28864
rect 4063 28800 4079 28864
rect 4143 28800 4159 28864
rect 4223 28800 4231 28864
rect 3911 27776 4231 28800
rect 3911 27712 3919 27776
rect 3983 27712 3999 27776
rect 4063 27712 4079 27776
rect 4143 27712 4159 27776
rect 4223 27712 4231 27776
rect 3911 26688 4231 27712
rect 3911 26624 3919 26688
rect 3983 26624 3999 26688
rect 4063 26624 4079 26688
rect 4143 26624 4159 26688
rect 4223 26624 4231 26688
rect 3911 25600 4231 26624
rect 3911 25536 3919 25600
rect 3983 25536 3999 25600
rect 4063 25536 4079 25600
rect 4143 25536 4159 25600
rect 4223 25536 4231 25600
rect 3911 24512 4231 25536
rect 3911 24448 3919 24512
rect 3983 24448 3999 24512
rect 4063 24448 4079 24512
rect 4143 24448 4159 24512
rect 4223 24448 4231 24512
rect 3911 23424 4231 24448
rect 3911 23360 3919 23424
rect 3983 23360 3999 23424
rect 4063 23360 4079 23424
rect 4143 23360 4159 23424
rect 4223 23360 4231 23424
rect 3911 22336 4231 23360
rect 3911 22272 3919 22336
rect 3983 22272 3999 22336
rect 4063 22272 4079 22336
rect 4143 22272 4159 22336
rect 4223 22272 4231 22336
rect 3911 21248 4231 22272
rect 3911 21184 3919 21248
rect 3983 21184 3999 21248
rect 4063 21184 4079 21248
rect 4143 21184 4159 21248
rect 4223 21184 4231 21248
rect 3911 20160 4231 21184
rect 4478 21045 4538 30227
rect 4662 25941 4722 31315
rect 4843 30428 4909 30429
rect 4843 30364 4844 30428
rect 4908 30364 4909 30428
rect 4843 30363 4909 30364
rect 4659 25940 4725 25941
rect 4659 25876 4660 25940
rect 4724 25876 4725 25940
rect 4659 25875 4725 25876
rect 4846 23493 4906 30363
rect 5398 29749 5458 34443
rect 5395 29748 5461 29749
rect 5395 29684 5396 29748
rect 5460 29684 5461 29748
rect 5395 29683 5461 29684
rect 5395 29068 5461 29069
rect 5395 29004 5396 29068
rect 5460 29010 5461 29068
rect 5582 29010 5642 35123
rect 5460 29004 5642 29010
rect 5395 29003 5642 29004
rect 5398 28950 5642 29003
rect 5027 28524 5093 28525
rect 5027 28460 5028 28524
rect 5092 28460 5093 28524
rect 5027 28459 5093 28460
rect 4843 23492 4909 23493
rect 4843 23428 4844 23492
rect 4908 23428 4909 23492
rect 4843 23427 4909 23428
rect 4659 22812 4725 22813
rect 4659 22748 4660 22812
rect 4724 22748 4725 22812
rect 4659 22747 4725 22748
rect 4475 21044 4541 21045
rect 4475 20980 4476 21044
rect 4540 20980 4541 21044
rect 4475 20979 4541 20980
rect 3911 20096 3919 20160
rect 3983 20096 3999 20160
rect 4063 20096 4079 20160
rect 4143 20096 4159 20160
rect 4223 20096 4231 20160
rect 3911 19072 4231 20096
rect 3911 19008 3919 19072
rect 3983 19008 3999 19072
rect 4063 19008 4079 19072
rect 4143 19008 4159 19072
rect 4223 19008 4231 19072
rect 3911 17984 4231 19008
rect 3911 17920 3919 17984
rect 3983 17920 3999 17984
rect 4063 17920 4079 17984
rect 4143 17920 4159 17984
rect 4223 17920 4231 17984
rect 3911 16896 4231 17920
rect 3911 16832 3919 16896
rect 3983 16832 3999 16896
rect 4063 16832 4079 16896
rect 4143 16832 4159 16896
rect 4223 16832 4231 16896
rect 3555 16284 3621 16285
rect 3555 16220 3556 16284
rect 3620 16220 3621 16284
rect 3555 16219 3621 16220
rect 3911 15808 4231 16832
rect 3911 15744 3919 15808
rect 3983 15744 3999 15808
rect 4063 15744 4079 15808
rect 4143 15744 4159 15808
rect 4223 15744 4231 15808
rect 3371 15604 3437 15605
rect 3371 15540 3372 15604
rect 3436 15540 3437 15604
rect 3371 15539 3437 15540
rect 3374 12205 3434 15539
rect 3911 14720 4231 15744
rect 4662 15197 4722 22747
rect 4843 18188 4909 18189
rect 4843 18124 4844 18188
rect 4908 18124 4909 18188
rect 4843 18123 4909 18124
rect 4659 15196 4725 15197
rect 4659 15132 4660 15196
rect 4724 15132 4725 15196
rect 4659 15131 4725 15132
rect 3911 14656 3919 14720
rect 3983 14656 3999 14720
rect 4063 14656 4079 14720
rect 4143 14656 4159 14720
rect 4223 14656 4231 14720
rect 3911 13632 4231 14656
rect 3911 13568 3919 13632
rect 3983 13568 3999 13632
rect 4063 13568 4079 13632
rect 4143 13568 4159 13632
rect 4223 13568 4231 13632
rect 3555 13292 3621 13293
rect 3555 13228 3556 13292
rect 3620 13228 3621 13292
rect 3555 13227 3621 13228
rect 3371 12204 3437 12205
rect 3371 12140 3372 12204
rect 3436 12140 3437 12204
rect 3371 12139 3437 12140
rect 3003 9620 3069 9621
rect 3003 9556 3004 9620
rect 3068 9556 3069 9620
rect 3003 9555 3069 9556
rect 3558 5813 3618 13227
rect 3911 12544 4231 13568
rect 3911 12480 3919 12544
rect 3983 12480 3999 12544
rect 4063 12480 4079 12544
rect 4143 12480 4159 12544
rect 4223 12480 4231 12544
rect 3911 11456 4231 12480
rect 3911 11392 3919 11456
rect 3983 11392 3999 11456
rect 4063 11392 4079 11456
rect 4143 11392 4159 11456
rect 4223 11392 4231 11456
rect 3911 10368 4231 11392
rect 3911 10304 3919 10368
rect 3983 10304 3999 10368
rect 4063 10304 4079 10368
rect 4143 10304 4159 10368
rect 4223 10304 4231 10368
rect 3911 9280 4231 10304
rect 3911 9216 3919 9280
rect 3983 9216 3999 9280
rect 4063 9216 4079 9280
rect 4143 9216 4159 9280
rect 4223 9216 4231 9280
rect 3911 8192 4231 9216
rect 3911 8128 3919 8192
rect 3983 8128 3999 8192
rect 4063 8128 4079 8192
rect 4143 8128 4159 8192
rect 4223 8128 4231 8192
rect 3911 7104 4231 8128
rect 3911 7040 3919 7104
rect 3983 7040 3999 7104
rect 4063 7040 4079 7104
rect 4143 7040 4159 7104
rect 4223 7040 4231 7104
rect 3911 6016 4231 7040
rect 4662 6901 4722 15131
rect 4659 6900 4725 6901
rect 4659 6836 4660 6900
rect 4724 6836 4725 6900
rect 4659 6835 4725 6836
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3555 5812 3621 5813
rect 3555 5748 3556 5812
rect 3620 5748 3621 5812
rect 3555 5747 3621 5748
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 2635 2548 2701 2549
rect 2635 2484 2636 2548
rect 2700 2484 2701 2548
rect 2635 2483 2701 2484
rect 1163 2412 1229 2413
rect 1163 2348 1164 2412
rect 1228 2348 1229 2412
rect 1163 2347 1229 2348
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 611 1188 677 1189
rect 611 1124 612 1188
rect 676 1124 677 1188
rect 611 1123 677 1124
rect 3911 1040 4231 1600
rect 4846 1325 4906 18123
rect 5030 11797 5090 28459
rect 5398 21997 5458 28950
rect 5947 27436 6013 27437
rect 5947 27372 5948 27436
rect 6012 27372 6013 27436
rect 5947 27371 6013 27372
rect 5579 24852 5645 24853
rect 5579 24788 5580 24852
rect 5644 24788 5645 24852
rect 5579 24787 5645 24788
rect 5395 21996 5461 21997
rect 5395 21932 5396 21996
rect 5460 21932 5461 21996
rect 5395 21931 5461 21932
rect 5398 20909 5458 21931
rect 5395 20908 5461 20909
rect 5395 20844 5396 20908
rect 5460 20844 5461 20908
rect 5395 20843 5461 20844
rect 5395 18460 5461 18461
rect 5395 18396 5396 18460
rect 5460 18396 5461 18460
rect 5395 18395 5461 18396
rect 5398 13973 5458 18395
rect 5395 13972 5461 13973
rect 5395 13908 5396 13972
rect 5460 13908 5461 13972
rect 5395 13907 5461 13908
rect 5027 11796 5093 11797
rect 5027 11732 5028 11796
rect 5092 11732 5093 11796
rect 5027 11731 5093 11732
rect 5582 1325 5642 24787
rect 5950 23493 6010 27371
rect 6134 26213 6194 41515
rect 6131 26212 6197 26213
rect 6131 26148 6132 26212
rect 6196 26148 6197 26212
rect 6131 26147 6197 26148
rect 6131 25668 6197 25669
rect 6131 25604 6132 25668
rect 6196 25604 6197 25668
rect 6131 25603 6197 25604
rect 5947 23492 6013 23493
rect 5947 23428 5948 23492
rect 6012 23428 6013 23492
rect 5947 23427 6013 23428
rect 6134 21861 6194 25603
rect 6131 21860 6197 21861
rect 6131 21796 6132 21860
rect 6196 21796 6197 21860
rect 6131 21795 6197 21796
rect 5947 14788 6013 14789
rect 5947 14724 5948 14788
rect 6012 14724 6013 14788
rect 5947 14723 6013 14724
rect 5950 13565 6010 14723
rect 6131 14652 6197 14653
rect 6131 14588 6132 14652
rect 6196 14588 6197 14652
rect 6131 14587 6197 14588
rect 5947 13564 6013 13565
rect 5947 13500 5948 13564
rect 6012 13500 6013 13564
rect 5947 13499 6013 13500
rect 4843 1324 4909 1325
rect 4843 1260 4844 1324
rect 4908 1260 4909 1324
rect 4843 1259 4909 1260
rect 5579 1324 5645 1325
rect 5579 1260 5580 1324
rect 5644 1260 5645 1324
rect 5579 1259 5645 1260
rect 6134 1189 6194 14587
rect 6318 10029 6378 41787
rect 6878 41376 7198 42400
rect 9845 43008 10165 43568
rect 9845 42944 9853 43008
rect 9917 42944 9933 43008
rect 9997 42944 10013 43008
rect 10077 42944 10093 43008
rect 10157 42944 10165 43008
rect 7603 42260 7669 42261
rect 7603 42196 7604 42260
rect 7668 42196 7669 42260
rect 7603 42195 7669 42196
rect 6878 41312 6886 41376
rect 6950 41312 6966 41376
rect 7030 41312 7046 41376
rect 7110 41312 7126 41376
rect 7190 41312 7198 41376
rect 6878 40288 7198 41312
rect 6878 40224 6886 40288
rect 6950 40224 6966 40288
rect 7030 40224 7046 40288
rect 7110 40224 7126 40288
rect 7190 40224 7198 40288
rect 6878 39200 7198 40224
rect 6878 39136 6886 39200
rect 6950 39136 6966 39200
rect 7030 39136 7046 39200
rect 7110 39136 7126 39200
rect 7190 39136 7198 39200
rect 6878 38112 7198 39136
rect 6878 38048 6886 38112
rect 6950 38048 6966 38112
rect 7030 38048 7046 38112
rect 7110 38048 7126 38112
rect 7190 38048 7198 38112
rect 6683 37364 6749 37365
rect 6683 37300 6684 37364
rect 6748 37300 6749 37364
rect 6683 37299 6749 37300
rect 6686 35461 6746 37299
rect 6878 37024 7198 38048
rect 6878 36960 6886 37024
rect 6950 36960 6966 37024
rect 7030 36960 7046 37024
rect 7110 36960 7126 37024
rect 7190 36960 7198 37024
rect 6878 35936 7198 36960
rect 6878 35872 6886 35936
rect 6950 35872 6966 35936
rect 7030 35872 7046 35936
rect 7110 35872 7126 35936
rect 7190 35872 7198 35936
rect 6683 35460 6749 35461
rect 6683 35396 6684 35460
rect 6748 35396 6749 35460
rect 6683 35395 6749 35396
rect 6499 25940 6565 25941
rect 6499 25876 6500 25940
rect 6564 25876 6565 25940
rect 6499 25875 6565 25876
rect 6502 23493 6562 25875
rect 6499 23492 6565 23493
rect 6499 23428 6500 23492
rect 6564 23428 6565 23492
rect 6499 23427 6565 23428
rect 6686 22110 6746 35395
rect 6502 22050 6746 22110
rect 6878 34848 7198 35872
rect 6878 34784 6886 34848
rect 6950 34784 6966 34848
rect 7030 34784 7046 34848
rect 7110 34784 7126 34848
rect 7190 34784 7198 34848
rect 6878 33760 7198 34784
rect 6878 33696 6886 33760
rect 6950 33696 6966 33760
rect 7030 33696 7046 33760
rect 7110 33696 7126 33760
rect 7190 33696 7198 33760
rect 6878 32672 7198 33696
rect 6878 32608 6886 32672
rect 6950 32608 6966 32672
rect 7030 32608 7046 32672
rect 7110 32608 7126 32672
rect 7190 32608 7198 32672
rect 6878 31584 7198 32608
rect 6878 31520 6886 31584
rect 6950 31520 6966 31584
rect 7030 31520 7046 31584
rect 7110 31520 7126 31584
rect 7190 31520 7198 31584
rect 6878 30496 7198 31520
rect 7419 31380 7485 31381
rect 7419 31316 7420 31380
rect 7484 31316 7485 31380
rect 7419 31315 7485 31316
rect 6878 30432 6886 30496
rect 6950 30432 6966 30496
rect 7030 30432 7046 30496
rect 7110 30432 7126 30496
rect 7190 30432 7198 30496
rect 6878 29408 7198 30432
rect 6878 29344 6886 29408
rect 6950 29344 6966 29408
rect 7030 29344 7046 29408
rect 7110 29344 7126 29408
rect 7190 29344 7198 29408
rect 6878 28320 7198 29344
rect 6878 28256 6886 28320
rect 6950 28256 6966 28320
rect 7030 28256 7046 28320
rect 7110 28256 7126 28320
rect 7190 28256 7198 28320
rect 6878 27232 7198 28256
rect 6878 27168 6886 27232
rect 6950 27168 6966 27232
rect 7030 27168 7046 27232
rect 7110 27168 7126 27232
rect 7190 27168 7198 27232
rect 6878 26144 7198 27168
rect 6878 26080 6886 26144
rect 6950 26080 6966 26144
rect 7030 26080 7046 26144
rect 7110 26080 7126 26144
rect 7190 26080 7198 26144
rect 6878 25056 7198 26080
rect 6878 24992 6886 25056
rect 6950 24992 6966 25056
rect 7030 24992 7046 25056
rect 7110 24992 7126 25056
rect 7190 24992 7198 25056
rect 6878 23968 7198 24992
rect 6878 23904 6886 23968
rect 6950 23904 6966 23968
rect 7030 23904 7046 23968
rect 7110 23904 7126 23968
rect 7190 23904 7198 23968
rect 6878 22880 7198 23904
rect 6878 22816 6886 22880
rect 6950 22816 6966 22880
rect 7030 22816 7046 22880
rect 7110 22816 7126 22880
rect 7190 22816 7198 22880
rect 6315 10028 6381 10029
rect 6315 9964 6316 10028
rect 6380 9964 6381 10028
rect 6315 9963 6381 9964
rect 6502 1325 6562 22050
rect 6878 21792 7198 22816
rect 6878 21728 6886 21792
rect 6950 21728 6966 21792
rect 7030 21728 7046 21792
rect 7110 21728 7126 21792
rect 7190 21728 7198 21792
rect 6878 20704 7198 21728
rect 6878 20640 6886 20704
rect 6950 20640 6966 20704
rect 7030 20640 7046 20704
rect 7110 20640 7126 20704
rect 7190 20640 7198 20704
rect 6878 19616 7198 20640
rect 6878 19552 6886 19616
rect 6950 19552 6966 19616
rect 7030 19552 7046 19616
rect 7110 19552 7126 19616
rect 7190 19552 7198 19616
rect 6878 18528 7198 19552
rect 6878 18464 6886 18528
rect 6950 18464 6966 18528
rect 7030 18464 7046 18528
rect 7110 18464 7126 18528
rect 7190 18464 7198 18528
rect 6878 17440 7198 18464
rect 6878 17376 6886 17440
rect 6950 17376 6966 17440
rect 7030 17376 7046 17440
rect 7110 17376 7126 17440
rect 7190 17376 7198 17440
rect 6878 16352 7198 17376
rect 6878 16288 6886 16352
rect 6950 16288 6966 16352
rect 7030 16288 7046 16352
rect 7110 16288 7126 16352
rect 7190 16288 7198 16352
rect 6878 15264 7198 16288
rect 6878 15200 6886 15264
rect 6950 15200 6966 15264
rect 7030 15200 7046 15264
rect 7110 15200 7126 15264
rect 7190 15200 7198 15264
rect 6878 14176 7198 15200
rect 6878 14112 6886 14176
rect 6950 14112 6966 14176
rect 7030 14112 7046 14176
rect 7110 14112 7126 14176
rect 7190 14112 7198 14176
rect 6878 13088 7198 14112
rect 6878 13024 6886 13088
rect 6950 13024 6966 13088
rect 7030 13024 7046 13088
rect 7110 13024 7126 13088
rect 7190 13024 7198 13088
rect 6878 12000 7198 13024
rect 6878 11936 6886 12000
rect 6950 11936 6966 12000
rect 7030 11936 7046 12000
rect 7110 11936 7126 12000
rect 7190 11936 7198 12000
rect 6878 10912 7198 11936
rect 7422 11117 7482 31315
rect 7606 31245 7666 42195
rect 7787 42124 7853 42125
rect 7787 42060 7788 42124
rect 7852 42060 7853 42124
rect 7787 42059 7853 42060
rect 8707 42124 8773 42125
rect 8707 42060 8708 42124
rect 8772 42060 8773 42124
rect 8707 42059 8773 42060
rect 7603 31244 7669 31245
rect 7603 31180 7604 31244
rect 7668 31180 7669 31244
rect 7603 31179 7669 31180
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 6878 10848 6886 10912
rect 6950 10848 6966 10912
rect 7030 10848 7046 10912
rect 7110 10848 7126 10912
rect 7190 10848 7198 10912
rect 6878 9824 7198 10848
rect 6878 9760 6886 9824
rect 6950 9760 6966 9824
rect 7030 9760 7046 9824
rect 7110 9760 7126 9824
rect 7190 9760 7198 9824
rect 6878 8736 7198 9760
rect 6878 8672 6886 8736
rect 6950 8672 6966 8736
rect 7030 8672 7046 8736
rect 7110 8672 7126 8736
rect 7190 8672 7198 8736
rect 6878 7648 7198 8672
rect 6878 7584 6886 7648
rect 6950 7584 6966 7648
rect 7030 7584 7046 7648
rect 7110 7584 7126 7648
rect 7190 7584 7198 7648
rect 6878 6560 7198 7584
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 7790 2277 7850 42059
rect 8155 41852 8221 41853
rect 8155 41788 8156 41852
rect 8220 41788 8221 41852
rect 8155 41787 8221 41788
rect 7971 16556 8037 16557
rect 7971 16492 7972 16556
rect 8036 16492 8037 16556
rect 7971 16491 8037 16492
rect 7787 2276 7853 2277
rect 7787 2212 7788 2276
rect 7852 2212 7853 2276
rect 7787 2211 7853 2212
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 6499 1324 6565 1325
rect 6499 1260 6500 1324
rect 6564 1260 6565 1324
rect 6499 1259 6565 1260
rect 6131 1188 6197 1189
rect 6131 1124 6132 1188
rect 6196 1124 6197 1188
rect 6131 1123 6197 1124
rect 6878 1120 7198 2144
rect 7974 1325 8034 16491
rect 8158 2277 8218 41787
rect 8523 41716 8589 41717
rect 8523 41652 8524 41716
rect 8588 41652 8589 41716
rect 8523 41651 8589 41652
rect 8526 2277 8586 41651
rect 8155 2276 8221 2277
rect 8155 2212 8156 2276
rect 8220 2212 8221 2276
rect 8155 2211 8221 2212
rect 8523 2276 8589 2277
rect 8523 2212 8524 2276
rect 8588 2212 8589 2276
rect 8523 2211 8589 2212
rect 8710 1325 8770 42059
rect 9845 41920 10165 42944
rect 12812 43552 13132 43568
rect 12812 43488 12820 43552
rect 12884 43488 12900 43552
rect 12964 43488 12980 43552
rect 13044 43488 13060 43552
rect 13124 43488 13132 43552
rect 11835 42940 11901 42941
rect 11835 42876 11836 42940
rect 11900 42876 11901 42940
rect 11835 42875 11901 42876
rect 12203 42940 12269 42941
rect 12203 42876 12204 42940
rect 12268 42876 12269 42940
rect 12203 42875 12269 42876
rect 12571 42940 12637 42941
rect 12571 42876 12572 42940
rect 12636 42876 12637 42940
rect 12571 42875 12637 42876
rect 9845 41856 9853 41920
rect 9917 41856 9933 41920
rect 9997 41856 10013 41920
rect 10077 41856 10093 41920
rect 10157 41856 10165 41920
rect 9443 41852 9509 41853
rect 9443 41788 9444 41852
rect 9508 41788 9509 41852
rect 9443 41787 9509 41788
rect 8891 37364 8957 37365
rect 8891 37300 8892 37364
rect 8956 37300 8957 37364
rect 8891 37299 8957 37300
rect 8894 2277 8954 37299
rect 9259 26484 9325 26485
rect 9259 26420 9260 26484
rect 9324 26420 9325 26484
rect 9259 26419 9325 26420
rect 9262 21861 9322 26419
rect 9259 21860 9325 21861
rect 9259 21796 9260 21860
rect 9324 21796 9325 21860
rect 9259 21795 9325 21796
rect 9262 20365 9322 21795
rect 9259 20364 9325 20365
rect 9259 20300 9260 20364
rect 9324 20300 9325 20364
rect 9259 20299 9325 20300
rect 9446 2685 9506 41787
rect 9845 40832 10165 41856
rect 9845 40768 9853 40832
rect 9917 40768 9933 40832
rect 9997 40768 10013 40832
rect 10077 40768 10093 40832
rect 10157 40768 10165 40832
rect 9845 39744 10165 40768
rect 9845 39680 9853 39744
rect 9917 39680 9933 39744
rect 9997 39680 10013 39744
rect 10077 39680 10093 39744
rect 10157 39680 10165 39744
rect 9627 38724 9693 38725
rect 9627 38660 9628 38724
rect 9692 38660 9693 38724
rect 9627 38659 9693 38660
rect 9630 33013 9690 38659
rect 9845 38656 10165 39680
rect 9845 38592 9853 38656
rect 9917 38592 9933 38656
rect 9997 38592 10013 38656
rect 10077 38592 10093 38656
rect 10157 38592 10165 38656
rect 9845 37568 10165 38592
rect 11099 37772 11165 37773
rect 11099 37708 11100 37772
rect 11164 37708 11165 37772
rect 11099 37707 11165 37708
rect 9845 37504 9853 37568
rect 9917 37504 9933 37568
rect 9997 37504 10013 37568
rect 10077 37504 10093 37568
rect 10157 37504 10165 37568
rect 9845 36480 10165 37504
rect 9845 36416 9853 36480
rect 9917 36416 9933 36480
rect 9997 36416 10013 36480
rect 10077 36416 10093 36480
rect 10157 36416 10165 36480
rect 9845 35392 10165 36416
rect 10547 35868 10613 35869
rect 10547 35804 10548 35868
rect 10612 35804 10613 35868
rect 10547 35803 10613 35804
rect 9845 35328 9853 35392
rect 9917 35328 9933 35392
rect 9997 35328 10013 35392
rect 10077 35328 10093 35392
rect 10157 35328 10165 35392
rect 9845 34304 10165 35328
rect 9845 34240 9853 34304
rect 9917 34240 9933 34304
rect 9997 34240 10013 34304
rect 10077 34240 10093 34304
rect 10157 34240 10165 34304
rect 9845 33216 10165 34240
rect 9845 33152 9853 33216
rect 9917 33152 9933 33216
rect 9997 33152 10013 33216
rect 10077 33152 10093 33216
rect 10157 33152 10165 33216
rect 9627 33012 9693 33013
rect 9627 32948 9628 33012
rect 9692 32948 9693 33012
rect 9627 32947 9693 32948
rect 9845 32128 10165 33152
rect 10363 32876 10429 32877
rect 10363 32812 10364 32876
rect 10428 32812 10429 32876
rect 10363 32811 10429 32812
rect 9845 32064 9853 32128
rect 9917 32064 9933 32128
rect 9997 32064 10013 32128
rect 10077 32064 10093 32128
rect 10157 32064 10165 32128
rect 9845 31040 10165 32064
rect 9845 30976 9853 31040
rect 9917 30976 9933 31040
rect 9997 30976 10013 31040
rect 10077 30976 10093 31040
rect 10157 30976 10165 31040
rect 9845 29952 10165 30976
rect 9845 29888 9853 29952
rect 9917 29888 9933 29952
rect 9997 29888 10013 29952
rect 10077 29888 10093 29952
rect 10157 29888 10165 29952
rect 9845 28864 10165 29888
rect 9845 28800 9853 28864
rect 9917 28800 9933 28864
rect 9997 28800 10013 28864
rect 10077 28800 10093 28864
rect 10157 28800 10165 28864
rect 9845 27776 10165 28800
rect 10366 28797 10426 32811
rect 10550 29341 10610 35803
rect 10915 33556 10981 33557
rect 10915 33492 10916 33556
rect 10980 33492 10981 33556
rect 10915 33491 10981 33492
rect 10547 29340 10613 29341
rect 10547 29276 10548 29340
rect 10612 29276 10613 29340
rect 10547 29275 10613 29276
rect 10363 28796 10429 28797
rect 10363 28732 10364 28796
rect 10428 28732 10429 28796
rect 10363 28731 10429 28732
rect 9845 27712 9853 27776
rect 9917 27712 9933 27776
rect 9997 27712 10013 27776
rect 10077 27712 10093 27776
rect 10157 27712 10165 27776
rect 9845 26688 10165 27712
rect 9845 26624 9853 26688
rect 9917 26624 9933 26688
rect 9997 26624 10013 26688
rect 10077 26624 10093 26688
rect 10157 26624 10165 26688
rect 9845 25600 10165 26624
rect 9845 25536 9853 25600
rect 9917 25536 9933 25600
rect 9997 25536 10013 25600
rect 10077 25536 10093 25600
rect 10157 25536 10165 25600
rect 9845 24512 10165 25536
rect 10366 25397 10426 28731
rect 10731 25804 10797 25805
rect 10731 25740 10732 25804
rect 10796 25740 10797 25804
rect 10731 25739 10797 25740
rect 10363 25396 10429 25397
rect 10363 25332 10364 25396
rect 10428 25332 10429 25396
rect 10363 25331 10429 25332
rect 9845 24448 9853 24512
rect 9917 24448 9933 24512
rect 9997 24448 10013 24512
rect 10077 24448 10093 24512
rect 10157 24448 10165 24512
rect 9845 23424 10165 24448
rect 9845 23360 9853 23424
rect 9917 23360 9933 23424
rect 9997 23360 10013 23424
rect 10077 23360 10093 23424
rect 10157 23360 10165 23424
rect 9845 22336 10165 23360
rect 9845 22272 9853 22336
rect 9917 22272 9933 22336
rect 9997 22272 10013 22336
rect 10077 22272 10093 22336
rect 10157 22272 10165 22336
rect 9845 21248 10165 22272
rect 9845 21184 9853 21248
rect 9917 21184 9933 21248
rect 9997 21184 10013 21248
rect 10077 21184 10093 21248
rect 10157 21184 10165 21248
rect 9845 20160 10165 21184
rect 9845 20096 9853 20160
rect 9917 20096 9933 20160
rect 9997 20096 10013 20160
rect 10077 20096 10093 20160
rect 10157 20096 10165 20160
rect 9845 19072 10165 20096
rect 10366 19685 10426 25331
rect 10363 19684 10429 19685
rect 10363 19620 10364 19684
rect 10428 19620 10429 19684
rect 10363 19619 10429 19620
rect 9845 19008 9853 19072
rect 9917 19008 9933 19072
rect 9997 19008 10013 19072
rect 10077 19008 10093 19072
rect 10157 19008 10165 19072
rect 9845 17984 10165 19008
rect 9845 17920 9853 17984
rect 9917 17920 9933 17984
rect 9997 17920 10013 17984
rect 10077 17920 10093 17984
rect 10157 17920 10165 17984
rect 9845 16896 10165 17920
rect 10734 17917 10794 25739
rect 10918 24309 10978 33491
rect 10915 24308 10981 24309
rect 10915 24244 10916 24308
rect 10980 24244 10981 24308
rect 10915 24243 10981 24244
rect 11102 22541 11162 37707
rect 11467 35324 11533 35325
rect 11467 35260 11468 35324
rect 11532 35260 11533 35324
rect 11467 35259 11533 35260
rect 11470 30701 11530 35259
rect 11467 30700 11533 30701
rect 11467 30636 11468 30700
rect 11532 30636 11533 30700
rect 11467 30635 11533 30636
rect 11283 26756 11349 26757
rect 11283 26692 11284 26756
rect 11348 26692 11349 26756
rect 11283 26691 11349 26692
rect 11099 22540 11165 22541
rect 11099 22476 11100 22540
rect 11164 22476 11165 22540
rect 11099 22475 11165 22476
rect 11286 19350 11346 26691
rect 11651 23220 11717 23221
rect 11651 23156 11652 23220
rect 11716 23156 11717 23220
rect 11651 23155 11717 23156
rect 11467 22540 11533 22541
rect 11467 22476 11468 22540
rect 11532 22476 11533 22540
rect 11467 22475 11533 22476
rect 10918 19290 11346 19350
rect 10731 17916 10797 17917
rect 10731 17852 10732 17916
rect 10796 17852 10797 17916
rect 10731 17851 10797 17852
rect 9845 16832 9853 16896
rect 9917 16832 9933 16896
rect 9997 16832 10013 16896
rect 10077 16832 10093 16896
rect 10157 16832 10165 16896
rect 9845 15808 10165 16832
rect 9845 15744 9853 15808
rect 9917 15744 9933 15808
rect 9997 15744 10013 15808
rect 10077 15744 10093 15808
rect 10157 15744 10165 15808
rect 9845 14720 10165 15744
rect 9845 14656 9853 14720
rect 9917 14656 9933 14720
rect 9997 14656 10013 14720
rect 10077 14656 10093 14720
rect 10157 14656 10165 14720
rect 9845 13632 10165 14656
rect 10918 13701 10978 19290
rect 10915 13700 10981 13701
rect 10915 13636 10916 13700
rect 10980 13636 10981 13700
rect 10915 13635 10981 13636
rect 9845 13568 9853 13632
rect 9917 13568 9933 13632
rect 9997 13568 10013 13632
rect 10077 13568 10093 13632
rect 10157 13568 10165 13632
rect 9845 12544 10165 13568
rect 10547 12748 10613 12749
rect 10547 12684 10548 12748
rect 10612 12684 10613 12748
rect 10547 12683 10613 12684
rect 9845 12480 9853 12544
rect 9917 12480 9933 12544
rect 9997 12480 10013 12544
rect 10077 12480 10093 12544
rect 10157 12480 10165 12544
rect 9845 11456 10165 12480
rect 9845 11392 9853 11456
rect 9917 11392 9933 11456
rect 9997 11392 10013 11456
rect 10077 11392 10093 11456
rect 10157 11392 10165 11456
rect 9845 10368 10165 11392
rect 9845 10304 9853 10368
rect 9917 10304 9933 10368
rect 9997 10304 10013 10368
rect 10077 10304 10093 10368
rect 10157 10304 10165 10368
rect 9845 9280 10165 10304
rect 9845 9216 9853 9280
rect 9917 9216 9933 9280
rect 9997 9216 10013 9280
rect 10077 9216 10093 9280
rect 10157 9216 10165 9280
rect 9845 8192 10165 9216
rect 9845 8128 9853 8192
rect 9917 8128 9933 8192
rect 9997 8128 10013 8192
rect 10077 8128 10093 8192
rect 10157 8128 10165 8192
rect 9845 7104 10165 8128
rect 9845 7040 9853 7104
rect 9917 7040 9933 7104
rect 9997 7040 10013 7104
rect 10077 7040 10093 7104
rect 10157 7040 10165 7104
rect 9845 6016 10165 7040
rect 10550 6085 10610 12683
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 10547 6084 10613 6085
rect 10547 6020 10548 6084
rect 10612 6020 10613 6084
rect 10547 6019 10613 6020
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 8891 2276 8957 2277
rect 8891 2212 8892 2276
rect 8956 2212 8957 2276
rect 8891 2211 8957 2212
rect 9845 1664 10165 2688
rect 10550 2413 10610 6019
rect 10918 3365 10978 11051
rect 11470 10709 11530 22475
rect 11654 19005 11714 23155
rect 11651 19004 11717 19005
rect 11651 18940 11652 19004
rect 11716 18940 11717 19004
rect 11651 18939 11717 18940
rect 11654 15197 11714 18939
rect 11651 15196 11717 15197
rect 11651 15132 11652 15196
rect 11716 15132 11717 15196
rect 11651 15131 11717 15132
rect 11651 12748 11717 12749
rect 11651 12684 11652 12748
rect 11716 12684 11717 12748
rect 11651 12683 11717 12684
rect 11467 10708 11533 10709
rect 11467 10644 11468 10708
rect 11532 10644 11533 10708
rect 11467 10643 11533 10644
rect 11654 5949 11714 12683
rect 11838 11117 11898 42875
rect 12019 31788 12085 31789
rect 12019 31724 12020 31788
rect 12084 31724 12085 31788
rect 12019 31723 12085 31724
rect 12022 22949 12082 31723
rect 12206 24717 12266 42875
rect 12203 24716 12269 24717
rect 12203 24652 12204 24716
rect 12268 24652 12269 24716
rect 12203 24651 12269 24652
rect 12019 22948 12085 22949
rect 12019 22884 12020 22948
rect 12084 22884 12085 22948
rect 12019 22883 12085 22884
rect 12019 17916 12085 17917
rect 12019 17852 12020 17916
rect 12084 17852 12085 17916
rect 12019 17851 12085 17852
rect 11835 11116 11901 11117
rect 11835 11052 11836 11116
rect 11900 11052 11901 11116
rect 11835 11051 11901 11052
rect 11651 5948 11717 5949
rect 11651 5884 11652 5948
rect 11716 5884 11717 5948
rect 11651 5883 11717 5884
rect 10915 3364 10981 3365
rect 10915 3300 10916 3364
rect 10980 3300 10981 3364
rect 10915 3299 10981 3300
rect 12022 2413 12082 17851
rect 12387 13292 12453 13293
rect 12387 13228 12388 13292
rect 12452 13228 12453 13292
rect 12387 13227 12453 13228
rect 12390 12450 12450 13227
rect 12206 12390 12450 12450
rect 12206 9890 12266 12390
rect 12574 10573 12634 42875
rect 12812 42464 13132 43488
rect 15779 43008 16099 43568
rect 15779 42944 15787 43008
rect 15851 42944 15867 43008
rect 15931 42944 15947 43008
rect 16011 42944 16027 43008
rect 16091 42944 16099 43008
rect 13859 42940 13925 42941
rect 13859 42876 13860 42940
rect 13924 42876 13925 42940
rect 13859 42875 13925 42876
rect 14411 42940 14477 42941
rect 14411 42876 14412 42940
rect 14476 42876 14477 42940
rect 14411 42875 14477 42876
rect 14963 42940 15029 42941
rect 14963 42876 14964 42940
rect 15028 42876 15029 42940
rect 14963 42875 15029 42876
rect 15515 42940 15581 42941
rect 15515 42876 15516 42940
rect 15580 42876 15581 42940
rect 15515 42875 15581 42876
rect 12812 42400 12820 42464
rect 12884 42400 12900 42464
rect 12964 42400 12980 42464
rect 13044 42400 13060 42464
rect 13124 42400 13132 42464
rect 12812 41376 13132 42400
rect 12812 41312 12820 41376
rect 12884 41312 12900 41376
rect 12964 41312 12980 41376
rect 13044 41312 13060 41376
rect 13124 41312 13132 41376
rect 12812 40288 13132 41312
rect 12812 40224 12820 40288
rect 12884 40224 12900 40288
rect 12964 40224 12980 40288
rect 13044 40224 13060 40288
rect 13124 40224 13132 40288
rect 12812 39200 13132 40224
rect 12812 39136 12820 39200
rect 12884 39136 12900 39200
rect 12964 39136 12980 39200
rect 13044 39136 13060 39200
rect 13124 39136 13132 39200
rect 12812 38112 13132 39136
rect 12812 38048 12820 38112
rect 12884 38048 12900 38112
rect 12964 38048 12980 38112
rect 13044 38048 13060 38112
rect 13124 38048 13132 38112
rect 12812 37024 13132 38048
rect 12812 36960 12820 37024
rect 12884 36960 12900 37024
rect 12964 36960 12980 37024
rect 13044 36960 13060 37024
rect 13124 36960 13132 37024
rect 12812 35936 13132 36960
rect 12812 35872 12820 35936
rect 12884 35872 12900 35936
rect 12964 35872 12980 35936
rect 13044 35872 13060 35936
rect 13124 35872 13132 35936
rect 12812 34848 13132 35872
rect 13307 35052 13373 35053
rect 13307 34988 13308 35052
rect 13372 34988 13373 35052
rect 13307 34987 13373 34988
rect 12812 34784 12820 34848
rect 12884 34784 12900 34848
rect 12964 34784 12980 34848
rect 13044 34784 13060 34848
rect 13124 34784 13132 34848
rect 12812 33760 13132 34784
rect 12812 33696 12820 33760
rect 12884 33696 12900 33760
rect 12964 33696 12980 33760
rect 13044 33696 13060 33760
rect 13124 33696 13132 33760
rect 12812 32672 13132 33696
rect 12812 32608 12820 32672
rect 12884 32608 12900 32672
rect 12964 32608 12980 32672
rect 13044 32608 13060 32672
rect 13124 32608 13132 32672
rect 12812 31584 13132 32608
rect 12812 31520 12820 31584
rect 12884 31520 12900 31584
rect 12964 31520 12980 31584
rect 13044 31520 13060 31584
rect 13124 31520 13132 31584
rect 12812 30496 13132 31520
rect 12812 30432 12820 30496
rect 12884 30432 12900 30496
rect 12964 30432 12980 30496
rect 13044 30432 13060 30496
rect 13124 30432 13132 30496
rect 12812 29408 13132 30432
rect 12812 29344 12820 29408
rect 12884 29344 12900 29408
rect 12964 29344 12980 29408
rect 13044 29344 13060 29408
rect 13124 29344 13132 29408
rect 12812 28320 13132 29344
rect 12812 28256 12820 28320
rect 12884 28256 12900 28320
rect 12964 28256 12980 28320
rect 13044 28256 13060 28320
rect 13124 28256 13132 28320
rect 12812 27232 13132 28256
rect 12812 27168 12820 27232
rect 12884 27168 12900 27232
rect 12964 27168 12980 27232
rect 13044 27168 13060 27232
rect 13124 27168 13132 27232
rect 12812 26144 13132 27168
rect 12812 26080 12820 26144
rect 12884 26080 12900 26144
rect 12964 26080 12980 26144
rect 13044 26080 13060 26144
rect 13124 26080 13132 26144
rect 12812 25056 13132 26080
rect 12812 24992 12820 25056
rect 12884 24992 12900 25056
rect 12964 24992 12980 25056
rect 13044 24992 13060 25056
rect 13124 24992 13132 25056
rect 12812 23968 13132 24992
rect 12812 23904 12820 23968
rect 12884 23904 12900 23968
rect 12964 23904 12980 23968
rect 13044 23904 13060 23968
rect 13124 23904 13132 23968
rect 12812 22880 13132 23904
rect 12812 22816 12820 22880
rect 12884 22816 12900 22880
rect 12964 22816 12980 22880
rect 13044 22816 13060 22880
rect 13124 22816 13132 22880
rect 12812 21792 13132 22816
rect 12812 21728 12820 21792
rect 12884 21728 12900 21792
rect 12964 21728 12980 21792
rect 13044 21728 13060 21792
rect 13124 21728 13132 21792
rect 12812 20704 13132 21728
rect 12812 20640 12820 20704
rect 12884 20640 12900 20704
rect 12964 20640 12980 20704
rect 13044 20640 13060 20704
rect 13124 20640 13132 20704
rect 12812 19616 13132 20640
rect 12812 19552 12820 19616
rect 12884 19552 12900 19616
rect 12964 19552 12980 19616
rect 13044 19552 13060 19616
rect 13124 19552 13132 19616
rect 12812 18528 13132 19552
rect 12812 18464 12820 18528
rect 12884 18464 12900 18528
rect 12964 18464 12980 18528
rect 13044 18464 13060 18528
rect 13124 18464 13132 18528
rect 12812 17440 13132 18464
rect 12812 17376 12820 17440
rect 12884 17376 12900 17440
rect 12964 17376 12980 17440
rect 13044 17376 13060 17440
rect 13124 17376 13132 17440
rect 12812 16352 13132 17376
rect 12812 16288 12820 16352
rect 12884 16288 12900 16352
rect 12964 16288 12980 16352
rect 13044 16288 13060 16352
rect 13124 16288 13132 16352
rect 12812 15264 13132 16288
rect 12812 15200 12820 15264
rect 12884 15200 12900 15264
rect 12964 15200 12980 15264
rect 13044 15200 13060 15264
rect 13124 15200 13132 15264
rect 12812 14176 13132 15200
rect 12812 14112 12820 14176
rect 12884 14112 12900 14176
rect 12964 14112 12980 14176
rect 13044 14112 13060 14176
rect 13124 14112 13132 14176
rect 12812 13088 13132 14112
rect 12812 13024 12820 13088
rect 12884 13024 12900 13088
rect 12964 13024 12980 13088
rect 13044 13024 13060 13088
rect 13124 13024 13132 13088
rect 12812 12000 13132 13024
rect 12812 11936 12820 12000
rect 12884 11936 12900 12000
rect 12964 11936 12980 12000
rect 13044 11936 13060 12000
rect 13124 11936 13132 12000
rect 12812 10912 13132 11936
rect 12812 10848 12820 10912
rect 12884 10848 12900 10912
rect 12964 10848 12980 10912
rect 13044 10848 13060 10912
rect 13124 10848 13132 10912
rect 12571 10572 12637 10573
rect 12571 10508 12572 10572
rect 12636 10508 12637 10572
rect 12571 10507 12637 10508
rect 12206 9830 12634 9890
rect 12203 9756 12269 9757
rect 12203 9692 12204 9756
rect 12268 9692 12269 9756
rect 12203 9691 12269 9692
rect 12206 4045 12266 9691
rect 12203 4044 12269 4045
rect 12203 3980 12204 4044
rect 12268 3980 12269 4044
rect 12203 3979 12269 3980
rect 12574 3365 12634 9830
rect 12812 9824 13132 10848
rect 12812 9760 12820 9824
rect 12884 9760 12900 9824
rect 12964 9760 12980 9824
rect 13044 9760 13060 9824
rect 13124 9760 13132 9824
rect 12812 8736 13132 9760
rect 12812 8672 12820 8736
rect 12884 8672 12900 8736
rect 12964 8672 12980 8736
rect 13044 8672 13060 8736
rect 13124 8672 13132 8736
rect 12812 7648 13132 8672
rect 12812 7584 12820 7648
rect 12884 7584 12900 7648
rect 12964 7584 12980 7648
rect 13044 7584 13060 7648
rect 13124 7584 13132 7648
rect 12812 6560 13132 7584
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12571 3364 12637 3365
rect 12571 3300 12572 3364
rect 12636 3300 12637 3364
rect 12571 3299 12637 3300
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 10547 2412 10613 2413
rect 10547 2348 10548 2412
rect 10612 2348 10613 2412
rect 10547 2347 10613 2348
rect 12019 2412 12085 2413
rect 12019 2348 12020 2412
rect 12084 2348 12085 2412
rect 12019 2347 12085 2348
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 7971 1324 8037 1325
rect 7971 1260 7972 1324
rect 8036 1260 8037 1324
rect 7971 1259 8037 1260
rect 8707 1324 8773 1325
rect 8707 1260 8708 1324
rect 8772 1260 8773 1324
rect 8707 1259 8773 1260
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 1040 10165 1600
rect 12812 2208 13132 3232
rect 13310 2685 13370 34987
rect 13491 29612 13557 29613
rect 13491 29548 13492 29612
rect 13556 29548 13557 29612
rect 13491 29547 13557 29548
rect 13494 23493 13554 29547
rect 13675 28524 13741 28525
rect 13675 28460 13676 28524
rect 13740 28460 13741 28524
rect 13675 28459 13741 28460
rect 13491 23492 13557 23493
rect 13491 23428 13492 23492
rect 13556 23428 13557 23492
rect 13491 23427 13557 23428
rect 13678 23357 13738 28459
rect 13675 23356 13741 23357
rect 13675 23292 13676 23356
rect 13740 23292 13741 23356
rect 13675 23291 13741 23292
rect 13675 22948 13741 22949
rect 13675 22884 13676 22948
rect 13740 22884 13741 22948
rect 13675 22883 13741 22884
rect 13678 18733 13738 22883
rect 13675 18732 13741 18733
rect 13675 18668 13676 18732
rect 13740 18668 13741 18732
rect 13675 18667 13741 18668
rect 13862 8261 13922 42875
rect 14414 15469 14474 42875
rect 14595 18052 14661 18053
rect 14595 17988 14596 18052
rect 14660 17988 14661 18052
rect 14595 17987 14661 17988
rect 14411 15468 14477 15469
rect 14411 15404 14412 15468
rect 14476 15404 14477 15468
rect 14411 15403 14477 15404
rect 13859 8260 13925 8261
rect 13859 8196 13860 8260
rect 13924 8196 13925 8260
rect 13859 8195 13925 8196
rect 14598 4045 14658 17987
rect 14966 7309 15026 42875
rect 15518 18053 15578 42875
rect 15779 41920 16099 42944
rect 15779 41856 15787 41920
rect 15851 41856 15867 41920
rect 15931 41856 15947 41920
rect 16011 41856 16027 41920
rect 16091 41856 16099 41920
rect 15779 40832 16099 41856
rect 18746 43552 19066 43568
rect 18746 43488 18754 43552
rect 18818 43488 18834 43552
rect 18898 43488 18914 43552
rect 18978 43488 18994 43552
rect 19058 43488 19066 43552
rect 18746 42464 19066 43488
rect 18746 42400 18754 42464
rect 18818 42400 18834 42464
rect 18898 42400 18914 42464
rect 18978 42400 18994 42464
rect 19058 42400 19066 42464
rect 17539 41852 17605 41853
rect 17539 41788 17540 41852
rect 17604 41788 17605 41852
rect 17539 41787 17605 41788
rect 16435 41716 16501 41717
rect 16435 41652 16436 41716
rect 16500 41652 16501 41716
rect 16435 41651 16501 41652
rect 17355 41716 17421 41717
rect 17355 41652 17356 41716
rect 17420 41652 17421 41716
rect 17355 41651 17421 41652
rect 15779 40768 15787 40832
rect 15851 40768 15867 40832
rect 15931 40768 15947 40832
rect 16011 40768 16027 40832
rect 16091 40768 16099 40832
rect 15779 39744 16099 40768
rect 15779 39680 15787 39744
rect 15851 39680 15867 39744
rect 15931 39680 15947 39744
rect 16011 39680 16027 39744
rect 16091 39680 16099 39744
rect 15779 38656 16099 39680
rect 15779 38592 15787 38656
rect 15851 38592 15867 38656
rect 15931 38592 15947 38656
rect 16011 38592 16027 38656
rect 16091 38592 16099 38656
rect 15779 37568 16099 38592
rect 15779 37504 15787 37568
rect 15851 37504 15867 37568
rect 15931 37504 15947 37568
rect 16011 37504 16027 37568
rect 16091 37504 16099 37568
rect 15779 36480 16099 37504
rect 15779 36416 15787 36480
rect 15851 36416 15867 36480
rect 15931 36416 15947 36480
rect 16011 36416 16027 36480
rect 16091 36416 16099 36480
rect 15779 35392 16099 36416
rect 15779 35328 15787 35392
rect 15851 35328 15867 35392
rect 15931 35328 15947 35392
rect 16011 35328 16027 35392
rect 16091 35328 16099 35392
rect 15779 34304 16099 35328
rect 15779 34240 15787 34304
rect 15851 34240 15867 34304
rect 15931 34240 15947 34304
rect 16011 34240 16027 34304
rect 16091 34240 16099 34304
rect 15779 33216 16099 34240
rect 15779 33152 15787 33216
rect 15851 33152 15867 33216
rect 15931 33152 15947 33216
rect 16011 33152 16027 33216
rect 16091 33152 16099 33216
rect 15779 32128 16099 33152
rect 15779 32064 15787 32128
rect 15851 32064 15867 32128
rect 15931 32064 15947 32128
rect 16011 32064 16027 32128
rect 16091 32064 16099 32128
rect 15779 31040 16099 32064
rect 15779 30976 15787 31040
rect 15851 30976 15867 31040
rect 15931 30976 15947 31040
rect 16011 30976 16027 31040
rect 16091 30976 16099 31040
rect 15779 29952 16099 30976
rect 15779 29888 15787 29952
rect 15851 29888 15867 29952
rect 15931 29888 15947 29952
rect 16011 29888 16027 29952
rect 16091 29888 16099 29952
rect 15779 28864 16099 29888
rect 16251 29068 16317 29069
rect 16251 29004 16252 29068
rect 16316 29004 16317 29068
rect 16251 29003 16317 29004
rect 15779 28800 15787 28864
rect 15851 28800 15867 28864
rect 15931 28800 15947 28864
rect 16011 28800 16027 28864
rect 16091 28800 16099 28864
rect 15779 27776 16099 28800
rect 16254 27845 16314 29003
rect 16251 27844 16317 27845
rect 16251 27780 16252 27844
rect 16316 27780 16317 27844
rect 16251 27779 16317 27780
rect 15779 27712 15787 27776
rect 15851 27712 15867 27776
rect 15931 27712 15947 27776
rect 16011 27712 16027 27776
rect 16091 27712 16099 27776
rect 15779 26688 16099 27712
rect 15779 26624 15787 26688
rect 15851 26624 15867 26688
rect 15931 26624 15947 26688
rect 16011 26624 16027 26688
rect 16091 26624 16099 26688
rect 15779 25600 16099 26624
rect 15779 25536 15787 25600
rect 15851 25536 15867 25600
rect 15931 25536 15947 25600
rect 16011 25536 16027 25600
rect 16091 25536 16099 25600
rect 15779 24512 16099 25536
rect 15779 24448 15787 24512
rect 15851 24448 15867 24512
rect 15931 24448 15947 24512
rect 16011 24448 16027 24512
rect 16091 24448 16099 24512
rect 15779 23424 16099 24448
rect 15779 23360 15787 23424
rect 15851 23360 15867 23424
rect 15931 23360 15947 23424
rect 16011 23360 16027 23424
rect 16091 23360 16099 23424
rect 15779 22336 16099 23360
rect 15779 22272 15787 22336
rect 15851 22272 15867 22336
rect 15931 22272 15947 22336
rect 16011 22272 16027 22336
rect 16091 22272 16099 22336
rect 15779 21248 16099 22272
rect 15779 21184 15787 21248
rect 15851 21184 15867 21248
rect 15931 21184 15947 21248
rect 16011 21184 16027 21248
rect 16091 21184 16099 21248
rect 15779 20160 16099 21184
rect 15779 20096 15787 20160
rect 15851 20096 15867 20160
rect 15931 20096 15947 20160
rect 16011 20096 16027 20160
rect 16091 20096 16099 20160
rect 15779 19072 16099 20096
rect 15779 19008 15787 19072
rect 15851 19008 15867 19072
rect 15931 19008 15947 19072
rect 16011 19008 16027 19072
rect 16091 19008 16099 19072
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 15779 17984 16099 19008
rect 15779 17920 15787 17984
rect 15851 17920 15867 17984
rect 15931 17920 15947 17984
rect 16011 17920 16027 17984
rect 16091 17920 16099 17984
rect 15779 16896 16099 17920
rect 15779 16832 15787 16896
rect 15851 16832 15867 16896
rect 15931 16832 15947 16896
rect 16011 16832 16027 16896
rect 16091 16832 16099 16896
rect 15515 16012 15581 16013
rect 15515 15948 15516 16012
rect 15580 15948 15581 16012
rect 15515 15947 15581 15948
rect 15518 10845 15578 15947
rect 15779 15808 16099 16832
rect 15779 15744 15787 15808
rect 15851 15744 15867 15808
rect 15931 15744 15947 15808
rect 16011 15744 16027 15808
rect 16091 15744 16099 15808
rect 15779 14720 16099 15744
rect 16251 15196 16317 15197
rect 16251 15132 16252 15196
rect 16316 15132 16317 15196
rect 16251 15131 16317 15132
rect 15779 14656 15787 14720
rect 15851 14656 15867 14720
rect 15931 14656 15947 14720
rect 16011 14656 16027 14720
rect 16091 14656 16099 14720
rect 15779 13632 16099 14656
rect 15779 13568 15787 13632
rect 15851 13568 15867 13632
rect 15931 13568 15947 13632
rect 16011 13568 16027 13632
rect 16091 13568 16099 13632
rect 15779 12544 16099 13568
rect 15779 12480 15787 12544
rect 15851 12480 15867 12544
rect 15931 12480 15947 12544
rect 16011 12480 16027 12544
rect 16091 12480 16099 12544
rect 15779 11456 16099 12480
rect 15779 11392 15787 11456
rect 15851 11392 15867 11456
rect 15931 11392 15947 11456
rect 16011 11392 16027 11456
rect 16091 11392 16099 11456
rect 15515 10844 15581 10845
rect 15515 10780 15516 10844
rect 15580 10780 15581 10844
rect 15515 10779 15581 10780
rect 15779 10368 16099 11392
rect 16254 10981 16314 15131
rect 16251 10980 16317 10981
rect 16251 10916 16252 10980
rect 16316 10916 16317 10980
rect 16251 10915 16317 10916
rect 15779 10304 15787 10368
rect 15851 10304 15867 10368
rect 15931 10304 15947 10368
rect 16011 10304 16027 10368
rect 16091 10304 16099 10368
rect 15779 9280 16099 10304
rect 16254 9757 16314 10915
rect 16251 9756 16317 9757
rect 16251 9692 16252 9756
rect 16316 9692 16317 9756
rect 16251 9691 16317 9692
rect 15779 9216 15787 9280
rect 15851 9216 15867 9280
rect 15931 9216 15947 9280
rect 16011 9216 16027 9280
rect 16091 9216 16099 9280
rect 15779 8192 16099 9216
rect 15779 8128 15787 8192
rect 15851 8128 15867 8192
rect 15931 8128 15947 8192
rect 16011 8128 16027 8192
rect 16091 8128 16099 8192
rect 14963 7308 15029 7309
rect 14963 7244 14964 7308
rect 15028 7244 15029 7308
rect 14963 7243 15029 7244
rect 15779 7104 16099 8128
rect 15779 7040 15787 7104
rect 15851 7040 15867 7104
rect 15931 7040 15947 7104
rect 16011 7040 16027 7104
rect 16091 7040 16099 7104
rect 15779 6016 16099 7040
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 14595 4044 14661 4045
rect 14595 3980 14596 4044
rect 14660 3980 14661 4044
rect 14595 3979 14661 3980
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 13307 2684 13373 2685
rect 13307 2620 13308 2684
rect 13372 2620 13373 2684
rect 13307 2619 13373 2620
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 16438 1325 16498 41651
rect 16619 29204 16685 29205
rect 16619 29140 16620 29204
rect 16684 29140 16685 29204
rect 16619 29139 16685 29140
rect 16622 25261 16682 29139
rect 16803 28796 16869 28797
rect 16803 28732 16804 28796
rect 16868 28732 16869 28796
rect 16803 28731 16869 28732
rect 16619 25260 16685 25261
rect 16619 25196 16620 25260
rect 16684 25196 16685 25260
rect 16619 25195 16685 25196
rect 16806 21725 16866 28731
rect 17171 28660 17237 28661
rect 17171 28596 17172 28660
rect 17236 28596 17237 28660
rect 17171 28595 17237 28596
rect 16803 21724 16869 21725
rect 16803 21660 16804 21724
rect 16868 21660 16869 21724
rect 16803 21659 16869 21660
rect 17174 19005 17234 28595
rect 17171 19004 17237 19005
rect 17171 18940 17172 19004
rect 17236 18940 17237 19004
rect 17171 18939 17237 18940
rect 16987 18188 17053 18189
rect 16987 18124 16988 18188
rect 17052 18124 17053 18188
rect 16987 18123 17053 18124
rect 16990 5133 17050 18123
rect 16987 5132 17053 5133
rect 16987 5068 16988 5132
rect 17052 5068 17053 5132
rect 16987 5067 17053 5068
rect 17358 2685 17418 41651
rect 17542 27709 17602 41787
rect 18459 41716 18525 41717
rect 18459 41652 18460 41716
rect 18524 41652 18525 41716
rect 18459 41651 18525 41652
rect 18275 41444 18341 41445
rect 18275 41380 18276 41444
rect 18340 41380 18341 41444
rect 18275 41379 18341 41380
rect 17907 37908 17973 37909
rect 17907 37844 17908 37908
rect 17972 37844 17973 37908
rect 17907 37843 17973 37844
rect 17539 27708 17605 27709
rect 17539 27644 17540 27708
rect 17604 27644 17605 27708
rect 17539 27643 17605 27644
rect 17539 23084 17605 23085
rect 17539 23020 17540 23084
rect 17604 23020 17605 23084
rect 17539 23019 17605 23020
rect 17542 3773 17602 23019
rect 17723 17780 17789 17781
rect 17723 17716 17724 17780
rect 17788 17716 17789 17780
rect 17723 17715 17789 17716
rect 17539 3772 17605 3773
rect 17539 3708 17540 3772
rect 17604 3708 17605 3772
rect 17539 3707 17605 3708
rect 17355 2684 17421 2685
rect 17355 2620 17356 2684
rect 17420 2620 17421 2684
rect 17355 2619 17421 2620
rect 17726 2413 17786 17715
rect 17910 7581 17970 37843
rect 17907 7580 17973 7581
rect 17907 7516 17908 7580
rect 17972 7516 17973 7580
rect 17907 7515 17973 7516
rect 18278 4045 18338 41379
rect 18275 4044 18341 4045
rect 18275 3980 18276 4044
rect 18340 3980 18341 4044
rect 18275 3979 18341 3980
rect 18462 2685 18522 41651
rect 18746 41376 19066 42400
rect 21713 43008 22033 43568
rect 21713 42944 21721 43008
rect 21785 42944 21801 43008
rect 21865 42944 21881 43008
rect 21945 42944 21961 43008
rect 22025 42944 22033 43008
rect 21713 41920 22033 42944
rect 21713 41856 21721 41920
rect 21785 41856 21801 41920
rect 21865 41856 21881 41920
rect 21945 41856 21961 41920
rect 22025 41856 22033 41920
rect 19379 41716 19445 41717
rect 19379 41652 19380 41716
rect 19444 41652 19445 41716
rect 19379 41651 19445 41652
rect 18746 41312 18754 41376
rect 18818 41312 18834 41376
rect 18898 41312 18914 41376
rect 18978 41312 18994 41376
rect 19058 41312 19066 41376
rect 18746 40288 19066 41312
rect 18746 40224 18754 40288
rect 18818 40224 18834 40288
rect 18898 40224 18914 40288
rect 18978 40224 18994 40288
rect 19058 40224 19066 40288
rect 18746 39200 19066 40224
rect 18746 39136 18754 39200
rect 18818 39136 18834 39200
rect 18898 39136 18914 39200
rect 18978 39136 18994 39200
rect 19058 39136 19066 39200
rect 18746 38112 19066 39136
rect 18746 38048 18754 38112
rect 18818 38048 18834 38112
rect 18898 38048 18914 38112
rect 18978 38048 18994 38112
rect 19058 38048 19066 38112
rect 18746 37024 19066 38048
rect 18746 36960 18754 37024
rect 18818 36960 18834 37024
rect 18898 36960 18914 37024
rect 18978 36960 18994 37024
rect 19058 36960 19066 37024
rect 18746 35936 19066 36960
rect 18746 35872 18754 35936
rect 18818 35872 18834 35936
rect 18898 35872 18914 35936
rect 18978 35872 18994 35936
rect 19058 35872 19066 35936
rect 18746 34848 19066 35872
rect 18746 34784 18754 34848
rect 18818 34784 18834 34848
rect 18898 34784 18914 34848
rect 18978 34784 18994 34848
rect 19058 34784 19066 34848
rect 18746 33760 19066 34784
rect 18746 33696 18754 33760
rect 18818 33696 18834 33760
rect 18898 33696 18914 33760
rect 18978 33696 18994 33760
rect 19058 33696 19066 33760
rect 18746 32672 19066 33696
rect 18746 32608 18754 32672
rect 18818 32608 18834 32672
rect 18898 32608 18914 32672
rect 18978 32608 18994 32672
rect 19058 32608 19066 32672
rect 18746 31584 19066 32608
rect 18746 31520 18754 31584
rect 18818 31520 18834 31584
rect 18898 31520 18914 31584
rect 18978 31520 18994 31584
rect 19058 31520 19066 31584
rect 18746 30496 19066 31520
rect 18746 30432 18754 30496
rect 18818 30432 18834 30496
rect 18898 30432 18914 30496
rect 18978 30432 18994 30496
rect 19058 30432 19066 30496
rect 18746 29408 19066 30432
rect 18746 29344 18754 29408
rect 18818 29344 18834 29408
rect 18898 29344 18914 29408
rect 18978 29344 18994 29408
rect 19058 29344 19066 29408
rect 18746 28320 19066 29344
rect 18746 28256 18754 28320
rect 18818 28256 18834 28320
rect 18898 28256 18914 28320
rect 18978 28256 18994 28320
rect 19058 28256 19066 28320
rect 18746 27232 19066 28256
rect 18746 27168 18754 27232
rect 18818 27168 18834 27232
rect 18898 27168 18914 27232
rect 18978 27168 18994 27232
rect 19058 27168 19066 27232
rect 18746 26144 19066 27168
rect 18746 26080 18754 26144
rect 18818 26080 18834 26144
rect 18898 26080 18914 26144
rect 18978 26080 18994 26144
rect 19058 26080 19066 26144
rect 18746 25056 19066 26080
rect 18746 24992 18754 25056
rect 18818 24992 18834 25056
rect 18898 24992 18914 25056
rect 18978 24992 18994 25056
rect 19058 24992 19066 25056
rect 18746 23968 19066 24992
rect 18746 23904 18754 23968
rect 18818 23904 18834 23968
rect 18898 23904 18914 23968
rect 18978 23904 18994 23968
rect 19058 23904 19066 23968
rect 18746 22880 19066 23904
rect 18746 22816 18754 22880
rect 18818 22816 18834 22880
rect 18898 22816 18914 22880
rect 18978 22816 18994 22880
rect 19058 22816 19066 22880
rect 18746 21792 19066 22816
rect 18746 21728 18754 21792
rect 18818 21728 18834 21792
rect 18898 21728 18914 21792
rect 18978 21728 18994 21792
rect 19058 21728 19066 21792
rect 18746 20704 19066 21728
rect 18746 20640 18754 20704
rect 18818 20640 18834 20704
rect 18898 20640 18914 20704
rect 18978 20640 18994 20704
rect 19058 20640 19066 20704
rect 18746 19616 19066 20640
rect 18746 19552 18754 19616
rect 18818 19552 18834 19616
rect 18898 19552 18914 19616
rect 18978 19552 18994 19616
rect 19058 19552 19066 19616
rect 18746 18528 19066 19552
rect 18746 18464 18754 18528
rect 18818 18464 18834 18528
rect 18898 18464 18914 18528
rect 18978 18464 18994 18528
rect 19058 18464 19066 18528
rect 18746 17440 19066 18464
rect 18746 17376 18754 17440
rect 18818 17376 18834 17440
rect 18898 17376 18914 17440
rect 18978 17376 18994 17440
rect 19058 17376 19066 17440
rect 18746 16352 19066 17376
rect 18746 16288 18754 16352
rect 18818 16288 18834 16352
rect 18898 16288 18914 16352
rect 18978 16288 18994 16352
rect 19058 16288 19066 16352
rect 18746 15264 19066 16288
rect 18746 15200 18754 15264
rect 18818 15200 18834 15264
rect 18898 15200 18914 15264
rect 18978 15200 18994 15264
rect 19058 15200 19066 15264
rect 18746 14176 19066 15200
rect 18746 14112 18754 14176
rect 18818 14112 18834 14176
rect 18898 14112 18914 14176
rect 18978 14112 18994 14176
rect 19058 14112 19066 14176
rect 18746 13088 19066 14112
rect 18746 13024 18754 13088
rect 18818 13024 18834 13088
rect 18898 13024 18914 13088
rect 18978 13024 18994 13088
rect 19058 13024 19066 13088
rect 18746 12000 19066 13024
rect 18746 11936 18754 12000
rect 18818 11936 18834 12000
rect 18898 11936 18914 12000
rect 18978 11936 18994 12000
rect 19058 11936 19066 12000
rect 18746 10912 19066 11936
rect 19382 11117 19442 41651
rect 21713 40832 22033 41856
rect 21713 40768 21721 40832
rect 21785 40768 21801 40832
rect 21865 40768 21881 40832
rect 21945 40768 21961 40832
rect 22025 40768 22033 40832
rect 21713 39744 22033 40768
rect 24680 43552 25000 43568
rect 24680 43488 24688 43552
rect 24752 43488 24768 43552
rect 24832 43488 24848 43552
rect 24912 43488 24928 43552
rect 24992 43488 25000 43552
rect 24680 42464 25000 43488
rect 24680 42400 24688 42464
rect 24752 42400 24768 42464
rect 24832 42400 24848 42464
rect 24912 42400 24928 42464
rect 24992 42400 25000 42464
rect 24680 41376 25000 42400
rect 24680 41312 24688 41376
rect 24752 41312 24768 41376
rect 24832 41312 24848 41376
rect 24912 41312 24928 41376
rect 24992 41312 25000 41376
rect 24680 40288 25000 41312
rect 24680 40224 24688 40288
rect 24752 40224 24768 40288
rect 24832 40224 24848 40288
rect 24912 40224 24928 40288
rect 24992 40224 25000 40288
rect 22875 40220 22941 40221
rect 22875 40156 22876 40220
rect 22940 40156 22941 40220
rect 22875 40155 22941 40156
rect 21713 39680 21721 39744
rect 21785 39680 21801 39744
rect 21865 39680 21881 39744
rect 21945 39680 21961 39744
rect 22025 39680 22033 39744
rect 19563 38724 19629 38725
rect 19563 38660 19564 38724
rect 19628 38660 19629 38724
rect 19563 38659 19629 38660
rect 19379 11116 19445 11117
rect 19379 11052 19380 11116
rect 19444 11052 19445 11116
rect 19379 11051 19445 11052
rect 18746 10848 18754 10912
rect 18818 10848 18834 10912
rect 18898 10848 18914 10912
rect 18978 10848 18994 10912
rect 19058 10848 19066 10912
rect 18746 9824 19066 10848
rect 18746 9760 18754 9824
rect 18818 9760 18834 9824
rect 18898 9760 18914 9824
rect 18978 9760 18994 9824
rect 19058 9760 19066 9824
rect 18746 8736 19066 9760
rect 18746 8672 18754 8736
rect 18818 8672 18834 8736
rect 18898 8672 18914 8736
rect 18978 8672 18994 8736
rect 19058 8672 19066 8736
rect 18746 7648 19066 8672
rect 18746 7584 18754 7648
rect 18818 7584 18834 7648
rect 18898 7584 18914 7648
rect 18978 7584 18994 7648
rect 19058 7584 19066 7648
rect 18746 6560 19066 7584
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 19195 3772 19261 3773
rect 19195 3708 19196 3772
rect 19260 3708 19261 3772
rect 19195 3707 19261 3708
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18459 2684 18525 2685
rect 18459 2620 18460 2684
rect 18524 2620 18525 2684
rect 18459 2619 18525 2620
rect 17723 2412 17789 2413
rect 17723 2348 17724 2412
rect 17788 2348 17789 2412
rect 17723 2347 17789 2348
rect 18746 2208 19066 3232
rect 19198 2685 19258 3707
rect 19566 2685 19626 38659
rect 21713 38656 22033 39680
rect 22878 39130 22938 40155
rect 21713 38592 21721 38656
rect 21785 38592 21801 38656
rect 21865 38592 21881 38656
rect 21945 38592 21961 38656
rect 22025 38592 22033 38656
rect 21713 37568 22033 38592
rect 21713 37504 21721 37568
rect 21785 37504 21801 37568
rect 21865 37504 21881 37568
rect 21945 37504 21961 37568
rect 22025 37504 22033 37568
rect 21713 36480 22033 37504
rect 21713 36416 21721 36480
rect 21785 36416 21801 36480
rect 21865 36416 21881 36480
rect 21945 36416 21961 36480
rect 22025 36416 22033 36480
rect 21713 35392 22033 36416
rect 21713 35328 21721 35392
rect 21785 35328 21801 35392
rect 21865 35328 21881 35392
rect 21945 35328 21961 35392
rect 22025 35328 22033 35392
rect 21713 34304 22033 35328
rect 21713 34240 21721 34304
rect 21785 34240 21801 34304
rect 21865 34240 21881 34304
rect 21945 34240 21961 34304
rect 22025 34240 22033 34304
rect 19931 33420 19997 33421
rect 19931 33356 19932 33420
rect 19996 33356 19997 33420
rect 19931 33355 19997 33356
rect 19747 33284 19813 33285
rect 19747 33220 19748 33284
rect 19812 33220 19813 33284
rect 19747 33219 19813 33220
rect 19750 17917 19810 33219
rect 19747 17916 19813 17917
rect 19747 17852 19748 17916
rect 19812 17852 19813 17916
rect 19747 17851 19813 17852
rect 19934 2685 19994 33355
rect 21713 33216 22033 34240
rect 21713 33152 21721 33216
rect 21785 33152 21801 33216
rect 21865 33152 21881 33216
rect 21945 33152 21961 33216
rect 22025 33152 22033 33216
rect 21713 32128 22033 33152
rect 21713 32064 21721 32128
rect 21785 32064 21801 32128
rect 21865 32064 21881 32128
rect 21945 32064 21961 32128
rect 22025 32064 22033 32128
rect 21035 31244 21101 31245
rect 21035 31180 21036 31244
rect 21100 31180 21101 31244
rect 21035 31179 21101 31180
rect 21038 29010 21098 31179
rect 21713 31040 22033 32064
rect 21713 30976 21721 31040
rect 21785 30976 21801 31040
rect 21865 30976 21881 31040
rect 21945 30976 21961 31040
rect 22025 30976 22033 31040
rect 21587 30428 21653 30429
rect 21587 30364 21588 30428
rect 21652 30364 21653 30428
rect 21587 30363 21653 30364
rect 20486 28950 21098 29010
rect 20486 19350 20546 28950
rect 20667 27980 20733 27981
rect 20667 27916 20668 27980
rect 20732 27916 20733 27980
rect 20667 27915 20733 27916
rect 20670 25258 20730 27915
rect 20851 27708 20917 27709
rect 20851 27644 20852 27708
rect 20916 27644 20917 27708
rect 20851 27643 20917 27644
rect 20854 26893 20914 27643
rect 20851 26892 20917 26893
rect 20851 26828 20852 26892
rect 20916 26828 20917 26892
rect 20851 26827 20917 26828
rect 21590 25261 21650 30363
rect 21713 29952 22033 30976
rect 21713 29888 21721 29952
rect 21785 29888 21801 29952
rect 21865 29888 21881 29952
rect 21945 29888 21961 29952
rect 22025 29888 22033 29952
rect 21713 28864 22033 29888
rect 21713 28800 21721 28864
rect 21785 28800 21801 28864
rect 21865 28800 21881 28864
rect 21945 28800 21961 28864
rect 22025 28800 22033 28864
rect 21713 27776 22033 28800
rect 21713 27712 21721 27776
rect 21785 27712 21801 27776
rect 21865 27712 21881 27776
rect 21945 27712 21961 27776
rect 22025 27712 22033 27776
rect 21713 26688 22033 27712
rect 21713 26624 21721 26688
rect 21785 26624 21801 26688
rect 21865 26624 21881 26688
rect 21945 26624 21961 26688
rect 22025 26624 22033 26688
rect 21713 25600 22033 26624
rect 21713 25536 21721 25600
rect 21785 25536 21801 25600
rect 21865 25536 21881 25600
rect 21945 25536 21961 25600
rect 22025 25536 22033 25600
rect 21587 25260 21653 25261
rect 20670 25198 20914 25258
rect 20486 19290 20730 19350
rect 20299 16420 20365 16421
rect 20299 16356 20300 16420
rect 20364 16356 20365 16420
rect 20299 16355 20365 16356
rect 20302 9893 20362 16355
rect 20299 9892 20365 9893
rect 20299 9828 20300 9892
rect 20364 9828 20365 9892
rect 20299 9827 20365 9828
rect 19195 2684 19261 2685
rect 19195 2620 19196 2684
rect 19260 2620 19261 2684
rect 19195 2619 19261 2620
rect 19563 2684 19629 2685
rect 19563 2620 19564 2684
rect 19628 2620 19629 2684
rect 19563 2619 19629 2620
rect 19931 2684 19997 2685
rect 19931 2620 19932 2684
rect 19996 2620 19997 2684
rect 19931 2619 19997 2620
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 16435 1324 16501 1325
rect 16435 1260 16436 1324
rect 16500 1260 16501 1324
rect 16435 1259 16501 1260
rect 18746 1120 19066 2144
rect 20670 2005 20730 19290
rect 20854 18189 20914 25198
rect 21587 25196 21588 25260
rect 21652 25196 21653 25260
rect 21587 25195 21653 25196
rect 21713 24512 22033 25536
rect 21713 24448 21721 24512
rect 21785 24448 21801 24512
rect 21865 24448 21881 24512
rect 21945 24448 21961 24512
rect 22025 24448 22033 24512
rect 21403 23628 21469 23629
rect 21403 23564 21404 23628
rect 21468 23564 21469 23628
rect 21403 23563 21469 23564
rect 20851 18188 20917 18189
rect 20851 18124 20852 18188
rect 20916 18124 20917 18188
rect 20851 18123 20917 18124
rect 20851 18052 20917 18053
rect 20851 17988 20852 18052
rect 20916 17988 20917 18052
rect 20851 17987 20917 17988
rect 20854 11389 20914 17987
rect 21219 17508 21285 17509
rect 21219 17444 21220 17508
rect 21284 17444 21285 17508
rect 21219 17443 21285 17444
rect 21222 12341 21282 17443
rect 21219 12340 21285 12341
rect 21219 12276 21220 12340
rect 21284 12276 21285 12340
rect 21219 12275 21285 12276
rect 20851 11388 20917 11389
rect 20851 11324 20852 11388
rect 20916 11324 20917 11388
rect 20851 11323 20917 11324
rect 21406 6221 21466 23563
rect 21713 23424 22033 24448
rect 21713 23360 21721 23424
rect 21785 23360 21801 23424
rect 21865 23360 21881 23424
rect 21945 23360 21961 23424
rect 22025 23360 22033 23424
rect 21713 22336 22033 23360
rect 21713 22272 21721 22336
rect 21785 22272 21801 22336
rect 21865 22272 21881 22336
rect 21945 22272 21961 22336
rect 22025 22272 22033 22336
rect 21713 21248 22033 22272
rect 21713 21184 21721 21248
rect 21785 21184 21801 21248
rect 21865 21184 21881 21248
rect 21945 21184 21961 21248
rect 22025 21184 22033 21248
rect 21713 20160 22033 21184
rect 21713 20096 21721 20160
rect 21785 20096 21801 20160
rect 21865 20096 21881 20160
rect 21945 20096 21961 20160
rect 22025 20096 22033 20160
rect 21713 19072 22033 20096
rect 21713 19008 21721 19072
rect 21785 19008 21801 19072
rect 21865 19008 21881 19072
rect 21945 19008 21961 19072
rect 22025 19008 22033 19072
rect 21713 17984 22033 19008
rect 21713 17920 21721 17984
rect 21785 17920 21801 17984
rect 21865 17920 21881 17984
rect 21945 17920 21961 17984
rect 22025 17920 22033 17984
rect 21713 16896 22033 17920
rect 21713 16832 21721 16896
rect 21785 16832 21801 16896
rect 21865 16832 21881 16896
rect 21945 16832 21961 16896
rect 22025 16832 22033 16896
rect 21713 15808 22033 16832
rect 21713 15744 21721 15808
rect 21785 15744 21801 15808
rect 21865 15744 21881 15808
rect 21945 15744 21961 15808
rect 22025 15744 22033 15808
rect 21713 14720 22033 15744
rect 21713 14656 21721 14720
rect 21785 14656 21801 14720
rect 21865 14656 21881 14720
rect 21945 14656 21961 14720
rect 22025 14656 22033 14720
rect 21713 13632 22033 14656
rect 22326 39070 22938 39130
rect 24680 39200 25000 40224
rect 24680 39136 24688 39200
rect 24752 39136 24768 39200
rect 24832 39136 24848 39200
rect 24912 39136 24928 39200
rect 24992 39136 25000 39200
rect 22326 13701 22386 39070
rect 22507 38996 22573 38997
rect 22507 38932 22508 38996
rect 22572 38932 22573 38996
rect 22507 38931 22573 38932
rect 22510 19957 22570 38931
rect 24680 38112 25000 39136
rect 24680 38048 24688 38112
rect 24752 38048 24768 38112
rect 24832 38048 24848 38112
rect 24912 38048 24928 38112
rect 24992 38048 25000 38112
rect 24680 37024 25000 38048
rect 24680 36960 24688 37024
rect 24752 36960 24768 37024
rect 24832 36960 24848 37024
rect 24912 36960 24928 37024
rect 24992 36960 25000 37024
rect 22875 36004 22941 36005
rect 22875 35940 22876 36004
rect 22940 35940 22941 36004
rect 22875 35939 22941 35940
rect 22507 19956 22573 19957
rect 22507 19892 22508 19956
rect 22572 19892 22573 19956
rect 22507 19891 22573 19892
rect 22691 19820 22757 19821
rect 22691 19756 22692 19820
rect 22756 19756 22757 19820
rect 22691 19755 22757 19756
rect 22323 13700 22389 13701
rect 22323 13636 22324 13700
rect 22388 13636 22389 13700
rect 22323 13635 22389 13636
rect 21713 13568 21721 13632
rect 21785 13568 21801 13632
rect 21865 13568 21881 13632
rect 21945 13568 21961 13632
rect 22025 13568 22033 13632
rect 21713 12544 22033 13568
rect 21713 12480 21721 12544
rect 21785 12480 21801 12544
rect 21865 12480 21881 12544
rect 21945 12480 21961 12544
rect 22025 12480 22033 12544
rect 21713 11456 22033 12480
rect 21713 11392 21721 11456
rect 21785 11392 21801 11456
rect 21865 11392 21881 11456
rect 21945 11392 21961 11456
rect 22025 11392 22033 11456
rect 21713 10368 22033 11392
rect 21713 10304 21721 10368
rect 21785 10304 21801 10368
rect 21865 10304 21881 10368
rect 21945 10304 21961 10368
rect 22025 10304 22033 10368
rect 21713 9280 22033 10304
rect 21713 9216 21721 9280
rect 21785 9216 21801 9280
rect 21865 9216 21881 9280
rect 21945 9216 21961 9280
rect 22025 9216 22033 9280
rect 21713 8192 22033 9216
rect 21713 8128 21721 8192
rect 21785 8128 21801 8192
rect 21865 8128 21881 8192
rect 21945 8128 21961 8192
rect 22025 8128 22033 8192
rect 21713 7104 22033 8128
rect 21713 7040 21721 7104
rect 21785 7040 21801 7104
rect 21865 7040 21881 7104
rect 21945 7040 21961 7104
rect 22025 7040 22033 7104
rect 21403 6220 21469 6221
rect 21403 6156 21404 6220
rect 21468 6156 21469 6220
rect 21403 6155 21469 6156
rect 21713 6016 22033 7040
rect 22139 6764 22205 6765
rect 22139 6700 22140 6764
rect 22204 6700 22205 6764
rect 22139 6699 22205 6700
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 22142 3229 22202 6699
rect 22694 5541 22754 19755
rect 22878 5541 22938 35939
rect 24680 35936 25000 36960
rect 24680 35872 24688 35936
rect 24752 35872 24768 35936
rect 24832 35872 24848 35936
rect 24912 35872 24928 35936
rect 24992 35872 25000 35936
rect 24680 34848 25000 35872
rect 24680 34784 24688 34848
rect 24752 34784 24768 34848
rect 24832 34784 24848 34848
rect 24912 34784 24928 34848
rect 24992 34784 25000 34848
rect 24680 33760 25000 34784
rect 24680 33696 24688 33760
rect 24752 33696 24768 33760
rect 24832 33696 24848 33760
rect 24912 33696 24928 33760
rect 24992 33696 25000 33760
rect 24680 32672 25000 33696
rect 24680 32608 24688 32672
rect 24752 32608 24768 32672
rect 24832 32608 24848 32672
rect 24912 32608 24928 32672
rect 24992 32608 25000 32672
rect 24680 31584 25000 32608
rect 24680 31520 24688 31584
rect 24752 31520 24768 31584
rect 24832 31520 24848 31584
rect 24912 31520 24928 31584
rect 24992 31520 25000 31584
rect 24680 30496 25000 31520
rect 24680 30432 24688 30496
rect 24752 30432 24768 30496
rect 24832 30432 24848 30496
rect 24912 30432 24928 30496
rect 24992 30432 25000 30496
rect 24680 29408 25000 30432
rect 24680 29344 24688 29408
rect 24752 29344 24768 29408
rect 24832 29344 24848 29408
rect 24912 29344 24928 29408
rect 24992 29344 25000 29408
rect 24680 28320 25000 29344
rect 24680 28256 24688 28320
rect 24752 28256 24768 28320
rect 24832 28256 24848 28320
rect 24912 28256 24928 28320
rect 24992 28256 25000 28320
rect 24680 27232 25000 28256
rect 24680 27168 24688 27232
rect 24752 27168 24768 27232
rect 24832 27168 24848 27232
rect 24912 27168 24928 27232
rect 24992 27168 25000 27232
rect 24680 26144 25000 27168
rect 24680 26080 24688 26144
rect 24752 26080 24768 26144
rect 24832 26080 24848 26144
rect 24912 26080 24928 26144
rect 24992 26080 25000 26144
rect 24680 25056 25000 26080
rect 24680 24992 24688 25056
rect 24752 24992 24768 25056
rect 24832 24992 24848 25056
rect 24912 24992 24928 25056
rect 24992 24992 25000 25056
rect 24680 23968 25000 24992
rect 24680 23904 24688 23968
rect 24752 23904 24768 23968
rect 24832 23904 24848 23968
rect 24912 23904 24928 23968
rect 24992 23904 25000 23968
rect 24680 22880 25000 23904
rect 24680 22816 24688 22880
rect 24752 22816 24768 22880
rect 24832 22816 24848 22880
rect 24912 22816 24928 22880
rect 24992 22816 25000 22880
rect 24680 21792 25000 22816
rect 24680 21728 24688 21792
rect 24752 21728 24768 21792
rect 24832 21728 24848 21792
rect 24912 21728 24928 21792
rect 24992 21728 25000 21792
rect 24680 20704 25000 21728
rect 24680 20640 24688 20704
rect 24752 20640 24768 20704
rect 24832 20640 24848 20704
rect 24912 20640 24928 20704
rect 24992 20640 25000 20704
rect 24680 19616 25000 20640
rect 24680 19552 24688 19616
rect 24752 19552 24768 19616
rect 24832 19552 24848 19616
rect 24912 19552 24928 19616
rect 24992 19552 25000 19616
rect 24680 18528 25000 19552
rect 24680 18464 24688 18528
rect 24752 18464 24768 18528
rect 24832 18464 24848 18528
rect 24912 18464 24928 18528
rect 24992 18464 25000 18528
rect 24680 17440 25000 18464
rect 24680 17376 24688 17440
rect 24752 17376 24768 17440
rect 24832 17376 24848 17440
rect 24912 17376 24928 17440
rect 24992 17376 25000 17440
rect 24680 16352 25000 17376
rect 24680 16288 24688 16352
rect 24752 16288 24768 16352
rect 24832 16288 24848 16352
rect 24912 16288 24928 16352
rect 24992 16288 25000 16352
rect 24680 15264 25000 16288
rect 24680 15200 24688 15264
rect 24752 15200 24768 15264
rect 24832 15200 24848 15264
rect 24912 15200 24928 15264
rect 24992 15200 25000 15264
rect 24680 14176 25000 15200
rect 24680 14112 24688 14176
rect 24752 14112 24768 14176
rect 24832 14112 24848 14176
rect 24912 14112 24928 14176
rect 24992 14112 25000 14176
rect 24680 13088 25000 14112
rect 24680 13024 24688 13088
rect 24752 13024 24768 13088
rect 24832 13024 24848 13088
rect 24912 13024 24928 13088
rect 24992 13024 25000 13088
rect 24680 12000 25000 13024
rect 24680 11936 24688 12000
rect 24752 11936 24768 12000
rect 24832 11936 24848 12000
rect 24912 11936 24928 12000
rect 24992 11936 25000 12000
rect 24680 10912 25000 11936
rect 24680 10848 24688 10912
rect 24752 10848 24768 10912
rect 24832 10848 24848 10912
rect 24912 10848 24928 10912
rect 24992 10848 25000 10912
rect 24680 9824 25000 10848
rect 24680 9760 24688 9824
rect 24752 9760 24768 9824
rect 24832 9760 24848 9824
rect 24912 9760 24928 9824
rect 24992 9760 25000 9824
rect 24680 8736 25000 9760
rect 24680 8672 24688 8736
rect 24752 8672 24768 8736
rect 24832 8672 24848 8736
rect 24912 8672 24928 8736
rect 24992 8672 25000 8736
rect 24680 7648 25000 8672
rect 24680 7584 24688 7648
rect 24752 7584 24768 7648
rect 24832 7584 24848 7648
rect 24912 7584 24928 7648
rect 24992 7584 25000 7648
rect 24680 6560 25000 7584
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 22691 5540 22757 5541
rect 22691 5476 22692 5540
rect 22756 5476 22757 5540
rect 22691 5475 22757 5476
rect 22875 5540 22941 5541
rect 22875 5476 22876 5540
rect 22940 5476 22941 5540
rect 22875 5475 22941 5476
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 22139 3228 22205 3229
rect 22139 3164 22140 3228
rect 22204 3164 22205 3228
rect 22139 3163 22205 3164
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 20667 2004 20733 2005
rect 20667 1940 20668 2004
rect 20732 1940 20733 2004
rect 20667 1939 20733 1940
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 21713 1040 22033 1600
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
use sky130_fd_sc_hd__clkbuf_1  _000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _001_
timestamp 1688980957
transform 1 0 23276 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp 1688980957
transform 1 0 23184 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp 1688980957
transform 1 0 23184 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _004_
timestamp 1688980957
transform 1 0 23368 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp 1688980957
transform 1 0 23276 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp 1688980957
transform 1 0 23920 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp 1688980957
transform 1 0 22816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp 1688980957
transform 1 0 23552 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _009_
timestamp 1688980957
transform 1 0 21620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp 1688980957
transform 1 0 23092 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp 1688980957
transform 1 0 23644 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp 1688980957
transform 1 0 23092 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp 1688980957
transform 1 0 23736 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _015_
timestamp 1688980957
transform 1 0 20792 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _016_
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp 1688980957
transform 1 0 22816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _018_
timestamp 1688980957
transform 1 0 22356 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp 1688980957
transform 1 0 20608 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp 1688980957
transform 1 0 21620 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp 1688980957
transform 1 0 23368 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp 1688980957
transform 1 0 23644 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp 1688980957
transform 1 0 19780 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp 1688980957
transform 1 0 20056 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp 1688980957
transform 1 0 23460 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp 1688980957
transform 1 0 21160 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1688980957
transform 1 0 21344 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform 1 0 22356 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 20240 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1688980957
transform 1 0 20516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1688980957
transform 1 0 20332 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 23000 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 22080 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 20792 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1688980957
transform 1 0 17296 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1688980957
transform 1 0 22356 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 21160 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 21620 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform 1 0 21068 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform 1 0 20884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 22080 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1688980957
transform 1 0 20608 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1688980957
transform 1 0 23092 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1688980957
transform 1 0 12696 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp 1688980957
transform 1 0 15272 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 8372 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 3036 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 2760 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 3404 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 2852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 4416 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 4692 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 5428 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 6164 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 5152 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 5796 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 7176 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 7544 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 7820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 8096 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 10580 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 13340 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 11592 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 12420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 18308 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 18584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 16744 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform 1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 5336 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1688980957
transform 1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 7084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 3036 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 1472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1688980957
transform 1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1688980957
transform 1 0 1472 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1688980957
transform 1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1688980957
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 3036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 1472 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 5428 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform 1 0 3220 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform 1 0 3220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1688980957
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 4324 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 6992 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 23552 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 4508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 5336 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 5888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 7636 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 22724 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 23092 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 23184 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 23460 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 23092 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 22264 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 22632 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 18768 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 20976 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 18952 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 20056 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 22816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 21896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 19872 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 22080 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 22448 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 19320 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 20608 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 23184 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 23552 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 23736 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 23460 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 23460 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 23644 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 23552 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 23736 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 23460 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 21160 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 23368 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 22816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 23368 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 23184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 19872 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 23092 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 21620 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 19596 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 23644 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 23000 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 20424 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 22816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 20884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 20240 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 19964 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 21160 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 20332 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_39
timestamp 1688980957
transform 1 0 4692 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_61
timestamp 1688980957
transform 1 0 6716 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_75
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_21
timestamp 1688980957
transform 1 0 3036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_139
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_253
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_11
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_42 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_88
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_129
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_159
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_163
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_234
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_19 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_34
timestamp 1688980957
transform 1 0 4232 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_116
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_135
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_159
timestamp 1688980957
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_20
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_37
timestamp 1688980957
transform 1 0 4508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_64
timestamp 1688980957
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_106
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_114
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_156
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_168
timestamp 1688980957
transform 1 0 16560 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_180
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_38
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_50
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_128
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_183
timestamp 1688980957
transform 1 0 17940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_199
timestamp 1688980957
transform 1 0 19412 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_250
timestamp 1688980957
transform 1 0 24104 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_35
timestamp 1688980957
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_52
timestamp 1688980957
transform 1 0 5888 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_64
timestamp 1688980957
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_170
timestamp 1688980957
transform 1 0 16744 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_230
timestamp 1688980957
transform 1 0 22264 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_72
timestamp 1688980957
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_84
timestamp 1688980957
transform 1 0 8832 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_103
timestamp 1688980957
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_14
timestamp 1688980957
transform 1 0 2392 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_52
timestamp 1688980957
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_125
timestamp 1688980957
transform 1 0 12604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 1688980957
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_212
timestamp 1688980957
transform 1 0 20608 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_238
timestamp 1688980957
transform 1 0 23000 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_29
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_165
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_177
timestamp 1688980957
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_184
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_196
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_208
timestamp 1688980957
transform 1 0 20240 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_11
timestamp 1688980957
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_35
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_52
timestamp 1688980957
transform 1 0 5888 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_64
timestamp 1688980957
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_76
timestamp 1688980957
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_118
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_238
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1688980957
transform 1 0 23736 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_129
timestamp 1688980957
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 1688980957
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_201
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_228
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_245
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_35
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_190
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_207
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_229
timestamp 1688980957
transform 1 0 22172 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_83
timestamp 1688980957
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_131
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_135
timestamp 1688980957
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_238
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_35
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_47
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_59
timestamp 1688980957
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_67
timestamp 1688980957
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_186
timestamp 1688980957
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 1688980957
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_217
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_24
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_143
timestamp 1688980957
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_218
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_234
timestamp 1688980957
transform 1 0 22632 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_253
timestamp 1688980957
transform 1 0 24380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_71
timestamp 1688980957
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_129
timestamp 1688980957
transform 1 0 12972 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_180
timestamp 1688980957
transform 1 0 17664 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_186
timestamp 1688980957
transform 1 0 18216 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_190
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_205
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_229
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_250
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_72
timestamp 1688980957
transform 1 0 7728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_84
timestamp 1688980957
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_103
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_108
timestamp 1688980957
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_152
timestamp 1688980957
transform 1 0 15088 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 1688980957
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_177
timestamp 1688980957
transform 1 0 17388 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_231
timestamp 1688980957
transform 1 0 22356 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_250
timestamp 1688980957
transform 1 0 24104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_254
timestamp 1688980957
transform 1 0 24472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_17
timestamp 1688980957
transform 1 0 2668 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_58
timestamp 1688980957
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_106
timestamp 1688980957
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_118
timestamp 1688980957
transform 1 0 11960 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_200
timestamp 1688980957
transform 1 0 19504 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_217
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_229
timestamp 1688980957
transform 1 0 22172 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_7
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_143
timestamp 1688980957
transform 1 0 14260 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_199
timestamp 1688980957
transform 1 0 19412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_211
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_219
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_238
timestamp 1688980957
transform 1 0 23000 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_129
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_159
timestamp 1688980957
transform 1 0 15732 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_203
timestamp 1688980957
transform 1 0 19780 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_49
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_72
timestamp 1688980957
transform 1 0 7728 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_130
timestamp 1688980957
transform 1 0 13064 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_154
timestamp 1688980957
transform 1 0 15272 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_185
timestamp 1688980957
transform 1 0 18124 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_246
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_253
timestamp 1688980957
transform 1 0 24380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_44
timestamp 1688980957
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_56
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_68
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_80
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_92
timestamp 1688980957
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_123
timestamp 1688980957
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_183
timestamp 1688980957
transform 1 0 17940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_193
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_61
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_162
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_202
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_214
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_248
timestamp 1688980957
transform 1 0 23920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_39
timestamp 1688980957
transform 1 0 4692 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_218
timestamp 1688980957
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_224
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_50
timestamp 1688980957
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_86
timestamp 1688980957
transform 1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_131
timestamp 1688980957
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_154
timestamp 1688980957
transform 1 0 15272 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_190
timestamp 1688980957
transform 1 0 18584 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_198
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_240
timestamp 1688980957
transform 1 0 23184 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_44
timestamp 1688980957
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_185
timestamp 1688980957
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_190
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_212
timestamp 1688980957
transform 1 0 20608 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_224
timestamp 1688980957
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_99
timestamp 1688980957
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_134
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_142
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_159
timestamp 1688980957
transform 1 0 15732 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_204
timestamp 1688980957
transform 1 0 19872 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_215
timestamp 1688980957
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_253
timestamp 1688980957
transform 1 0 24380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_35
timestamp 1688980957
transform 1 0 4324 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_183
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_222
timestamp 1688980957
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_230
timestamp 1688980957
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_250
timestamp 1688980957
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_30
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_38
timestamp 1688980957
transform 1 0 4600 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_75
timestamp 1688980957
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_87
timestamp 1688980957
transform 1 0 9108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_95
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_124
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_184
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_196
timestamp 1688980957
transform 1 0 19136 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_203
timestamp 1688980957
transform 1 0 19780 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_209
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_214
timestamp 1688980957
transform 1 0 20792 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_219
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_240
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_50
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_69
timestamp 1688980957
transform 1 0 7452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_118
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_156
timestamp 1688980957
transform 1 0 15456 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_168
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_192
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_29
timestamp 1688980957
transform 1 0 3772 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_131
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_139
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_173
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_207
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_219
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_24
timestamp 1688980957
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_44
timestamp 1688980957
transform 1 0 5152 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_56
timestamp 1688980957
transform 1 0 6256 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_64
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_80
timestamp 1688980957
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_137
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_204
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_208
timestamp 1688980957
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_220
timestamp 1688980957
transform 1 0 21344 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_232
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_241
timestamp 1688980957
transform 1 0 23276 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_128
timestamp 1688980957
transform 1 0 12880 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_184
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_235
timestamp 1688980957
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_239
timestamp 1688980957
transform 1 0 23092 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_32
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_78
timestamp 1688980957
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_113
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_250
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_18
timestamp 1688980957
transform 1 0 2760 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_143
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_159
timestamp 1688980957
transform 1 0 15732 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_196
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_208
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_220
timestamp 1688980957
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_254
timestamp 1688980957
transform 1 0 24472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_68
timestamp 1688980957
transform 1 0 7360 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_115
timestamp 1688980957
transform 1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_147
timestamp 1688980957
transform 1 0 14628 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_169
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_187
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_200
timestamp 1688980957
transform 1 0 19504 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_208
timestamp 1688980957
transform 1 0 20240 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_212
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_216
timestamp 1688980957
transform 1 0 20976 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_228
timestamp 1688980957
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_232
timestamp 1688980957
transform 1 0 22448 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_24
timestamp 1688980957
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_36
timestamp 1688980957
transform 1 0 4416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_54
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_75
timestamp 1688980957
transform 1 0 8004 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_96
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_131
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_147
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_196
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_200
timestamp 1688980957
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_228
timestamp 1688980957
transform 1 0 22080 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_240
timestamp 1688980957
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_32
timestamp 1688980957
transform 1 0 4048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_36
timestamp 1688980957
transform 1 0 4416 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_55
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_75
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17664 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_213
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_217
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_225
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_234
timestamp 1688980957
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_238
timestamp 1688980957
transform 1 0 23000 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_48
timestamp 1688980957
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_72
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_80
timestamp 1688980957
transform 1 0 8464 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_150
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_190
timestamp 1688980957
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_214
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_220
timestamp 1688980957
transform 1 0 21344 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_24
timestamp 1688980957
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_78
timestamp 1688980957
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_99
timestamp 1688980957
transform 1 0 10212 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_119
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_131
timestamp 1688980957
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_168
timestamp 1688980957
transform 1 0 16560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_180
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_191
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_200
timestamp 1688980957
transform 1 0 19504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_205
timestamp 1688980957
transform 1 0 19964 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_211
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_247
timestamp 1688980957
transform 1 0 23828 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_13
timestamp 1688980957
transform 1 0 2300 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_33
timestamp 1688980957
transform 1 0 4140 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_120
timestamp 1688980957
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_124
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_146
timestamp 1688980957
transform 1 0 14536 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_233
timestamp 1688980957
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_239
timestamp 1688980957
transform 1 0 23092 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_21
timestamp 1688980957
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_68
timestamp 1688980957
transform 1 0 7360 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_75
timestamp 1688980957
transform 1 0 8004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_118
timestamp 1688980957
transform 1 0 11960 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_124
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_187
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_206
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_212
timestamp 1688980957
transform 1 0 20608 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_218
timestamp 1688980957
transform 1 0 21160 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_230
timestamp 1688980957
transform 1 0 22264 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_77
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_95
timestamp 1688980957
transform 1 0 9844 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_159
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_199
timestamp 1688980957
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_203
timestamp 1688980957
transform 1 0 19780 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_228
timestamp 1688980957
transform 1 0 22080 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_247
timestamp 1688980957
transform 1 0 23828 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_12
timestamp 1688980957
transform 1 0 2208 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_62
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_66
timestamp 1688980957
transform 1 0 7176 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_82
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_128
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_200
timestamp 1688980957
transform 1 0 19504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_204
timestamp 1688980957
transform 1 0 19872 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_208
timestamp 1688980957
transform 1 0 20240 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_224
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_241
timestamp 1688980957
transform 1 0 23276 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_107
timestamp 1688980957
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_128
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_151
timestamp 1688980957
transform 1 0 14996 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_234
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_241
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_32
timestamp 1688980957
transform 1 0 4048 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_44
timestamp 1688980957
transform 1 0 5152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_56
timestamp 1688980957
transform 1 0 6256 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_74
timestamp 1688980957
transform 1 0 7912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_82
timestamp 1688980957
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_129
timestamp 1688980957
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_172
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_200
timestamp 1688980957
transform 1 0 19504 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_224
timestamp 1688980957
transform 1 0 21712 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_232
timestamp 1688980957
transform 1 0 22448 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_238
timestamp 1688980957
transform 1 0 23000 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_242
timestamp 1688980957
transform 1 0 23368 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_7
timestamp 1688980957
transform 1 0 1748 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_29
timestamp 1688980957
transform 1 0 3772 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_52
timestamp 1688980957
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_87
timestamp 1688980957
transform 1 0 9108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_99
timestamp 1688980957
transform 1 0 10212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1688980957
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_190
timestamp 1688980957
transform 1 0 18584 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_202
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_214
timestamp 1688980957
transform 1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_240
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_247
timestamp 1688980957
transform 1 0 23828 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_21
timestamp 1688980957
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_73
timestamp 1688980957
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_103
timestamp 1688980957
transform 1 0 10580 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_111
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_128
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_149
timestamp 1688980957
transform 1 0 14812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_154
timestamp 1688980957
transform 1 0 15272 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_162
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_208
timestamp 1688980957
transform 1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_214
timestamp 1688980957
transform 1 0 20792 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_247
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_34
timestamp 1688980957
transform 1 0 4232 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1688980957
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_72
timestamp 1688980957
transform 1 0 7728 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_84
timestamp 1688980957
transform 1 0 8832 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_96
timestamp 1688980957
transform 1 0 9936 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_148
timestamp 1688980957
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_152
timestamp 1688980957
transform 1 0 15088 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_198
timestamp 1688980957
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_231
timestamp 1688980957
transform 1 0 22356 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_45
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_57
timestamp 1688980957
transform 1 0 6348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_100
timestamp 1688980957
transform 1 0 10304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_114
timestamp 1688980957
transform 1 0 11592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_130
timestamp 1688980957
transform 1 0 13064 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_156
timestamp 1688980957
transform 1 0 15456 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_183
timestamp 1688980957
transform 1 0 17940 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_187
timestamp 1688980957
transform 1 0 18308 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_191
timestamp 1688980957
transform 1 0 18676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_200
timestamp 1688980957
transform 1 0 19504 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_220
timestamp 1688980957
transform 1 0 21344 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_232
timestamp 1688980957
transform 1 0 22448 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_246
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_11
timestamp 1688980957
transform 1 0 2116 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_30
timestamp 1688980957
transform 1 0 3864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_38
timestamp 1688980957
transform 1 0 4600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_83
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_87
timestamp 1688980957
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_117
timestamp 1688980957
transform 1 0 11868 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_123
timestamp 1688980957
transform 1 0 12420 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_139
timestamp 1688980957
transform 1 0 13892 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_159
timestamp 1688980957
transform 1 0 15732 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_184
timestamp 1688980957
transform 1 0 18032 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_192
timestamp 1688980957
transform 1 0 18768 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_211
timestamp 1688980957
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_248
timestamp 1688980957
transform 1 0 23920 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_39
timestamp 1688980957
transform 1 0 4692 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_58
timestamp 1688980957
transform 1 0 6440 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_62
timestamp 1688980957
transform 1 0 6808 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_101
timestamp 1688980957
transform 1 0 10396 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_178
timestamp 1688980957
transform 1 0 17480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_190
timestamp 1688980957
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_215
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_226
timestamp 1688980957
transform 1 0 21896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_234
timestamp 1688980957
transform 1 0 22632 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_240
timestamp 1688980957
transform 1 0 23184 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_247
timestamp 1688980957
transform 1 0 23828 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_31
timestamp 1688980957
transform 1 0 3956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_48
timestamp 1688980957
transform 1 0 5520 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_61
timestamp 1688980957
transform 1 0 6716 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_77
timestamp 1688980957
transform 1 0 8188 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_89
timestamp 1688980957
transform 1 0 9292 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_95
timestamp 1688980957
transform 1 0 9844 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_154
timestamp 1688980957
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 1688980957
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_198
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_7
timestamp 1688980957
transform 1 0 1748 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_32
timestamp 1688980957
transform 1 0 4048 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_49
timestamp 1688980957
transform 1 0 5612 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 1688980957
transform 1 0 7728 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_100
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_154
timestamp 1688980957
transform 1 0 15272 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_158
timestamp 1688980957
transform 1 0 15640 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_207
timestamp 1688980957
transform 1 0 20148 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_211
timestamp 1688980957
transform 1 0 20516 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_215
timestamp 1688980957
transform 1 0 20884 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_227
timestamp 1688980957
transform 1 0 21988 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_231
timestamp 1688980957
transform 1 0 22356 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_235
timestamp 1688980957
transform 1 0 22724 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_242
timestamp 1688980957
transform 1 0 23368 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_49
timestamp 1688980957
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_75
timestamp 1688980957
transform 1 0 8004 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_79
timestamp 1688980957
transform 1 0 8372 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_98
timestamp 1688980957
transform 1 0 10120 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_117
timestamp 1688980957
transform 1 0 11868 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_142
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_150
timestamp 1688980957
transform 1 0 14904 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_187
timestamp 1688980957
transform 1 0 18308 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_192
timestamp 1688980957
transform 1 0 18768 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_222
timestamp 1688980957
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_229
timestamp 1688980957
transform 1 0 22172 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_233
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_240
timestamp 1688980957
transform 1 0 23184 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_247
timestamp 1688980957
transform 1 0 23828 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_24
timestamp 1688980957
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_42
timestamp 1688980957
transform 1 0 4968 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_50
timestamp 1688980957
transform 1 0 5704 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_66
timestamp 1688980957
transform 1 0 7176 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_78
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_105
timestamp 1688980957
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_156
timestamp 1688980957
transform 1 0 15456 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_178
timestamp 1688980957
transform 1 0 17480 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_190
timestamp 1688980957
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_203
timestamp 1688980957
transform 1 0 19780 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_226
timestamp 1688980957
transform 1 0 21896 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_238
timestamp 1688980957
transform 1 0 23000 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_242
timestamp 1688980957
transform 1 0 23368 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_41
timestamp 1688980957
transform 1 0 4876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_53
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_90
timestamp 1688980957
transform 1 0 9384 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_96
timestamp 1688980957
transform 1 0 9936 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_157
timestamp 1688980957
transform 1 0 15548 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_165
timestamp 1688980957
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_212
timestamp 1688980957
transform 1 0 20608 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_228
timestamp 1688980957
transform 1 0 22080 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_9
timestamp 1688980957
transform 1 0 1932 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_38
timestamp 1688980957
transform 1 0 4600 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_58
timestamp 1688980957
transform 1 0 6440 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_93
timestamp 1688980957
transform 1 0 9660 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_132
timestamp 1688980957
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_162
timestamp 1688980957
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_174
timestamp 1688980957
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_178
timestamp 1688980957
transform 1 0 17480 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_194
timestamp 1688980957
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_225
timestamp 1688980957
transform 1 0 21804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_232
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_239
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_37
timestamp 1688980957
transform 1 0 4508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_90
timestamp 1688980957
transform 1 0 9384 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_106
timestamp 1688980957
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_201
timestamp 1688980957
transform 1 0 19596 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_248
timestamp 1688980957
transform 1 0 23920 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_24
timestamp 1688980957
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_52
timestamp 1688980957
transform 1 0 5888 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_60
timestamp 1688980957
transform 1 0 6624 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_100
timestamp 1688980957
transform 1 0 10304 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_112
timestamp 1688980957
transform 1 0 11408 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_156
timestamp 1688980957
transform 1 0 15456 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_160
timestamp 1688980957
transform 1 0 15824 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_179
timestamp 1688980957
transform 1 0 17572 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_183
timestamp 1688980957
transform 1 0 17940 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_188
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_223
timestamp 1688980957
transform 1 0 21620 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_237
timestamp 1688980957
transform 1 0 22908 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_24
timestamp 1688980957
transform 1 0 3312 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_72
timestamp 1688980957
transform 1 0 7728 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_80
timestamp 1688980957
transform 1 0 8464 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_87
timestamp 1688980957
transform 1 0 9108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_141
timestamp 1688980957
transform 1 0 14076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_157
timestamp 1688980957
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_165
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_179
timestamp 1688980957
transform 1 0 17572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_191
timestamp 1688980957
transform 1 0 18676 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_243
timestamp 1688980957
transform 1 0 23460 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_248
timestamp 1688980957
transform 1 0 23920 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_9
timestamp 1688980957
transform 1 0 1932 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_62
timestamp 1688980957
transform 1 0 6808 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_74
timestamp 1688980957
transform 1 0 7912 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_93
timestamp 1688980957
transform 1 0 9660 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_131
timestamp 1688980957
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_156
timestamp 1688980957
transform 1 0 15456 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_173
timestamp 1688980957
transform 1 0 17020 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_188
timestamp 1688980957
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_203
timestamp 1688980957
transform 1 0 19780 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_207
timestamp 1688980957
transform 1 0 20148 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_213
timestamp 1688980957
transform 1 0 20700 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_217
timestamp 1688980957
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_229
timestamp 1688980957
transform 1 0 22172 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_246
timestamp 1688980957
transform 1 0 23736 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_31
timestamp 1688980957
transform 1 0 3956 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_73
timestamp 1688980957
transform 1 0 7820 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_108
timestamp 1688980957
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_146
timestamp 1688980957
transform 1 0 14536 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_158
timestamp 1688980957
transform 1 0 15640 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_166
timestamp 1688980957
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_177
timestamp 1688980957
transform 1 0 17388 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_201
timestamp 1688980957
transform 1 0 19596 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_213
timestamp 1688980957
transform 1 0 20700 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_220
timestamp 1688980957
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_228
timestamp 1688980957
transform 1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_242
timestamp 1688980957
transform 1 0 23368 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_25
timestamp 1688980957
transform 1 0 3404 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_67
timestamp 1688980957
transform 1 0 7268 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_79
timestamp 1688980957
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_173
timestamp 1688980957
transform 1 0 17020 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_215
timestamp 1688980957
transform 1 0 20884 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_219
timestamp 1688980957
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_226
timestamp 1688980957
transform 1 0 21896 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_230
timestamp 1688980957
transform 1 0 22264 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_234
timestamp 1688980957
transform 1 0 22632 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_96
timestamp 1688980957
transform 1 0 9936 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_108
timestamp 1688980957
transform 1 0 11040 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_128
timestamp 1688980957
transform 1 0 12880 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_140
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_152
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_164
timestamp 1688980957
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_177
timestamp 1688980957
transform 1 0 17388 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_182
timestamp 1688980957
transform 1 0 17848 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_197
timestamp 1688980957
transform 1 0 19228 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_204
timestamp 1688980957
transform 1 0 19872 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_218
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_233
timestamp 1688980957
transform 1 0 22540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_242
timestamp 1688980957
transform 1 0 23368 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_246
timestamp 1688980957
transform 1 0 23736 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_14
timestamp 1688980957
transform 1 0 2392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_35
timestamp 1688980957
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_54
timestamp 1688980957
transform 1 0 6072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_58
timestamp 1688980957
transform 1 0 6440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_81
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_124
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_136
timestamp 1688980957
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_214
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_222
timestamp 1688980957
transform 1 0 21528 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_229
timestamp 1688980957
transform 1 0 22172 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_54
timestamp 1688980957
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_72
timestamp 1688980957
transform 1 0 7728 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_80
timestamp 1688980957
transform 1 0 8464 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_101
timestamp 1688980957
transform 1 0 10396 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_109
timestamp 1688980957
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_134
timestamp 1688980957
transform 1 0 13432 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_146
timestamp 1688980957
transform 1 0 14536 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_158
timestamp 1688980957
transform 1 0 15640 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_166
timestamp 1688980957
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_250
timestamp 1688980957
transform 1 0 24104 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_25
timestamp 1688980957
transform 1 0 3404 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_44
timestamp 1688980957
transform 1 0 5152 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_67
timestamp 1688980957
transform 1 0 7268 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_79
timestamp 1688980957
transform 1 0 8372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_102
timestamp 1688980957
transform 1 0 10488 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_110
timestamp 1688980957
transform 1 0 11224 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_203
timestamp 1688980957
transform 1 0 19780 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_207
timestamp 1688980957
transform 1 0 20148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_219
timestamp 1688980957
transform 1 0 21252 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_227
timestamp 1688980957
transform 1 0 21988 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_231
timestamp 1688980957
transform 1 0 22356 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_244
timestamp 1688980957
transform 1 0 23552 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_75
timestamp 1688980957
transform 1 0 8004 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_91
timestamp 1688980957
transform 1 0 9476 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_103
timestamp 1688980957
transform 1 0 10580 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_128
timestamp 1688980957
transform 1 0 12880 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_140
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_152
timestamp 1688980957
transform 1 0 15088 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_164
timestamp 1688980957
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_209
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_216
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_220
timestamp 1688980957
transform 1 0 21344 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_241
timestamp 1688980957
transform 1 0 23276 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_248
timestamp 1688980957
transform 1 0 23920 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_25
timestamp 1688980957
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_118
timestamp 1688980957
transform 1 0 11960 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_137
timestamp 1688980957
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_216
timestamp 1688980957
transform 1 0 20976 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_220
timestamp 1688980957
transform 1 0 21344 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_234
timestamp 1688980957
transform 1 0 22632 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_239
timestamp 1688980957
transform 1 0 23092 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_243
timestamp 1688980957
transform 1 0 23460 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_33
timestamp 1688980957
transform 1 0 4140 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_37
timestamp 1688980957
transform 1 0 4508 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_65
timestamp 1688980957
transform 1 0 7084 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_103
timestamp 1688980957
transform 1 0 10580 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_109
timestamp 1688980957
transform 1 0 11132 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71_200
timestamp 1688980957
transform 1 0 19504 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_243
timestamp 1688980957
transform 1 0 23460 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_248
timestamp 1688980957
transform 1 0 23920 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_44
timestamp 1688980957
transform 1 0 5152 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_78
timestamp 1688980957
transform 1 0 8280 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_93
timestamp 1688980957
transform 1 0 9660 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_134
timestamp 1688980957
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_204
timestamp 1688980957
transform 1 0 19872 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_241
timestamp 1688980957
transform 1 0 23276 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_14
timestamp 1688980957
transform 1 0 2392 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_24
timestamp 1688980957
transform 1 0 3312 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_75
timestamp 1688980957
transform 1 0 8004 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_96
timestamp 1688980957
transform 1 0 9936 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_198
timestamp 1688980957
transform 1 0 19320 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_234
timestamp 1688980957
transform 1 0 22632 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_253
timestamp 1688980957
transform 1 0 24380 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_35
timestamp 1688980957
transform 1 0 4324 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_42
timestamp 1688980957
transform 1 0 4968 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_50
timestamp 1688980957
transform 1 0 5704 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_54
timestamp 1688980957
transform 1 0 6072 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_58
timestamp 1688980957
transform 1 0 6440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_62
timestamp 1688980957
transform 1 0 6808 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_69
timestamp 1688980957
transform 1 0 7452 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_82
timestamp 1688980957
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_108
timestamp 1688980957
transform 1 0 11040 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_120
timestamp 1688980957
transform 1 0 12144 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_132
timestamp 1688980957
transform 1 0 13248 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_190
timestamp 1688980957
transform 1 0 18584 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_204
timestamp 1688980957
transform 1 0 19872 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_214
timestamp 1688980957
transform 1 0 20792 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_227
timestamp 1688980957
transform 1 0 21988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_22
timestamp 1688980957
transform 1 0 3128 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_35
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_44
timestamp 1688980957
transform 1 0 5152 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_48
timestamp 1688980957
transform 1 0 5520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_60
timestamp 1688980957
transform 1 0 6624 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_84
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_91
timestamp 1688980957
transform 1 0 9476 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_99
timestamp 1688980957
transform 1 0 10212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_201
timestamp 1688980957
transform 1 0 19596 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_228
timestamp 1688980957
transform 1 0 22080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_247
timestamp 1688980957
transform 1 0 23828 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_254
timestamp 1688980957
transform 1 0 24472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_9
timestamp 1688980957
transform 1 0 1932 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_58
timestamp 1688980957
transform 1 0 6440 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_76
timestamp 1688980957
transform 1 0 8096 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_88
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_96
timestamp 1688980957
transform 1 0 9936 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_106
timestamp 1688980957
transform 1 0 10856 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_132
timestamp 1688980957
transform 1 0 13248 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_150
timestamp 1688980957
transform 1 0 14904 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_160
timestamp 1688980957
transform 1 0 15824 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_164
timestamp 1688980957
transform 1 0 16192 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_220
timestamp 1688980957
transform 1 0 21344 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_12
timestamp 1688980957
transform 1 0 2208 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_26
timestamp 1688980957
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_32
timestamp 1688980957
transform 1 0 4048 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_42
timestamp 1688980957
transform 1 0 4968 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_50
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_85
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_117
timestamp 1688980957
transform 1 0 11868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_130
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_145
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_155
timestamp 1688980957
transform 1 0 15364 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_173
timestamp 1688980957
transform 1 0 17020 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_194
timestamp 1688980957
transform 1 0 18952 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_203
timestamp 1688980957
transform 1 0 19780 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_247
timestamp 1688980957
transform 1 0 23828 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_253
timestamp 1688980957
transform 1 0 24380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform 1 0 3404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 2944 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 2300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 3220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 2760 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 2576 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 3680 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1688980957
transform 1 0 2760 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1688980957
transform 1 0 3036 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 3404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1748 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2760 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 2300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 2024 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 2208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 2944 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 3220 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input50
timestamp 1688980957
transform 1 0 2852 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input51
timestamp 1688980957
transform 1 0 3404 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 4876 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input54
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 3312 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 4968 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 5520 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1688980957
transform 1 0 4048 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input66 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input67
timestamp 1688980957
transform 1 0 2392 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input68
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input69
timestamp 1688980957
transform 1 0 4600 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input70
timestamp 1688980957
transform 1 0 2392 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input71
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input72
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input73
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 3312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input75
timestamp 1688980957
transform 1 0 3864 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input76
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1688980957
transform 1 0 2760 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input78
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 2760 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input80
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 21252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 18032 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input88
timestamp 1688980957
transform 1 0 24196 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1688980957
transform 1 0 18584 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1688980957
transform 1 0 21068 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input92
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input93
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input95
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input97
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 23000 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input103
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input104
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1688980957
transform 1 0 3496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input106
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input107
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1688980957
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1688980957
transform 1 0 4784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1688980957
transform 1 0 5244 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input119
timestamp 1688980957
transform 1 0 3036 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input128
timestamp 1688980957
transform 1 0 5336 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input129
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 5060 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 22724 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 21528 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1688980957
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1688980957
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1688980957
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 9936 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 10304 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1688980957
transform 1 0 10672 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1688980957
transform 1 0 11040 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input157
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1688980957
transform 1 0 11592 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1688980957
transform 1 0 11868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1688980957
transform 1 0 12328 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1688980957
transform 1 0 12696 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1688980957
transform 1 0 13616 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 14628 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 14352 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input169
timestamp 1688980957
transform 1 0 14628 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1688980957
transform 1 0 14996 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1688980957
transform 1 0 15548 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1688980957
transform 1 0 15456 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input173
timestamp 1688980957
transform 1 0 15824 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 20792 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 18768 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 19596 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 20516 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 19504 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 17940 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 16192 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input181
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input182
timestamp 1688980957
transform 1 0 16560 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 17572 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 17848 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 18124 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 18400 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 21068 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._0_
timestamp 1688980957
transform 1 0 24104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._1_
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._2_
timestamp 1688980957
transform 1 0 22448 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._3_
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22172 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 24288 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23000 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22448 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 22080 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21160 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22356 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 24196 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22448 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23184 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19596 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20240 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19136 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21804 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20056 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 20608 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20884 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22080 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22724 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23184 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21160 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20240 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19412 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17112 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17848 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 21620 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21988 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20976 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22080 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18124 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19320 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18952 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17572 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20240 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18400 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20608 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 22080 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 21436 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23000 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23460 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23368 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22356 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18124 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19320 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21160 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19044 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23000 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23276 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22080 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22632 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20516 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 21344 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20976 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19504 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20792 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18492 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19596 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19872 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19872 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19780 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19596 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19504 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23184 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22172 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23276 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22632 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 20148 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19688 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21252 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20700 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 20608 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19872 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 21252 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 23092 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 21528 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22724 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23000 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23276 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 22172 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 23092 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22356 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19596 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18952 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17480 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17664 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 23000 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 23368 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 22632 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 23736 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 12512 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 2300 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 4232 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 4876 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 5060 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 6072 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 1656 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 1932 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 9660 0 1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 12604 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 12052 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 1472 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 2300 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 11776 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 12328 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 17112 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 9936 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 2300 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 3496 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 8096 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 9108 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 11684 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 1840 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 4876 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 12880 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 13892 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 10856 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 3496 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 6900 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 10028 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 11684 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 4508 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 10028 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 15088 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 12604 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 3404 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 11868 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 12512 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 18032 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 16008 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 14628 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 6624 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 7268 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit0
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit2
timestamp 1688980957
transform 1 0 6624 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit3
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit4
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit5
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit6
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit7
timestamp 1688980957
transform 1 0 9200 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit8
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit10
timestamp 1688980957
transform 1 0 6808 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit11
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit12
timestamp 1688980957
transform 1 0 2300 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit13
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 11500 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 2208 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 2300 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 15180 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 12420 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 16192 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 17572 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit0
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit1
timestamp 1688980957
transform 1 0 17112 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit3
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit4
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit5
timestamp 1688980957
transform 1 0 3496 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit6
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit7
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit8
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit9
timestamp 1688980957
transform 1 0 16744 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit11
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit12
timestamp 1688980957
transform 1 0 1656 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit13
timestamp 1688980957
transform 1 0 2024 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit14
timestamp 1688980957
transform 1 0 6808 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit15
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit16
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit17
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit18
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit19
timestamp 1688980957
transform 1 0 6808 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit20
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit21
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit22
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit23
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit24
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit25
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit26
timestamp 1688980957
transform 1 0 4876 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit27
timestamp 1688980957
transform 1 0 5520 0 1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit28
timestamp 1688980957
transform 1 0 4876 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit29
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit30
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12604 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit0
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit2
timestamp 1688980957
transform 1 0 1840 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit3
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit5
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit6
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit7
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit8
timestamp 1688980957
transform 1 0 7452 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit9
timestamp 1688980957
transform 1 0 9200 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit10
timestamp 1688980957
transform 1 0 3956 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit11
timestamp 1688980957
transform 1 0 4508 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit12
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit13
timestamp 1688980957
transform 1 0 1564 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit14
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit15
timestamp 1688980957
transform 1 0 6440 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit16
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit17
timestamp 1688980957
transform 1 0 15364 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1840 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit19
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1656 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit21
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit22
timestamp 1688980957
transform 1 0 6716 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit23
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit24
timestamp 1688980957
transform 1 0 17204 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit25
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit26
timestamp 1688980957
transform 1 0 4324 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit27
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit28
timestamp 1688980957
transform 1 0 1656 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit29
timestamp 1688980957
transform 1 0 2208 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit30
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit31
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit0
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit1
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit2
timestamp 1688980957
transform 1 0 13432 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit3
timestamp 1688980957
transform 1 0 14168 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit4
timestamp 1688980957
transform 1 0 12512 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit6
timestamp 1688980957
transform 1 0 14904 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit7
timestamp 1688980957
transform 1 0 4784 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit8
timestamp 1688980957
transform 1 0 5428 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit9
timestamp 1688980957
transform 1 0 6900 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit10
timestamp 1688980957
transform 1 0 9936 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit11
timestamp 1688980957
transform 1 0 11040 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit12
timestamp 1688980957
transform 1 0 12512 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit13
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit14
timestamp 1688980957
transform 1 0 16928 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit15
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit16
timestamp 1688980957
transform 1 0 9844 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit17
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit18
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit19
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit20
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit21
timestamp 1688980957
transform 1 0 9200 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit22
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit23
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit24
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit25
timestamp 1688980957
transform 1 0 9384 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit26
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit27
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit28
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit29
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit30
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit31
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit0
timestamp 1688980957
transform 1 0 8464 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit1
timestamp 1688980957
transform 1 0 9476 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit2
timestamp 1688980957
transform 1 0 9200 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit3
timestamp 1688980957
transform 1 0 4692 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit4
timestamp 1688980957
transform 1 0 5428 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit5
timestamp 1688980957
transform 1 0 6532 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit6
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit7
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit8
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit9
timestamp 1688980957
transform 1 0 15180 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit10
timestamp 1688980957
transform 1 0 15916 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit11
timestamp 1688980957
transform 1 0 15640 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit12
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit13
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit14
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit15
timestamp 1688980957
transform 1 0 4876 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit16
timestamp 1688980957
transform 1 0 11776 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit17
timestamp 1688980957
transform 1 0 13156 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit18
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit19
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit20
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit21
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit22
timestamp 1688980957
transform 1 0 4784 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit23
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit24
timestamp 1688980957
transform 1 0 5796 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit25
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit26
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit27
timestamp 1688980957
transform 1 0 14168 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit28
timestamp 1688980957
transform 1 0 11960 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit29
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit30
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit31
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit0
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit1
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit2
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit3
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit4
timestamp 1688980957
transform 1 0 22724 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit5
timestamp 1688980957
transform 1 0 22724 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit6
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit7
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit8
timestamp 1688980957
transform 1 0 7728 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit9
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1472 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit12
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit13
timestamp 1688980957
transform 1 0 12052 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit14
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit15
timestamp 1688980957
transform 1 0 14168 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit16
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit17
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1656 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit22
timestamp 1688980957
transform 1 0 6808 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit23
timestamp 1688980957
transform 1 0 7360 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit24
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit25
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit26
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit27
timestamp 1688980957
transform 1 0 1472 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1564 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit30
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit31
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit0
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit1
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit2
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit3
timestamp 1688980957
transform 1 0 18216 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit4
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit5
timestamp 1688980957
transform 1 0 22356 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit6
timestamp 1688980957
transform 1 0 21252 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit7
timestamp 1688980957
transform 1 0 22356 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit8
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit9
timestamp 1688980957
transform 1 0 19964 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit10
timestamp 1688980957
transform 1 0 17572 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit11
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit12
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit13
timestamp 1688980957
transform 1 0 22448 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit14
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit15
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit16
timestamp 1688980957
transform 1 0 19872 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit17
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit18
timestamp 1688980957
transform 1 0 19596 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit19
timestamp 1688980957
transform 1 0 17940 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit20
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit21
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit22
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit23
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit24
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit25
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit26
timestamp 1688980957
transform 1 0 22724 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit27
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit28
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit29
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit30
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit31
timestamp 1688980957
transform 1 0 19136 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit24
timestamp 1688980957
transform 1 0 19320 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit25
timestamp 1688980957
transform 1 0 19228 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit26
timestamp 1688980957
transform 1 0 22264 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit27
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit28
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit29
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit30
timestamp 1688980957
transform 1 0 22448 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit31
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 3680 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 3864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._36_
timestamp 1688980957
transform 1 0 4324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._37_
timestamp 1688980957
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._38_
timestamp 1688980957
transform 1 0 4692 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._39_
timestamp 1688980957
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._40_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._41_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._42_
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._43_
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._44_
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._45_
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._46_
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._47_
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 8004 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2
timestamp 1688980957
transform 1 0 4968 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 14720 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 14996 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 16008 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 6348 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 6900 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 2852 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 13156 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 11776 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 17112 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 11224 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 2576 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 12788 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 2668 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 9936 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 11316 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 4324 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 9844 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 15732 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 11776 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 16652 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 3864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 1748 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 9844 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 10856 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 14260 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 4784 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 10396 0 1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 8464 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 11316 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 8740 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 3220 0 -1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 8004 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 7268 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 3312 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 8924 0 -1 40256
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 13064 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1472 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 11408 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 8648 0 -1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1472 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 6900 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 1564 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1840 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 4784 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 13892 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 11408 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 6164 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 14076 0 -1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 1748 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 2392 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 6256 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 14628 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 1748 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 1748 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 8096 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 14260 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 5428 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 5336 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 3496 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 2852 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 3680 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 5704 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 2392 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 11040 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 11316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 10580 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10488 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9016 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9200 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8280 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7912 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6992 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5060 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 9292 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 9108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 8832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6808 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 17020 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 17296 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 15548 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 15548 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 15824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14996 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 12788 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 13064 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 7452 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7636 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 13892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12512 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12788 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 10488 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 10488 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 4508 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 5704 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 6900 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 7176 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 7728 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 8004 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 9200 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 7084 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 7636 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 8188 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 8464 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 23552 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1688980957
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 23736 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 23368 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 23368 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1688980957
transform 1 0 23644 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 23552 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output206
timestamp 1688980957
transform 1 0 23736 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output209
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output213
timestamp 1688980957
transform 1 0 23552 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output216
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output217
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1688980957
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 23460 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output220
timestamp 1688980957
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1688980957
transform 1 0 24196 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1688980957
transform 1 0 24196 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1688980957
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output224
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1688980957
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output228
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1688980957
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output231
timestamp 1688980957
transform 1 0 23736 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1688980957
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1688980957
transform 1 0 24196 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1688980957
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output235
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1688980957
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output238
timestamp 1688980957
transform 1 0 23736 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output239
timestamp 1688980957
transform 1 0 23276 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 23920 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1688980957
transform 1 0 23920 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output242
timestamp 1688980957
transform 1 0 23092 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output243
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output244
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 22724 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1688980957
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1688980957
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1688980957
transform 1 0 24196 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1688980957
transform 1 0 19872 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 23276 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 22724 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 22080 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 22632 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 23276 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 21988 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 23828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 23184 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 22172 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output264
timestamp 1688980957
transform 1 0 20792 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1688980957
transform 1 0 21344 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output267
timestamp 1688980957
transform 1 0 22172 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 22724 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output269
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 20240 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 21160 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output273
timestamp 1688980957
transform 1 0 2944 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output278
timestamp 1688980957
transform 1 0 1932 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output279
timestamp 1688980957
transform 1 0 1656 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output282
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output283
timestamp 1688980957
transform 1 0 2392 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1688980957
transform 1 0 2760 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1688980957
transform 1 0 3956 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 3956 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output288
timestamp 1688980957
transform 1 0 4416 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output289
timestamp 1688980957
transform 1 0 4508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 4968 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1688980957
transform 1 0 4784 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output292
timestamp 1688980957
transform 1 0 5152 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output293
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output295
timestamp 1688980957
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1688980957
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output297
timestamp 1688980957
transform 1 0 9384 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output298
timestamp 1688980957
transform 1 0 9016 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output299
timestamp 1688980957
transform 1 0 9384 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output300
timestamp 1688980957
transform 1 0 5888 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1688980957
transform 1 0 5888 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output302
timestamp 1688980957
transform 1 0 6624 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 6624 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 7176 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1688980957
transform 1 0 7176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1688980957
transform 1 0 7544 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output308
timestamp 1688980957
transform 1 0 8280 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output309
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output310
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output311
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output314
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output318
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output319
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output320
timestamp 1688980957
transform 1 0 16100 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output321
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output322
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output323
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output325
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output326
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output328
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output329
timestamp 1688980957
transform 1 0 15548 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 19136 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output339
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output342
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 20516 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 2116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 2116 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 1564 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 1564 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 2852 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 1564 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 2116 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 3772 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 3220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 2300 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 2668 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 2668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 2116 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 24840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 24840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 24840 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 24840 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 24840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 24840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 24840 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 24840 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 24840 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 24840 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 24840 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 24840 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 24840 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 24840 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 24840 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 24840 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 24840 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 24840 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 24840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 24840 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 24840 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 24840 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 24840 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 24840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 24840 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 24840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 24840 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 24840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 24840 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 24840 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 24840 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 24840 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 24840 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 24840 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 24840 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 24840 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 24840 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 24840 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 24840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 24840 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 24840 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 24840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 24840 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 24840 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 17020 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 17388 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 18124 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 18492 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 18216 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 19136 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 16928 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 17204 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 17480 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 17756 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 18032 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 18308 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 18584 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 18676 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 19504 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 19044 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 19596 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 20056 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 20700 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 20884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 21436 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 22356 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 19780 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 23460 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 22356 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 23920 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 20240 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 20700 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 21712 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 21528 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 22172 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 22724 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 22632 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 21896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 23368 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 23736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 23368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 22448 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 23184 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23828 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 23920 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 24288 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 25840 9256 26000 9376 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 25840 9800 26000 9920 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 25840 10344 26000 10464 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 25840 10888 26000 11008 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s 0 17960 160 18080 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s 0 18232 160 18352 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s 0 18504 160 18624 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s 0 18776 160 18896 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s 0 21224 160 21344 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s 0 21496 160 21616 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s 0 21768 160 21888 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s 0 22040 160 22160 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s 0 22312 160 22432 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s 0 22584 160 22704 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s 0 22856 160 22976 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s 0 23128 160 23248 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s 0 19048 160 19168 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s 0 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s 0 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s 0 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s 0 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s 0 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s 0 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s 0 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s 0 27752 160 27872 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s 0 30472 160 30592 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s 0 30744 160 30864 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s 0 28024 160 28144 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s 0 28296 160 28416 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s 0 28568 160 28688 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s 0 28840 160 28960 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s 0 29112 160 29232 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s 0 29384 160 29504 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s 0 29656 160 29776 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s 0 29928 160 30048 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s 0 30200 160 30320 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s 0 23400 160 23520 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s 0 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s 0 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s 0 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s 0 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s 0 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s 0 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s 0 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s 0 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s 0 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s 0 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s 0 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s 0 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s 0 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s 0 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s 0 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 25840 15784 26000 15904 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 25840 16328 26000 16448 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 25840 16872 26000 16992 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 25840 17416 26000 17536 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 25840 13608 26000 13728 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 25840 14152 26000 14272 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 25840 14696 26000 14816 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 25840 15240 26000 15360 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 25840 11432 26000 11552 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 25840 11976 26000 12096 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 25840 12520 26000 12640 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 25840 13064 26000 13184 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 25840 24488 26000 24608 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 25840 25032 26000 25152 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 25840 25576 26000 25696 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 25840 26120 26000 26240 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 25840 22312 26000 22432 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 25840 22856 26000 22976 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 25840 23400 26000 23520 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 25840 23944 26000 24064 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 25840 20136 26000 20256 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 25840 20680 26000 20800 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 25840 21224 26000 21344 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 25840 21768 26000 21888 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 25840 17960 26000 18080 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 25840 18504 26000 18624 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 25840 19048 26000 19168 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 25840 19592 26000 19712 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s 0 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s 0 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s 0 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s 0 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s 0 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s 0 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s 0 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s 0 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s 0 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s 0 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s 0 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s 0 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s 0 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s 0 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s 0 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s 0 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s 0 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s 0 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s 0 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s 0 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s 0 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s 0 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s 0 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s 0 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s 0 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s 0 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s 0 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s 0 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s 0 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s 0 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s 0 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 25840 26664 26000 26784 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 25840 32104 26000 32224 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 25840 32648 26000 32768 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 25840 33192 26000 33312 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 25840 33736 26000 33856 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 25840 34280 26000 34400 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 25840 34824 26000 34944 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 25840 35368 26000 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 25840 35912 26000 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 25840 36456 26000 36576 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 25840 37000 26000 37120 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 25840 27208 26000 27328 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 25840 37544 26000 37664 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 25840 38088 26000 38208 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 25840 38632 26000 38752 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 25840 39176 26000 39296 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 25840 39720 26000 39840 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 25840 40264 26000 40384 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 25840 40808 26000 40928 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 25840 41352 26000 41472 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 25840 41896 26000 42016 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 25840 42440 26000 42560 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 25840 27752 26000 27872 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 25840 42984 26000 43104 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 25840 43528 26000 43648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 25840 28296 26000 28416 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 25840 28840 26000 28960 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 25840 29384 26000 29504 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 25840 29928 26000 30048 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 25840 30472 26000 30592 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 25840 31016 26000 31136 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 25840 31560 26000 31680 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 20350 44463 20406 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 23110 44463 23166 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 23386 44463 23442 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 23662 44463 23718 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 23938 44463 23994 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 24214 44463 24270 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 24490 44463 24546 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 24766 44463 24822 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 25042 44463 25098 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 25318 44463 25374 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 25594 44463 25650 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 20626 44463 20682 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 20902 44463 20958 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 21178 44463 21234 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 21454 44463 21510 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 21730 44463 21786 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 22006 44463 22062 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 22282 44463 22338 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 22558 44463 22614 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 22834 44463 22890 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 202 44463 258 44623 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 478 44463 534 44623 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 754 44463 810 44623 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 1030 44463 1086 44623 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 1306 44463 1362 44623 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 1582 44463 1638 44623 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 1858 44463 1914 44623 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 2134 44463 2190 44623 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 2410 44463 2466 44623 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 2686 44463 2742 44623 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 2962 44463 3018 44623 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 3238 44463 3294 44623 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 3514 44463 3570 44623 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 3790 44463 3846 44623 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 4066 44463 4122 44623 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 4342 44463 4398 44623 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 4618 44463 4674 44623 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 4894 44463 4950 44623 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 5170 44463 5226 44623 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 5446 44463 5502 44623 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 5722 44463 5778 44623 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 8482 44463 8538 44623 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8758 44463 8814 44623 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 9034 44463 9090 44623 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 9310 44463 9366 44623 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 9586 44463 9642 44623 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 9862 44463 9918 44623 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 5998 44463 6054 44623 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 6274 44463 6330 44623 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 6550 44463 6606 44623 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 6826 44463 6882 44623 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7102 44463 7158 44623 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7378 44463 7434 44623 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7654 44463 7710 44623 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 7930 44463 7986 44623 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 8206 44463 8262 44623 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 25840 7080 26000 7200 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 25840 7624 26000 7744 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 25840 8168 26000 8288 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 25840 8712 26000 8832 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 25840 4904 26000 5024 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 25840 5448 26000 5568 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 25840 5992 26000 6112 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 25840 6536 26000 6656 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 25840 2728 26000 2848 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 25840 3272 26000 3392 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 25840 3816 26000 3936 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 25840 4360 26000 4480 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 25840 552 26000 672 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 25840 1096 26000 1216 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 25840 1640 26000 1760 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 25840 2184 26000 2304 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 10138 44463 10194 44623 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 10414 44463 10470 44623 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 10690 44463 10746 44623 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 10966 44463 11022 44623 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 11242 44463 11298 44623 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 11518 44463 11574 44623 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 11794 44463 11850 44623 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 12070 44463 12126 44623 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 12346 44463 12402 44623 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 12622 44463 12678 44623 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 12898 44463 12954 44623 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 13174 44463 13230 44623 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 13450 44463 13506 44623 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 13726 44463 13782 44623 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 14002 44463 14058 44623 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 14278 44463 14334 44623 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 14554 44463 14610 44623 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 14830 44463 14886 44623 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 15106 44463 15162 44623 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 15382 44463 15438 44623 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 15658 44463 15714 44623 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 18418 44463 18474 44623 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 18694 44463 18750 44623 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 18970 44463 19026 44623 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 19246 44463 19302 44623 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 19522 44463 19578 44623 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 19798 44463 19854 44623 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 15934 44463 15990 44623 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 16210 44463 16266 44623 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 16486 44463 16542 44623 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 16762 44463 16818 44623 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 17038 44463 17094 44623 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 17314 44463 17370 44623 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 17590 44463 17646 44623 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 17866 44463 17922 44623 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 18142 44463 18198 44623 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 20074 44463 20130 44623 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 6878 1040 7198 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 9845 1040 10165 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 15779 1040 16099 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 21713 1040 22033 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s 0 4904 160 5024 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s 0 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s 0 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s 0 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s 0 5992 160 6112 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s 0 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s 0 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s 0 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s 0 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s 0 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s 0 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s 0 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s 0 8168 160 8288 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s 0 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s 0 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s 0 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s 0 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s 0 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s 0 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s 0 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s 0 14696 160 14816 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s 0 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s 0 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s 0 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s 0 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s 0 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s 0 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s 0 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s 0 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s 0 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s 0 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s 0 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s 0 10344 160 10464 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s 0 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s 0 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s 0 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s 0 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s 0 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s 0 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s 0 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s 0 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s 0 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s 0 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s 0 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s 0 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s 0 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s 0 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s 0 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 13052 43520 13052 43520 0 VGND
rlabel metal1 12972 42976 12972 42976 0 VPWR
rlabel metal1 24012 9146 24012 9146 0 Config_accessC_bit0
rlabel metal1 24748 7310 24748 7310 0 Config_accessC_bit1
rlabel metal2 23414 9775 23414 9775 0 Config_accessC_bit2
rlabel metal3 25572 10948 25572 10948 0 Config_accessC_bit3
rlabel metal3 682 18020 682 18020 0 E1END[0]
rlabel metal3 728 18292 728 18292 0 E1END[1]
rlabel metal3 820 18564 820 18564 0 E1END[2]
rlabel metal3 774 18836 774 18836 0 E1END[3]
rlabel metal3 682 21284 682 21284 0 E2END[0]
rlabel metal3 682 21556 682 21556 0 E2END[1]
rlabel metal3 728 21828 728 21828 0 E2END[2]
rlabel metal2 3588 21998 3588 21998 0 E2END[3]
rlabel metal3 820 22372 820 22372 0 E2END[4]
rlabel metal3 843 22644 843 22644 0 E2END[5]
rlabel metal3 728 22916 728 22916 0 E2END[6]
rlabel metal3 866 23188 866 23188 0 E2END[7]
rlabel metal2 3358 19227 3358 19227 0 E2MID[0]
rlabel metal3 958 19380 958 19380 0 E2MID[1]
rlabel metal3 728 19652 728 19652 0 E2MID[2]
rlabel metal3 498 19924 498 19924 0 E2MID[3]
rlabel metal3 452 20196 452 20196 0 E2MID[4]
rlabel metal3 774 20468 774 20468 0 E2MID[5]
rlabel metal3 728 20740 728 20740 0 E2MID[6]
rlabel metal3 728 21012 728 21012 0 E2MID[7]
rlabel metal3 452 27812 452 27812 0 E6END[0]
rlabel metal2 3726 30379 3726 30379 0 E6END[10]
rlabel metal3 728 30804 728 30804 0 E6END[11]
rlabel metal2 3174 28815 3174 28815 0 E6END[1]
rlabel metal3 452 28356 452 28356 0 E6END[2]
rlabel metal3 475 28628 475 28628 0 E6END[3]
rlabel metal2 3634 29019 3634 29019 0 E6END[4]
rlabel metal3 1740 29172 1740 29172 0 E6END[5]
rlabel metal3 728 29444 728 29444 0 E6END[6]
rlabel metal3 544 29716 544 29716 0 E6END[7]
rlabel metal3 475 29988 475 29988 0 E6END[8]
rlabel metal2 3818 30481 3818 30481 0 E6END[9]
rlabel metal3 452 23460 452 23460 0 EE4END[0]
rlabel metal2 3818 26265 3818 26265 0 EE4END[10]
rlabel metal3 682 26452 682 26452 0 EE4END[11]
rlabel metal3 774 26724 774 26724 0 EE4END[12]
rlabel metal3 958 26996 958 26996 0 EE4END[13]
rlabel metal3 659 27268 659 27268 0 EE4END[14]
rlabel metal3 567 27540 567 27540 0 EE4END[15]
rlabel metal3 590 23732 590 23732 0 EE4END[1]
rlabel metal3 774 24004 774 24004 0 EE4END[2]
rlabel metal3 912 24276 912 24276 0 EE4END[3]
rlabel metal3 636 24548 636 24548 0 EE4END[4]
rlabel metal3 1142 24820 1142 24820 0 EE4END[5]
rlabel metal3 682 25092 682 25092 0 EE4END[6]
rlabel metal3 728 25364 728 25364 0 EE4END[7]
rlabel metal2 2898 25993 2898 25993 0 EE4END[8]
rlabel metal2 3450 26129 3450 26129 0 EE4END[9]
rlabel metal2 24150 15759 24150 15759 0 FAB2RAM_A0_O0
rlabel metal3 25503 16388 25503 16388 0 FAB2RAM_A0_O1
rlabel metal3 25020 16932 25020 16932 0 FAB2RAM_A0_O2
rlabel metal1 24380 17306 24380 17306 0 FAB2RAM_A0_O3
rlabel metal3 25158 13668 25158 13668 0 FAB2RAM_A1_O0
rlabel metal3 25526 14212 25526 14212 0 FAB2RAM_A1_O1
rlabel metal3 24974 14756 24974 14756 0 FAB2RAM_A1_O2
rlabel metal1 24840 14450 24840 14450 0 FAB2RAM_A1_O3
rlabel metal3 24882 11492 24882 11492 0 FAB2RAM_C_O0
rlabel metal3 25572 12036 25572 12036 0 FAB2RAM_C_O1
rlabel metal3 25066 12580 25066 12580 0 FAB2RAM_C_O2
rlabel metal3 25687 13124 25687 13124 0 FAB2RAM_C_O3
rlabel metal3 25158 24548 25158 24548 0 FAB2RAM_D0_O0
rlabel metal3 25526 25092 25526 25092 0 FAB2RAM_D0_O1
rlabel metal3 25158 25636 25158 25636 0 FAB2RAM_D0_O2
rlabel metal3 25526 26180 25526 26180 0 FAB2RAM_D0_O3
rlabel metal1 24472 21658 24472 21658 0 FAB2RAM_D1_O0
rlabel metal3 25526 22916 25526 22916 0 FAB2RAM_D1_O1
rlabel metal3 25158 23460 25158 23460 0 FAB2RAM_D1_O2
rlabel metal3 25526 24004 25526 24004 0 FAB2RAM_D1_O3
rlabel metal1 24012 20026 24012 20026 0 FAB2RAM_D2_O0
rlabel metal1 24794 19278 24794 19278 0 FAB2RAM_D2_O1
rlabel metal3 24882 21284 24882 21284 0 FAB2RAM_D2_O2
rlabel metal3 25526 21828 25526 21828 0 FAB2RAM_D2_O3
rlabel metal3 25158 18020 25158 18020 0 FAB2RAM_D3_O0
rlabel metal3 25526 18564 25526 18564 0 FAB2RAM_D3_O1
rlabel metal3 24882 19108 24882 19108 0 FAB2RAM_D3_O2
rlabel metal1 24886 18734 24886 18734 0 FAB2RAM_D3_O3
rlabel metal3 1464 31076 1464 31076 0 FrameData[0]
rlabel metal3 774 33796 774 33796 0 FrameData[10]
rlabel metal2 3450 34867 3450 34867 0 FrameData[11]
rlabel metal3 1441 34340 1441 34340 0 FrameData[12]
rlabel metal3 452 34612 452 34612 0 FrameData[13]
rlabel metal3 774 34884 774 34884 0 FrameData[14]
rlabel metal2 3818 35649 3818 35649 0 FrameData[15]
rlabel metal3 866 35428 866 35428 0 FrameData[16]
rlabel metal2 2806 35972 2806 35972 0 FrameData[17]
rlabel via2 3634 35989 3634 35989 0 FrameData[18]
rlabel metal3 912 36244 912 36244 0 FrameData[19]
rlabel metal3 774 31348 774 31348 0 FrameData[1]
rlabel metal3 1050 36516 1050 36516 0 FrameData[20]
rlabel metal2 3174 38403 3174 38403 0 FrameData[21]
rlabel metal2 3910 37247 3910 37247 0 FrameData[22]
rlabel metal2 4922 37553 4922 37553 0 FrameData[23]
rlabel metal3 774 37604 774 37604 0 FrameData[24]
rlabel metal3 452 37876 452 37876 0 FrameData[25]
rlabel metal3 682 38148 682 38148 0 FrameData[26]
rlabel metal2 3082 38675 3082 38675 0 FrameData[27]
rlabel metal3 1441 38692 1441 38692 0 FrameData[28]
rlabel metal2 2806 39695 2806 39695 0 FrameData[29]
rlabel metal3 1970 31620 1970 31620 0 FrameData[2]
rlabel metal3 774 39236 774 39236 0 FrameData[30]
rlabel metal3 820 39508 820 39508 0 FrameData[31]
rlabel metal3 682 31892 682 31892 0 FrameData[3]
rlabel metal3 636 32164 636 32164 0 FrameData[4]
rlabel metal3 682 32436 682 32436 0 FrameData[5]
rlabel metal2 2806 33337 2806 33337 0 FrameData[6]
rlabel metal3 820 32980 820 32980 0 FrameData[7]
rlabel metal2 2898 33660 2898 33660 0 FrameData[8]
rlabel metal3 682 33524 682 33524 0 FrameData[9]
rlabel metal3 25158 26724 25158 26724 0 FrameData_O[0]
rlabel metal3 25158 32164 25158 32164 0 FrameData_O[10]
rlabel metal3 25572 32708 25572 32708 0 FrameData_O[11]
rlabel metal3 25158 33252 25158 33252 0 FrameData_O[12]
rlabel metal3 25572 33796 25572 33796 0 FrameData_O[13]
rlabel metal3 25503 34340 25503 34340 0 FrameData_O[14]
rlabel metal3 25572 34884 25572 34884 0 FrameData_O[15]
rlabel metal3 25158 35428 25158 35428 0 FrameData_O[16]
rlabel metal3 25526 35972 25526 35972 0 FrameData_O[17]
rlabel metal3 25158 36516 25158 36516 0 FrameData_O[18]
rlabel metal3 25503 37060 25503 37060 0 FrameData_O[19]
rlabel metal3 25526 27268 25526 27268 0 FrameData_O[1]
rlabel metal3 25158 37604 25158 37604 0 FrameData_O[20]
rlabel metal3 25572 38148 25572 38148 0 FrameData_O[21]
rlabel metal3 25158 38692 25158 38692 0 FrameData_O[22]
rlabel metal3 25572 39236 25572 39236 0 FrameData_O[23]
rlabel metal3 25158 39780 25158 39780 0 FrameData_O[24]
rlabel metal3 25526 40324 25526 40324 0 FrameData_O[25]
rlabel metal3 24790 40868 24790 40868 0 FrameData_O[26]
rlabel metal3 25572 41412 25572 41412 0 FrameData_O[27]
rlabel metal3 25020 41956 25020 41956 0 FrameData_O[28]
rlabel metal3 25526 42500 25526 42500 0 FrameData_O[29]
rlabel metal3 25158 27812 25158 27812 0 FrameData_O[2]
rlabel metal1 24748 41786 24748 41786 0 FrameData_O[30]
rlabel metal1 23184 42330 23184 42330 0 FrameData_O[31]
rlabel metal3 25526 28356 25526 28356 0 FrameData_O[3]
rlabel metal3 25158 28900 25158 28900 0 FrameData_O[4]
rlabel metal3 25526 29444 25526 29444 0 FrameData_O[5]
rlabel metal3 25158 29988 25158 29988 0 FrameData_O[6]
rlabel metal3 25526 30532 25526 30532 0 FrameData_O[7]
rlabel metal3 25158 31076 25158 31076 0 FrameData_O[8]
rlabel metal1 24702 31790 24702 31790 0 FrameData_O[9]
rlabel metal1 19734 1836 19734 1836 0 FrameStrobe[0]
rlabel metal1 23460 3502 23460 3502 0 FrameStrobe[10]
rlabel metal2 20562 1020 20562 1020 0 FrameStrobe[11]
rlabel metal2 23743 68 23743 68 0 FrameStrobe[12]
rlabel metal1 21758 5576 21758 5576 0 FrameStrobe[13]
rlabel metal2 24242 296 24242 296 0 FrameStrobe[14]
rlabel metal1 19734 3060 19734 3060 0 FrameStrobe[15]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[16]
rlabel metal2 19550 2244 19550 2244 0 FrameStrobe[17]
rlabel metal1 21298 1972 21298 1972 0 FrameStrobe[18]
rlabel metal2 21206 1122 21206 1122 0 FrameStrobe[19]
rlabel metal2 20654 908 20654 908 0 FrameStrobe[1]
rlabel metal1 20884 1938 20884 1938 0 FrameStrobe[2]
rlabel metal2 21206 262 21206 262 0 FrameStrobe[3]
rlabel metal2 21482 1248 21482 1248 0 FrameStrobe[4]
rlabel metal1 21436 1870 21436 1870 0 FrameStrobe[5]
rlabel metal2 22034 364 22034 364 0 FrameStrobe[6]
rlabel metal1 22494 3502 22494 3502 0 FrameStrobe[7]
rlabel metal2 22685 68 22685 68 0 FrameStrobe[8]
rlabel metal1 20654 2448 20654 2448 0 FrameStrobe[9]
rlabel metal1 20240 43418 20240 43418 0 FrameStrobe_O[0]
rlabel metal2 23138 43972 23138 43972 0 FrameStrobe_O[10]
rlabel metal1 23276 41242 23276 41242 0 FrameStrobe_O[11]
rlabel metal1 23092 41446 23092 41446 0 FrameStrobe_O[12]
rlabel metal1 23506 41786 23506 41786 0 FrameStrobe_O[13]
rlabel metal1 24196 42670 24196 42670 0 FrameStrobe_O[14]
rlabel metal1 24104 42330 24104 42330 0 FrameStrobe_O[15]
rlabel metal1 23184 42670 23184 42670 0 FrameStrobe_O[16]
rlabel metal1 24656 41242 24656 41242 0 FrameStrobe_O[17]
rlabel metal1 24518 41718 24518 41718 0 FrameStrobe_O[18]
rlabel metal1 24104 42126 24104 42126 0 FrameStrobe_O[19]
rlabel metal2 20654 43972 20654 43972 0 FrameStrobe_O[1]
rlabel metal1 21252 43146 21252 43146 0 FrameStrobe_O[2]
rlabel metal1 21620 43418 21620 43418 0 FrameStrobe_O[3]
rlabel metal1 22402 43384 22402 43384 0 FrameStrobe_O[4]
rlabel metal2 21758 43802 21758 43802 0 FrameStrobe_O[5]
rlabel metal2 22126 42959 22126 42959 0 FrameStrobe_O[6]
rlabel metal2 22310 43632 22310 43632 0 FrameStrobe_O[7]
rlabel metal2 22586 43870 22586 43870 0 FrameStrobe_O[8]
rlabel metal1 22862 42296 22862 42296 0 FrameStrobe_O[9]
rlabel metal1 24058 9554 24058 9554 0 Inst_Config_accessConfig_access.ConfigBits\[0\]
rlabel metal1 24518 8500 24518 8500 0 Inst_Config_accessConfig_access.ConfigBits\[1\]
rlabel metal1 22678 10540 22678 10540 0 Inst_Config_accessConfig_access.ConfigBits\[2\]
rlabel metal1 23644 11322 23644 11322 0 Inst_Config_accessConfig_access.ConfigBits\[3\]
rlabel metal2 19826 15164 19826 15164 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21942 17000 21942 17000 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23644 17850 23644 17850 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 22494 19380 22494 19380 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18062 16150 18062 16150 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 20966 17578 20966 17578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 15134 18360 15134 18360 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 20920 19822 20920 19822 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19826 16116 19826 16116 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22678 17714 22678 17714 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23552 16558 23552 16558 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal2 22126 20230 22126 20230 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18630 15674 18630 15674 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 20010 15436 20010 15436 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 19550 15436 19550 15436 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19826 14926 19826 14926 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 22218 17476 22218 17476 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21666 17204 21666 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21850 16694 21850 16694 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22172 16626 22172 16626 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 24334 17204 24334 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23138 16422 23138 16422 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 24288 16082 24288 16082 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 24012 16014 24012 16014 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21850 19380 21850 19380 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal2 22678 19822 22678 19822 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 22034 19312 22034 19312 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 22494 19278 22494 19278 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19182 13906 19182 13906 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 24242 14620 24242 14620 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23690 20570 23690 20570 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20378 19346 20378 19346 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18354 14314 18354 14314 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
rlabel via2 7866 21403 7866 21403 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
rlabel metal2 17158 25398 17158 25398 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18446 19822 18446 19822 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18722 14382 18722 14382 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23322 14348 23322 14348 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23368 19346 23368 19346 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20424 18734 20424 18734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18446 14416 18446 14416 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19642 13940 19642 13940 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18584 13498 18584 13498 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18906 13362 18906 13362 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23092 14994 23092 14994 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 22954 13940 22954 13940 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23920 14858 23920 14858 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 22862 14450 22862 14450 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 22954 20230 22954 20230 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23230 19278 23230 19278 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 24242 20604 24242 20604 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23966 20366 23966 20366 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 19642 18802 19642 18802 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20562 18870 20562 18870 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 20010 18938 20010 18938 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20930 19278 20930 19278 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 21850 14450 21850 14450 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20746 31178 20746 31178 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23046 37706 23046 37706 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel via1 21022 16422 21022 16422 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 20460 14994 20460 14994 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 8234 33031 8234 33031 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 21436 38930 21436 38930 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 19596 17170 19596 17170 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 22218 14586 22218 14586 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20700 31790 20700 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\]
rlabel metal2 23506 38556 23506 38556 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20700 17170 20700 17170 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21482 14348 21482 14348 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 22678 14348 22678 14348 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21758 14586 21758 14586 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22356 14450 22356 14450 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20102 31824 20102 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20700 31926 20700 31926 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20332 31790 20332 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21114 30906 21114 30906 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 22126 38522 22126 38522 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 22954 38420 22954 38420 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23046 37842 23046 37842 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23782 37944 23782 37944 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20102 17204 20102 17204 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20792 16082 20792 16082 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 20746 16762 20746 16762 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21160 16218 21160 16218 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 22218 29716 22218 29716 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20976 28050 20976 28050 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18814 35666 18814 35666 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19780 28934 19780 28934 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 21068 29614 21068 29614 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 5750 28152 5750 28152 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 14796 36074 14796 36074 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18262 28526 18262 28526 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 22310 30362 22310 30362 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20976 27438 20976 27438 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 18814 36108 18814 36108 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19274 27982 19274 27982 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21666 29580 21666 29580 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 22586 30090 22586 30090 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21942 29682 21942 29682 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 22402 29682 22402 29682 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20378 27574 20378 27574 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21022 27574 21022 27574 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21206 27914 21206 27914 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21574 27982 21574 27982 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18078 35054 18078 35054 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19550 35700 19550 35700 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18676 35258 18676 35258 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19366 35598 19366 35598 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 19274 28560 19274 28560 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19228 28730 19228 28730 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19550 28594 19550 28594 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19964 28594 19964 28594 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 21482 22372 21482 22372 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 23460 25262 23460 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18676 33490 18676 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19826 25874 19826 25874 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 20132 23018 20132 23018 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
rlabel metal2 4922 24208 4922 24208 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 17424 33490 17424 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 18998 26758 18998 26758 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 22356 21998 22356 21998 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23414 25398 23414 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19550 33388 19550 33388 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 19688 25262 19688 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 21436 22746 21436 22746 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 22448 22134 22448 22134 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 22172 22202 22172 22202 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21942 22406 21942 22406 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23046 25908 23046 25908 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23552 26010 23552 26010 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23322 25466 23322 25466 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23690 25398 23690 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18170 34000 18170 34000 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19320 33490 19320 33490 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18538 33422 18538 33422 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19090 33422 19090 33422 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 19274 25738 19274 25738 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20010 25398 20010 25398 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19734 25466 19734 25466 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20378 25806 20378 25806 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20884 21658 20884 21658 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 22678 27404 22678 27404 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20838 33966 20838 33966 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19274 30634 19274 30634 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17894 26316 17894 26316 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 21098 27370 21098 27370 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
rlabel via1 19361 34578 19361 34578 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 17802 30906 17802 30906 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20792 21862 20792 21862 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 22724 27642 22724 27642 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 21022 34612 21022 34612 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20102 30804 20102 30804 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 20010 20910 20010 20910 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 20746 21488 20746 21488 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20930 21114 20930 21114 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21482 21454 21482 21454 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 22908 27438 22908 27438 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23506 27506 23506 27506 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22954 27574 22954 27574 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23184 27506 23184 27506 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20056 34578 20056 34578 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 21574 34170 21574 34170 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 21114 34340 21114 34340 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21390 34034 21390 34034 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18538 31280 18538 31280 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19872 30702 19872 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18998 30906 18998 30906 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 19642 30770 19642 30770 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20010 23494 20010 23494 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 23138 22039 23138 22039 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23230 33490 23230 33490 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 21390 25670 21390 25670 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18068 23698 18068 23698 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 17250 24888 17250 24888 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 21344 33490 21344 33490 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 20138 24786 20138 24786 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 19274 24004 19274 24004 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 23874 23290 23874 23290 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 23046 33626 23046 33626 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 21758 24786 21758 24786 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19274 23120 19274 23120 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20010 24276 20010 24276 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19550 23154 19550 23154 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19918 23222 19918 23222 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23506 23732 23506 23732 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23414 23664 23414 23664 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 23414 22202 23414 22202 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel via1 23414 22073 23414 22073 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel via1 22218 32879 22218 32879 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 23874 33422 23874 33422 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 22862 33082 22862 33082 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23690 33422 23690 33422 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20930 24140 20930 24140 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21712 24922 21712 24922 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21252 24378 21252 24378 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 21620 24718 21620 24718 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 20378 7412 20378 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20194 10778 20194 10778 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23460 7514 23460 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 21850 9792 21850 9792 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18315 8466 18315 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
rlabel metal1 13754 11050 13754 11050 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
rlabel metal2 1886 16949 1886 16949 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
rlabel metal1 9384 9622 9384 9622 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
rlabel metal1 21804 7378 21804 7378 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
rlabel metal2 21114 10166 21114 10166 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 22494 7820 22494 7820 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 22586 9146 22586 9146 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 20792 6970 20792 6970 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21298 6766 21298 6766 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20332 7514 20332 7514 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 21114 7412 21114 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20240 10030 20240 10030 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20884 10642 20884 10642 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20240 10234 20240 10234 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 20746 10948 20746 10948 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 24012 7242 24012 7242 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 24150 6868 24150 6868 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 22862 8058 22862 8058 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 24058 7650 24058 7650 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21850 9520 21850 9520 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 22310 9622 22310 9622 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 22126 8908 22126 8908 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 22494 8466 22494 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19596 7854 19596 7854 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 21896 11662 21896 11662 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 23230 4454 23230 4454 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 22862 6222 22862 6222 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 16836 8058 16836 8058 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
rlabel metal1 2070 12274 2070 12274 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
rlabel metal1 3634 12750 3634 12750 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
rlabel metal1 20654 6324 20654 6324 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
rlabel metal1 19734 7514 19734 7514 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 23460 12206 23460 12206 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 22586 5236 22586 5236 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 21574 5848 21574 5848 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
rlabel metal2 18630 7412 18630 7412 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 20056 8058 20056 8058 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19458 7888 19458 7888 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19918 7786 19918 7786 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 22770 12036 22770 12036 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 23276 12206 23276 12206 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22402 11764 22402 11764 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 22954 11730 22954 11730 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 23506 6324 23506 6324 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 22351 1326 22351 1326 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 23598 5780 23598 5780 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 23092 1190 23092 1190 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 21252 6290 21252 6290 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 23414 6256 23414 6256 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 21528 6358 21528 6358 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 23046 6426 23046 6426 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 19366 5372 19366 5372 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20838 5134 20838 5134 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18998 11186 18998 11186 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19504 13294 19504 13294 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 8878 6188 8878 6188 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\]
rlabel metal2 20746 5151 20746 5151 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\]
rlabel metal1 18722 11288 18722 11288 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\]
rlabel metal2 20194 13090 20194 13090 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\]
rlabel metal2 20654 4148 20654 4148 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 21574 4250 21574 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 19136 10030 19136 10030 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 21574 12784 21574 12784 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 19228 4250 19228 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19734 4556 19734 4556 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19274 4794 19274 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19495 5202 19495 5202 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 20930 5066 20930 5066 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21436 4590 21436 4590 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 21114 4794 21114 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21436 4794 21436 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17940 10030 17940 10030 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 19918 10506 19918 10506 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18538 10234 18538 10234 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19228 11050 19228 11050 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20746 12614 20746 12614 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 21114 12954 21114 12954 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19918 13328 19918 13328 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20516 13226 20516 13226 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 18262 6086 18262 6086 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 23414 13396 23414 13396 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 21574 1394 21574 1394 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 21390 4080 21390 4080 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17940 6426 17940 6426 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\]
rlabel metal1 1564 14382 1564 14382 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\]
rlabel metal1 1104 10098 1104 10098 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\]
rlabel metal2 20838 3247 20838 3247 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\]
rlabel metal2 18814 4998 18814 4998 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 22494 13260 22494 13260 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 21942 4522 21942 4522 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 23920 2618 23920 2618 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
rlabel metal2 17710 4726 17710 4726 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18584 5202 18584 5202 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 18170 5746 18170 5746 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 18446 5780 18446 5780 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 23460 11866 23460 11866 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 22310 13736 22310 13736 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 22954 13498 22954 13498 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 23552 13974 23552 13974 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17434 3162 17434 3162 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 21712 3910 21712 3910 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 22448 4114 22448 4114 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21942 1190 21942 1190 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal4 22172 4964 22172 4964 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20286 4624 20286 4624 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 23920 3026 23920 3026 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20286 4216 20286 4216 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 12880 20366 12880 20366 0 Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
rlabel metal2 13570 20230 13570 20230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
rlabel metal2 5198 22236 5198 22236 0 Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 5428 21658 5428 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
rlabel metal1 9108 18394 9108 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
rlabel via1 9522 18683 9522 18683 0 Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
rlabel metal1 14628 18870 14628 18870 0 Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
rlabel metal1 15272 18394 15272 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 13478 27880 13478 27880 0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
rlabel metal2 14030 28220 14030 28220 0 Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
rlabel metal1 16146 26486 16146 26486 0 Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
rlabel metal2 5842 24990 5842 24990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
rlabel metal2 6394 24684 6394 24684 0 Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
rlabel metal2 7958 23324 7958 23324 0 Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 11086 30362 11086 30362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
rlabel via1 11914 30770 11914 30770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
rlabel metal1 13892 31314 13892 31314 0 Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
rlabel metal2 17296 21420 17296 21420 0 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
rlabel metal1 17940 21114 17940 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
rlabel metal1 18952 20978 18952 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
rlabel metal1 11546 5882 11546 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
rlabel metal2 12742 6086 12742 6086 0 Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
rlabel metal1 4462 17816 4462 17816 0 Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
rlabel metal2 5014 17850 5014 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
rlabel metal1 9656 11186 9656 11186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
rlabel metal1 10212 10778 10212 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
rlabel metal1 13524 4794 13524 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
rlabel metal1 14536 3706 14536 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
rlabel metal1 9338 6902 9338 6902 0 Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
rlabel metal1 10258 6834 10258 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
rlabel metal2 5014 5338 5014 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
rlabel metal2 5566 4998 5566 4998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
rlabel metal1 4508 9690 4508 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
rlabel metal2 5014 10268 5014 10268 0 Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
rlabel metal2 7406 5474 7406 5474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
rlabel metal1 7314 5882 7314 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
rlabel metal1 16008 5814 16008 5814 0 Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
rlabel metal1 17434 5338 17434 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
rlabel metal2 2438 12070 2438 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
rlabel metal1 3174 12274 3174 12274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
rlabel metal1 3082 3944 3082 3944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
rlabel metal2 3634 4556 3634 4556 0 Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
rlabel metal1 9568 3570 9568 3570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
rlabel metal1 10120 2074 10120 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
rlabel metal1 9016 5882 9016 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
rlabel metal2 10258 5780 10258 5780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
rlabel metal2 5014 6834 5014 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
rlabel metal2 5566 7140 5566 7140 0 Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
rlabel metal1 2392 17102 2392 17102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
rlabel metal2 2898 17884 2898 17884 0 Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
rlabel metal1 6440 7990 6440 7990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
rlabel metal2 7498 7684 7498 7684 0 Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
rlabel metal1 15456 4250 15456 4250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
rlabel metal2 16422 4964 16422 4964 0 Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
rlabel metal1 2438 14552 2438 14552 0 Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
rlabel metal1 3128 14042 3128 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
rlabel metal1 2576 2074 2576 2074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
rlabel metal1 3128 2618 3128 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
rlabel metal1 8280 3978 8280 3978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
rlabel metal1 9246 3162 9246 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
rlabel metal1 17986 7718 17986 7718 0 Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
rlabel metal1 17526 8568 17526 8568 0 Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
rlabel metal1 5474 14518 5474 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
rlabel metal1 6026 14042 6026 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
rlabel metal1 2576 9690 2576 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
rlabel metal1 3266 10098 3266 10098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
rlabel metal1 8280 8602 8280 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
rlabel metal1 8602 9146 8602 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
rlabel metal2 15870 10948 15870 10948 0 Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
rlabel metal1 16790 11186 16790 11186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
rlabel metal1 5980 11866 5980 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
rlabel metal1 6440 12274 6440 12274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
rlabel metal1 4416 12750 4416 12750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
rlabel metal1 4738 11866 4738 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
rlabel metal1 10442 13430 10442 13430 0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
rlabel metal1 11040 12954 11040 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
rlabel metal1 17563 11866 17563 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
rlabel metal1 17710 12274 17710 12274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
rlabel metal1 6164 9690 6164 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
rlabel metal1 7176 10098 7176 10098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
rlabel metal1 2438 17816 2438 17816 0 Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
rlabel metal2 2990 17850 2990 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
rlabel metal1 8280 12682 8280 12682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
rlabel metal2 9246 13260 9246 13260 0 Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
rlabel metal1 15962 8024 15962 8024 0 Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
rlabel metal1 16836 7922 16836 7922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
rlabel metal1 6992 14926 6992 14926 0 Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
rlabel metal1 7728 14586 7728 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
rlabel metal1 3036 7310 3036 7310 0 Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
rlabel metal1 3496 6970 3496 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
rlabel metal1 10258 8602 10258 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
rlabel metal1 10718 9146 10718 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
rlabel metal1 14950 14518 14950 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
rlabel metal1 15594 14042 15594 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
rlabel metal1 6118 39576 6118 39576 0 Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
rlabel metal2 6670 39916 6670 39916 0 Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
rlabel metal2 6026 39678 6026 39678 0 Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
rlabel metal1 6992 37978 6992 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
rlabel metal1 13156 13838 13156 13838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
rlabel metal2 13662 13668 13662 13668 0 Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
rlabel metal1 16698 13498 16698 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
rlabel metal1 17572 14042 17572 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
rlabel metal1 7590 11322 7590 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
rlabel metal1 8004 11866 8004 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
rlabel metal1 3680 15946 3680 15946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
rlabel metal1 4784 15674 4784 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
rlabel metal1 9660 15606 9660 15606 0 Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
rlabel metal1 10212 15130 10212 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
rlabel metal1 16422 16728 16422 16728 0 Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
rlabel metal1 17342 16626 17342 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
rlabel metal1 7728 15674 7728 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
rlabel metal2 8510 16422 8510 16422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
rlabel metal1 3450 20026 3450 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
rlabel metal2 4094 20604 4094 20604 0 Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
rlabel metal1 10488 17782 10488 17782 0 Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
rlabel metal1 11040 17306 11040 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
rlabel metal1 12519 25330 12519 25330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
rlabel metal2 12742 26282 12742 26282 0 Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
rlabel metal2 3266 28492 3266 28492 0 Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
rlabel metal1 3266 28118 3266 28118 0 Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
rlabel metal1 11040 36278 11040 36278 0 Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
rlabel metal2 12558 36414 12558 36414 0 Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
rlabel metal1 16468 28186 16468 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
rlabel via1 17249 28594 17249 28594 0 Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
rlabel metal2 13478 27982 13478 27982 0 Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
rlabel metal1 14260 26894 14260 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
rlabel metal2 3542 24276 3542 24276 0 Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
rlabel metal1 3542 22746 3542 22746 0 Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
rlabel metal1 10580 33014 10580 33014 0 Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
rlabel metal1 11132 32538 11132 32538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
rlabel metal1 17296 26894 17296 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
rlabel metal2 17894 27132 17894 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
rlabel metal2 11086 27132 11086 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
rlabel metal2 11914 27370 11914 27370 0 Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
rlabel metal1 4968 28390 4968 28390 0 Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
rlabel metal1 5520 27098 5520 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
rlabel metal1 10580 35190 10580 35190 0 Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
rlabel metal2 11086 34884 11086 34884 0 Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
rlabel metal1 16422 30872 16422 30872 0 Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
rlabel metal1 17204 30770 17204 30770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
rlabel metal1 13248 23630 13248 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
rlabel metal2 13846 23868 13846 23868 0 Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
rlabel metal1 3358 25364 3358 25364 0 Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
rlabel metal1 4416 25194 4416 25194 0 Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
rlabel metal2 12926 33184 12926 33184 0 Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
rlabel metal1 13340 33422 13340 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
rlabel metal1 17526 24922 17526 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
rlabel metal1 18492 24582 18492 24582 0 Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
rlabel metal1 16698 18938 16698 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
rlabel metal1 17296 19482 17296 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
rlabel metal1 7682 19958 7682 19958 0 Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
rlabel metal1 7820 18938 7820 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
rlabel metal2 5842 20060 5842 20060 0 Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
rlabel metal1 5750 19482 5750 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
rlabel metal2 15410 20774 15410 20774 0 Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
rlabel metal1 16054 20978 16054 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
rlabel metal2 15686 24038 15686 24038 0 Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
rlabel metal1 16468 24242 16468 24242 0 Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
rlabel metal1 7084 22406 7084 22406 0 Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
rlabel metal1 7544 21862 7544 21862 0 Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
rlabel metal1 7636 26214 7636 26214 0 Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
rlabel metal1 8050 25466 8050 25466 0 Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
rlabel metal1 14536 21658 14536 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
rlabel metal1 15226 22950 15226 22950 0 Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
rlabel metal1 12926 16218 12926 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
rlabel metal1 13478 17306 13478 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
rlabel metal1 2530 33388 2530 33388 0 Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
rlabel metal1 3404 33082 3404 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
rlabel metal1 12512 39882 12512 39882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
rlabel metal2 13386 39780 13386 39780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
rlabel metal1 18032 17850 18032 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
rlabel metal2 18354 18428 18354 18428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
rlabel metal1 10994 10132 10994 10132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
rlabel metal1 12742 9690 12742 9690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
rlabel metal1 3358 35156 3358 35156 0 Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
rlabel metal1 4462 34714 4462 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
rlabel metal2 9154 38250 9154 38250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
rlabel metal1 9338 37944 9338 37944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
rlabel metal1 13754 8058 13754 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
rlabel metal1 14444 8534 14444 8534 0 Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
rlabel metal2 12558 12070 12558 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
rlabel metal1 12466 12201 12466 12201 0 Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
rlabel metal1 3082 36618 3082 36618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
rlabel metal1 3818 36856 3818 36856 0 Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
rlabel metal1 8464 36550 8464 36550 0 Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
rlabel metal1 8602 35768 8602 35768 0 Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
rlabel metal2 13938 12070 13938 12070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
rlabel metal1 14812 12206 14812 12206 0 Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
rlabel metal2 11914 15130 11914 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
rlabel metal1 12190 14586 12190 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
rlabel metal2 3818 39916 3818 39916 0 Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
rlabel metal1 4462 39406 4462 39406 0 Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
rlabel metal2 7958 40154 7958 40154 0 Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
rlabel metal2 8418 39848 8418 39848 0 Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
rlabel metal1 13294 10506 13294 10506 0 Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
rlabel metal1 14582 10234 14582 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
rlabel metal1 11224 8058 11224 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
rlabel metal1 12190 8058 12190 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
rlabel metal1 2990 37740 2990 37740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
rlabel metal1 3910 37944 3910 37944 0 Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
rlabel metal2 9614 40426 9614 40426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
rlabel metal1 10028 39610 10028 39610 0 Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
rlabel metal1 13524 6970 13524 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
rlabel metal1 14214 6426 14214 6426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
rlabel metal1 10856 2618 10856 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
rlabel metal2 10350 3502 10350 3502 0 Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
rlabel metal2 3358 31076 3358 31076 0 Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
rlabel metal1 4922 30906 4922 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
rlabel metal2 5198 29852 5198 29852 0 Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
rlabel metal1 5796 29274 5796 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
rlabel metal2 11086 22950 11086 22950 0 Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
rlabel metal1 11132 23086 11132 23086 0 Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
rlabel metal2 6118 3162 6118 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
rlabel metal1 6900 2618 6900 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
rlabel metal1 6164 17034 6164 17034 0 Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
rlabel metal1 7222 17238 7222 17238 0 Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
rlabel metal1 9154 31654 9154 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
rlabel metal1 9522 30906 9522 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
rlabel metal2 12558 3740 12558 3740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
rlabel metal1 12834 3162 12834 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
rlabel metal2 12742 18666 12742 18666 0 Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
rlabel metal1 12190 18326 12190 18326 0 Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
rlabel metal1 2714 38794 2714 38794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
rlabel metal2 2346 39576 2346 39576 0 Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
rlabel metal2 10534 41015 10534 41015 0 Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
rlabel metal2 11086 40732 11086 40732 0 Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
rlabel metal1 13662 16660 13662 16660 0 Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
rlabel metal1 15042 16218 15042 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
rlabel metal2 8786 27302 8786 27302 0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 9614 27438 9614 27438 0 Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
rlabel metal1 2300 34714 2300 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
rlabel metal2 2714 35836 2714 35836 0 Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
rlabel metal2 12558 38624 12558 38624 0 Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
rlabel metal1 12880 37978 12880 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
rlabel metal1 14812 33014 14812 33014 0 Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
rlabel metal2 15318 33796 15318 33796 0 Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
rlabel metal2 9706 23834 9706 23834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
rlabel metal1 9476 22746 9476 22746 0 Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
rlabel metal1 2208 30158 2208 30158 0 Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 2714 30022 2714 30022 0 Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
rlabel metal1 2116 32334 2116 32334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
rlabel metal1 2530 31994 2530 31994 0 Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
rlabel metal1 7590 29784 7590 29784 0 Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
rlabel metal1 8280 29274 8280 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
rlabel metal1 2392 21658 2392 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
rlabel metal1 2300 21998 2300 21998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
rlabel metal2 2438 23766 2438 23766 0 Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
rlabel metal1 2254 24174 2254 24174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
rlabel metal1 2254 27302 2254 27302 0 Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
rlabel metal1 2530 26554 2530 26554 0 Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
rlabel metal2 8510 21284 8510 21284 0 Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
rlabel metal1 9430 21114 9430 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
rlabel metal2 9706 25194 9706 25194 0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
rlabel metal1 10350 25806 10350 25806 0 Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
rlabel metal1 10994 29138 10994 29138 0 Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
rlabel metal1 5612 36278 5612 36278 0 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
rlabel metal1 5980 35598 5980 35598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
rlabel metal1 7774 37230 7774 37230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
rlabel metal1 7452 34102 7452 34102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
rlabel metal2 8096 33490 8096 33490 0 Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
rlabel metal1 9338 34612 9338 34612 0 Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
rlabel metal2 16238 31518 16238 31518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
rlabel metal1 16882 31858 16882 31858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
rlabel metal1 17342 34612 17342 34612 0 Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
rlabel metal2 10994 20570 10994 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
rlabel metal1 10902 20026 10902 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
rlabel metal2 5566 33388 5566 33388 0 Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
rlabel metal1 5658 32878 5658 32878 0 Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
rlabel metal2 12834 35428 12834 35428 0 Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
rlabel metal1 12098 35768 12098 35768 0 Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
rlabel metal2 15134 32164 15134 32164 0 Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
rlabel metal2 14490 33694 14490 33694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
rlabel metal1 11270 22202 11270 22202 0 Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
rlabel metal2 12006 21794 12006 21794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
rlabel metal1 5842 27540 5842 27540 0 Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
rlabel metal1 6807 27370 6807 27370 0 Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
rlabel metal1 6808 31654 6808 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
rlabel metal1 7314 30906 7314 30906 0 Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
rlabel metal2 14950 29546 14950 29546 0 Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 14950 29206 14950 29206 0 Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
rlabel metal1 13064 18122 13064 18122 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
rlabel metal1 3174 33626 3174 33626 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
rlabel metal2 12374 38148 12374 38148 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
rlabel metal1 19619 18190 19619 18190 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
rlabel metal1 9430 23732 9430 23732 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
rlabel metal1 5026 7310 5026 7310 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
rlabel metal2 2346 32037 2346 32037 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
rlabel via1 16342 5746 16342 5746 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
rlabel metal2 2070 21199 2070 21199 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
rlabel metal2 6118 23970 6118 23970 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
rlabel metal2 2714 4998 2714 4998 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
rlabel metal1 8970 4046 8970 4046 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
rlabel via1 10454 9554 10454 9554 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
rlabel metal2 5290 35258 5290 35258 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
rlabel metal2 5796 20332 5796 20332 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
rlabel metal1 15594 29546 15594 29546 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
rlabel metal2 13386 14212 13386 14212 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
rlabel metal1 5762 24242 5762 24242 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
rlabel metal1 12650 33422 12650 33422 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
rlabel metal1 16928 8602 16928 8602 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
rlabel metal2 1058 19574 1058 19574 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
rlabel metal1 15686 16626 15686 16626 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
rlabel metal1 12558 12104 12558 12104 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
rlabel metal2 2714 17000 2714 17000 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
rlabel metal1 7832 16626 7832 16626 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
rlabel metal1 16284 14382 16284 14382 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
rlabel metal1 13202 25806 13202 25806 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
rlabel via1 4566 16082 4566 16082 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
rlabel via2 10442 27557 10442 27557 0 Inst_RAM_IO_switch_matrix.N1BEG0
rlabel metal2 3358 38148 3358 38148 0 Inst_RAM_IO_switch_matrix.N1BEG1
rlabel metal1 13018 42602 13018 42602 0 Inst_RAM_IO_switch_matrix.N1BEG2
rlabel metal1 16054 33082 16054 33082 0 Inst_RAM_IO_switch_matrix.N1BEG3
rlabel metal2 1150 27812 1150 27812 0 Inst_RAM_IO_switch_matrix.N2BEG0
rlabel metal2 1288 42092 1288 42092 0 Inst_RAM_IO_switch_matrix.N2BEG1
rlabel metal1 2576 42194 2576 42194 0 Inst_RAM_IO_switch_matrix.N2BEG2
rlabel metal1 8832 29818 8832 29818 0 Inst_RAM_IO_switch_matrix.N2BEG3
rlabel metal2 690 35896 690 35896 0 Inst_RAM_IO_switch_matrix.N2BEG4
rlabel metal2 414 32827 414 32827 0 Inst_RAM_IO_switch_matrix.N2BEG5
rlabel metal1 1610 41038 1610 41038 0 Inst_RAM_IO_switch_matrix.N2BEG6
rlabel metal1 9752 21658 9752 21658 0 Inst_RAM_IO_switch_matrix.N2BEG7
rlabel metal4 1012 22712 1012 22712 0 Inst_RAM_IO_switch_matrix.N2BEGb0
rlabel metal1 3818 31450 3818 31450 0 Inst_RAM_IO_switch_matrix.N2BEGb1
rlabel metal3 4163 34068 4163 34068 0 Inst_RAM_IO_switch_matrix.N2BEGb2
rlabel metal2 1012 27948 1012 27948 0 Inst_RAM_IO_switch_matrix.N2BEGb3
rlabel metal1 966 42670 966 42670 0 Inst_RAM_IO_switch_matrix.N2BEGb4
rlabel metal1 1288 19142 1288 19142 0 Inst_RAM_IO_switch_matrix.N2BEGb5
rlabel metal1 4968 31994 4968 31994 0 Inst_RAM_IO_switch_matrix.N2BEGb6
rlabel metal4 828 22440 828 22440 0 Inst_RAM_IO_switch_matrix.N2BEGb7
rlabel metal1 10626 42602 10626 42602 0 Inst_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 8648 37094 8648 37094 0 Inst_RAM_IO_switch_matrix.N4BEG1
rlabel metal2 9476 40188 9476 40188 0 Inst_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 16192 34714 16192 34714 0 Inst_RAM_IO_switch_matrix.N4BEG3
rlabel metal2 920 13124 920 13124 0 Inst_RAM_IO_switch_matrix.S1BEG0
rlabel metal2 18124 17238 18124 17238 0 Inst_RAM_IO_switch_matrix.S1BEG1
rlabel metal3 13133 2652 13133 2652 0 Inst_RAM_IO_switch_matrix.S1BEG2
rlabel metal3 21068 2448 21068 2448 0 Inst_RAM_IO_switch_matrix.S1BEG3
rlabel metal1 14306 2074 14306 2074 0 Inst_RAM_IO_switch_matrix.S2BEG0
rlabel via2 13294 2397 13294 2397 0 Inst_RAM_IO_switch_matrix.S2BEG1
rlabel via2 13570 1955 13570 1955 0 Inst_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 14628 2482 14628 2482 0 Inst_RAM_IO_switch_matrix.S2BEG3
rlabel metal2 14306 20230 14306 20230 0 Inst_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 14674 1870 14674 1870 0 Inst_RAM_IO_switch_matrix.S2BEG5
rlabel metal1 14582 18598 14582 18598 0 Inst_RAM_IO_switch_matrix.S2BEG6
rlabel metal2 15824 18598 15824 18598 0 Inst_RAM_IO_switch_matrix.S2BEG7
rlabel metal2 13846 2074 13846 2074 0 Inst_RAM_IO_switch_matrix.S2BEGb0
rlabel metal1 11362 2414 11362 2414 0 Inst_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 11546 2482 11546 2482 0 Inst_RAM_IO_switch_matrix.S2BEGb2
rlabel metal2 11546 1326 11546 1326 0 Inst_RAM_IO_switch_matrix.S2BEGb3
rlabel metal1 12282 2414 12282 2414 0 Inst_RAM_IO_switch_matrix.S2BEGb4
rlabel metal2 12466 15113 12466 15113 0 Inst_RAM_IO_switch_matrix.S2BEGb5
rlabel metal2 12466 24531 12466 24531 0 Inst_RAM_IO_switch_matrix.S2BEGb6
rlabel metal1 12880 1938 12880 1938 0 Inst_RAM_IO_switch_matrix.S2BEGb7
rlabel metal1 17158 7446 17158 7446 0 Inst_RAM_IO_switch_matrix.S4BEG0
rlabel metal3 18147 3740 18147 3740 0 Inst_RAM_IO_switch_matrix.S4BEG1
rlabel metal3 18952 18156 18952 18156 0 Inst_RAM_IO_switch_matrix.S4BEG2
rlabel metal1 19366 20774 19366 20774 0 Inst_RAM_IO_switch_matrix.S4BEG3
rlabel metal2 12650 5593 12650 5593 0 Inst_RAM_IO_switch_matrix.W1BEG0
rlabel metal2 6026 12580 6026 12580 0 Inst_RAM_IO_switch_matrix.W1BEG1
rlabel metal1 8602 11050 8602 11050 0 Inst_RAM_IO_switch_matrix.W1BEG2
rlabel metal1 14582 4658 14582 4658 0 Inst_RAM_IO_switch_matrix.W1BEG3
rlabel metal1 4278 6698 4278 6698 0 Inst_RAM_IO_switch_matrix.W2BEG0
rlabel metal1 6026 5338 6026 5338 0 Inst_RAM_IO_switch_matrix.W2BEG1
rlabel metal1 5612 6290 5612 6290 0 Inst_RAM_IO_switch_matrix.W2BEG2
rlabel metal1 8372 6290 8372 6290 0 Inst_RAM_IO_switch_matrix.W2BEG3
rlabel metal2 16606 5117 16606 5117 0 Inst_RAM_IO_switch_matrix.W2BEG4
rlabel metal1 4278 7888 4278 7888 0 Inst_RAM_IO_switch_matrix.W2BEG5
rlabel metal1 4416 4114 4416 4114 0 Inst_RAM_IO_switch_matrix.W2BEG6
rlabel metal1 2530 3060 2530 3060 0 Inst_RAM_IO_switch_matrix.W2BEG7
rlabel metal1 7958 6154 7958 6154 0 Inst_RAM_IO_switch_matrix.W2BEGb0
rlabel metal1 2806 7276 2806 7276 0 Inst_RAM_IO_switch_matrix.W2BEGb1
rlabel metal1 3818 8942 3818 8942 0 Inst_RAM_IO_switch_matrix.W2BEGb2
rlabel metal1 7728 8058 7728 8058 0 Inst_RAM_IO_switch_matrix.W2BEGb3
rlabel metal1 8418 5576 8418 5576 0 Inst_RAM_IO_switch_matrix.W2BEGb4
rlabel metal3 3450 11492 3450 11492 0 Inst_RAM_IO_switch_matrix.W2BEGb5
rlabel metal1 1702 4522 1702 4522 0 Inst_RAM_IO_switch_matrix.W2BEGb6
rlabel via2 2714 3485 2714 3485 0 Inst_RAM_IO_switch_matrix.W2BEGb7
rlabel metal1 8418 14280 8418 14280 0 Inst_RAM_IO_switch_matrix.W6BEG0
rlabel metal1 1518 39032 1518 39032 0 Inst_RAM_IO_switch_matrix.W6BEG1
rlabel metal1 3266 19380 3266 19380 0 Inst_RAM_IO_switch_matrix.W6BEG10
rlabel metal1 11684 17646 11684 17646 0 Inst_RAM_IO_switch_matrix.W6BEG11
rlabel metal1 2185 36822 2185 36822 0 Inst_RAM_IO_switch_matrix.W6BEG2
rlabel metal1 6668 15402 6668 15402 0 Inst_RAM_IO_switch_matrix.W6BEG3
rlabel via2 17802 14467 17802 14467 0 Inst_RAM_IO_switch_matrix.W6BEG4
rlabel metal2 1794 14671 1794 14671 0 Inst_RAM_IO_switch_matrix.W6BEG5
rlabel metal1 4508 16218 4508 16218 0 Inst_RAM_IO_switch_matrix.W6BEG6
rlabel metal1 10718 15674 10718 15674 0 Inst_RAM_IO_switch_matrix.W6BEG7
rlabel metal1 17664 16558 17664 16558 0 Inst_RAM_IO_switch_matrix.W6BEG8
rlabel metal1 6808 16762 6808 16762 0 Inst_RAM_IO_switch_matrix.W6BEG9
rlabel metal1 13386 6936 13386 6936 0 Inst_RAM_IO_switch_matrix.WW4BEG0
rlabel metal1 2070 13906 2070 13906 0 Inst_RAM_IO_switch_matrix.WW4BEG1
rlabel metal1 1610 17238 1610 17238 0 Inst_RAM_IO_switch_matrix.WW4BEG10
rlabel metal2 9522 13124 9522 13124 0 Inst_RAM_IO_switch_matrix.WW4BEG11
rlabel metal1 15962 7718 15962 7718 0 Inst_RAM_IO_switch_matrix.WW4BEG12
rlabel metal1 4094 14382 4094 14382 0 Inst_RAM_IO_switch_matrix.WW4BEG13
rlabel metal1 4232 7514 4232 7514 0 Inst_RAM_IO_switch_matrix.WW4BEG14
rlabel metal2 11270 10166 11270 10166 0 Inst_RAM_IO_switch_matrix.WW4BEG15
rlabel metal1 1702 9962 1702 9962 0 Inst_RAM_IO_switch_matrix.WW4BEG2
rlabel metal2 1610 9571 1610 9571 0 Inst_RAM_IO_switch_matrix.WW4BEG3
rlabel metal1 7314 11152 7314 11152 0 Inst_RAM_IO_switch_matrix.WW4BEG4
rlabel metal1 5658 11186 5658 11186 0 Inst_RAM_IO_switch_matrix.WW4BEG5
rlabel metal2 2116 11492 2116 11492 0 Inst_RAM_IO_switch_matrix.WW4BEG6
rlabel metal1 9338 13192 9338 13192 0 Inst_RAM_IO_switch_matrix.WW4BEG7
rlabel metal2 16606 11849 16606 11849 0 Inst_RAM_IO_switch_matrix.WW4BEG8
rlabel metal2 7590 10370 7590 10370 0 Inst_RAM_IO_switch_matrix.WW4BEG9
rlabel metal1 10810 25738 10810 25738 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
rlabel metal1 11040 26554 11040 26554 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
rlabel metal1 11086 28492 11086 28492 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 11546 28560 11546 28560 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 11178 28866 11178 28866 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
rlabel metal1 11178 29070 11178 29070 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
rlabel metal1 6440 35802 6440 35802 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
rlabel metal1 7038 36142 7038 36142 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
rlabel metal1 6992 36346 6992 36346 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 7728 36550 7728 36550 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7544 36890 7544 36890 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
rlabel metal1 8326 37298 8326 37298 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
rlabel metal1 9338 33456 9338 33456 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
rlabel metal1 8878 33490 8878 33490 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
rlabel metal1 9338 33626 9338 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 8878 33592 8878 33592 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 8970 34374 8970 34374 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
rlabel metal1 9108 34510 9108 34510 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
rlabel metal1 17296 31994 17296 31994 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
rlabel metal1 17480 29818 17480 29818 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
rlabel metal1 17020 33626 17020 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 17434 34170 17434 34170 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 16974 34442 16974 34442 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
rlabel metal1 17204 34510 17204 34510 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
rlabel metal1 14950 27438 14950 27438 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
rlabel metal1 15226 25874 15226 25874 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
rlabel metal1 15594 25908 15594 25908 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 16054 25840 16054 25840 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 15686 26180 15686 26180 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
rlabel metal1 16468 26010 16468 26010 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
rlabel metal1 7130 24174 7130 24174 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
rlabel metal1 7774 24174 7774 24174 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
rlabel metal1 7498 24242 7498 24242 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 8510 23732 8510 23732 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 7866 23120 7866 23120 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
rlabel metal1 8326 23086 8326 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
rlabel metal1 12558 30702 12558 30702 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
rlabel metal1 13018 30634 13018 30634 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
rlabel metal1 12834 31790 12834 31790 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 13386 30906 13386 30906 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 13386 31654 13386 31654 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
rlabel metal1 14950 30736 14950 30736 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
rlabel metal1 18492 21998 18492 21998 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
rlabel metal1 18676 21522 18676 21522 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
rlabel metal1 18446 21862 18446 21862 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 19458 20944 19458 20944 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 18722 20944 18722 20944 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
rlabel metal1 19228 20842 19228 20842 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
rlabel metal2 230 44193 230 44193 0 N1BEG[0]
rlabel metal2 506 43428 506 43428 0 N1BEG[1]
rlabel metal2 782 43156 782 43156 0 N1BEG[2]
rlabel metal2 1058 43258 1058 43258 0 N1BEG[3]
rlabel metal2 329 68 329 68 0 N1END[0]
rlabel metal2 506 1146 506 1146 0 N1END[1]
rlabel metal2 835 68 835 68 0 N1END[2]
rlabel metal1 1564 3094 1564 3094 0 N1END[3]
rlabel metal2 1334 43632 1334 43632 0 N2BEG[0]
rlabel metal2 1610 42986 1610 42986 0 N2BEG[1]
rlabel metal2 1886 43972 1886 43972 0 N2BEG[2]
rlabel metal2 2162 44057 2162 44057 0 N2BEG[3]
rlabel metal1 2668 41786 2668 41786 0 N2BEG[4]
rlabel metal2 2714 43581 2714 43581 0 N2BEG[5]
rlabel metal1 2898 43418 2898 43418 0 N2BEG[6]
rlabel metal2 3266 44057 3266 44057 0 N2BEG[7]
rlabel metal1 3266 42058 3266 42058 0 N2BEGb[0]
rlabel metal1 4002 42330 4002 42330 0 N2BEGb[1]
rlabel metal2 4094 43802 4094 43802 0 N2BEGb[2]
rlabel metal2 4370 43972 4370 43972 0 N2BEGb[3]
rlabel metal1 4692 42534 4692 42534 0 N2BEGb[4]
rlabel metal2 4922 43632 4922 43632 0 N2BEGb[5]
rlabel metal1 5106 42330 5106 42330 0 N2BEGb[6]
rlabel metal2 5474 44193 5474 44193 0 N2BEGb[7]
rlabel metal2 3641 68 3641 68 0 N2END[0]
rlabel metal2 3818 704 3818 704 0 N2END[1]
rlabel metal2 3995 68 3995 68 0 N2END[2]
rlabel metal2 4423 68 4423 68 0 N2END[3]
rlabel metal2 4593 68 4593 68 0 N2END[4]
rlabel metal2 4922 534 4922 534 0 N2END[5]
rlabel metal2 5251 68 5251 68 0 N2END[6]
rlabel metal2 5474 755 5474 755 0 N2END[7]
rlabel metal2 1334 755 1334 755 0 N2MID[0]
rlabel metal2 1709 68 1709 68 0 N2MID[1]
rlabel metal2 1985 68 1985 68 0 N2MID[2]
rlabel metal2 2261 68 2261 68 0 N2MID[3]
rlabel metal2 2438 398 2438 398 0 N2MID[4]
rlabel metal2 2714 1214 2714 1214 0 N2MID[5]
rlabel metal2 3043 68 3043 68 0 N2MID[6]
rlabel metal2 3266 1010 3266 1010 0 N2MID[7]
rlabel metal2 5750 43530 5750 43530 0 N4BEG[0]
rlabel metal1 8418 43418 8418 43418 0 N4BEG[10]
rlabel metal1 8740 42738 8740 42738 0 N4BEG[11]
rlabel metal1 8878 43418 8878 43418 0 N4BEG[12]
rlabel metal2 9338 43632 9338 43632 0 N4BEG[13]
rlabel metal1 9430 43418 9430 43418 0 N4BEG[14]
rlabel metal1 9844 43418 9844 43418 0 N4BEG[15]
rlabel metal2 6026 44057 6026 44057 0 N4BEG[1]
rlabel metal1 6210 43418 6210 43418 0 N4BEG[2]
rlabel metal2 6578 43921 6578 43921 0 N4BEG[3]
rlabel metal2 6854 44465 6854 44465 0 N4BEG[4]
rlabel metal2 7130 44125 7130 44125 0 N4BEG[5]
rlabel metal1 7728 42534 7728 42534 0 N4BEG[6]
rlabel metal1 7544 43418 7544 43418 0 N4BEG[7]
rlabel metal1 7866 43418 7866 43418 0 N4BEG[8]
rlabel metal2 8234 43428 8234 43428 0 N4BEG[9]
rlabel metal4 1196 22032 1196 22032 0 N4BEG_outbuf_0.A
rlabel metal2 5658 41820 5658 41820 0 N4BEG_outbuf_0.X
rlabel metal4 2484 12420 2484 12420 0 N4BEG_outbuf_1.A
rlabel metal1 6394 41616 6394 41616 0 N4BEG_outbuf_1.X
rlabel via2 9522 2635 9522 2635 0 N4BEG_outbuf_10.A
rlabel metal2 9154 42262 9154 42262 0 N4BEG_outbuf_10.X
rlabel metal2 8694 1411 8694 1411 0 N4BEG_outbuf_11.A
rlabel metal1 10166 42160 10166 42160 0 N4BEG_outbuf_11.X
rlabel metal3 6463 1156 6463 1156 0 N4BEG_outbuf_2.A
rlabel metal1 5382 41548 5382 41548 0 N4BEG_outbuf_2.X
rlabel metal2 12696 2108 12696 2108 0 N4BEG_outbuf_3.A
rlabel metal1 5888 41582 5888 41582 0 N4BEG_outbuf_3.X
rlabel metal2 7314 2210 7314 2210 0 N4BEG_outbuf_4.A
rlabel metal1 6164 42330 6164 42330 0 N4BEG_outbuf_4.X
rlabel via2 7958 1309 7958 1309 0 N4BEG_outbuf_5.A
rlabel metal1 7176 41582 7176 41582 0 N4BEG_outbuf_5.X
rlabel metal1 7728 2074 7728 2074 0 N4BEG_outbuf_6.A
rlabel metal1 7774 41616 7774 41616 0 N4BEG_outbuf_6.X
rlabel metal1 8096 2074 8096 2074 0 N4BEG_outbuf_7.A
rlabel metal1 8050 41650 8050 41650 0 N4BEG_outbuf_7.X
rlabel metal2 8418 2159 8418 2159 0 N4BEG_outbuf_8.A
rlabel metal1 8326 41684 8326 41684 0 N4BEG_outbuf_8.X
rlabel metal1 8832 2074 8832 2074 0 N4BEG_outbuf_9.A
rlabel metal2 7958 41253 7958 41253 0 N4BEG_outbuf_9.X
rlabel metal2 5750 670 5750 670 0 N4END[0]
rlabel metal2 8510 211 8510 211 0 N4END[10]
rlabel metal2 8786 143 8786 143 0 N4END[11]
rlabel metal2 9161 68 9161 68 0 N4END[12]
rlabel metal1 7590 2482 7590 2482 0 N4END[13]
rlabel metal2 9515 68 9515 68 0 N4END[14]
rlabel metal2 9890 704 9890 704 0 N4END[15]
rlabel metal2 6026 704 6026 704 0 N4END[1]
rlabel metal2 6355 68 6355 68 0 N4END[2]
rlabel metal2 6525 68 6525 68 0 N4END[3]
rlabel metal2 6755 68 6755 68 0 N4END[4]
rlabel metal2 7130 534 7130 534 0 N4END[5]
rlabel metal2 7406 1248 7406 1248 0 N4END[6]
rlabel metal2 7682 755 7682 755 0 N4END[7]
rlabel metal2 7958 619 7958 619 0 N4END[8]
rlabel metal2 8234 1180 8234 1180 0 N4END[9]
rlabel metal3 24836 7140 24836 7140 0 RAM2FAB_D0_I0
rlabel metal3 25572 7684 25572 7684 0 RAM2FAB_D0_I1
rlabel metal3 25204 8228 25204 8228 0 RAM2FAB_D0_I2
rlabel metal3 25503 8772 25503 8772 0 RAM2FAB_D0_I3
rlabel metal3 24951 4964 24951 4964 0 RAM2FAB_D1_I0
rlabel metal3 25802 5508 25802 5508 0 RAM2FAB_D1_I1
rlabel metal3 24790 6052 24790 6052 0 RAM2FAB_D1_I2
rlabel metal3 20884 6528 20884 6528 0 RAM2FAB_D1_I3
rlabel metal3 24284 2788 24284 2788 0 RAM2FAB_D2_I0
rlabel metal2 21298 3859 21298 3859 0 RAM2FAB_D2_I1
rlabel metal2 21482 4573 21482 4573 0 RAM2FAB_D2_I2
rlabel metal1 22034 4556 22034 4556 0 RAM2FAB_D2_I3
rlabel metal1 20286 3910 20286 3910 0 RAM2FAB_D3_I0
rlabel metal2 21068 5678 21068 5678 0 RAM2FAB_D3_I1
rlabel via2 21390 1411 21390 1411 0 RAM2FAB_D3_I2
rlabel metal1 17710 3026 17710 3026 0 RAM2FAB_D3_I3
rlabel metal2 10166 347 10166 347 0 S1BEG[0]
rlabel metal2 10495 68 10495 68 0 S1BEG[1]
rlabel metal2 10718 636 10718 636 0 S1BEG[2]
rlabel metal2 10994 908 10994 908 0 S1BEG[3]
rlabel metal2 10166 43904 10166 43904 0 S1END[0]
rlabel metal2 10442 43904 10442 43904 0 S1END[1]
rlabel metal2 10718 43904 10718 43904 0 S1END[2]
rlabel metal2 10994 43904 10994 43904 0 S1END[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 806 13754 806 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14306 908 14306 908 0 S2BEG[3]
rlabel metal2 14582 908 14582 908 0 S2BEG[4]
rlabel metal2 14858 806 14858 806 0 S2BEG[5]
rlabel metal2 15134 755 15134 755 0 S2BEG[6]
rlabel metal2 15410 942 15410 942 0 S2BEG[7]
rlabel metal2 11217 68 11217 68 0 S2BEGb[0]
rlabel metal2 11546 398 11546 398 0 S2BEGb[1]
rlabel metal2 11822 483 11822 483 0 S2BEGb[2]
rlabel metal2 12098 364 12098 364 0 S2BEGb[3]
rlabel metal2 12374 636 12374 636 0 S2BEGb[4]
rlabel metal2 12650 908 12650 908 0 S2BEGb[5]
rlabel metal2 12926 347 12926 347 0 S2BEGb[6]
rlabel metal2 13202 636 13202 636 0 S2BEGb[7]
rlabel metal2 11270 43904 11270 43904 0 S2END[0]
rlabel metal2 11546 44057 11546 44057 0 S2END[1]
rlabel metal2 11822 44329 11822 44329 0 S2END[2]
rlabel metal2 12098 43904 12098 43904 0 S2END[3]
rlabel metal2 12374 43938 12374 43938 0 S2END[4]
rlabel metal2 12650 43938 12650 43938 0 S2END[5]
rlabel metal2 12926 44125 12926 44125 0 S2END[6]
rlabel metal2 13202 44193 13202 44193 0 S2END[7]
rlabel metal2 13478 43938 13478 43938 0 S2MID[0]
rlabel metal2 13754 43632 13754 43632 0 S2MID[1]
rlabel metal2 14030 44057 14030 44057 0 S2MID[2]
rlabel metal2 14306 44057 14306 44057 0 S2MID[3]
rlabel metal2 14582 43938 14582 43938 0 S2MID[4]
rlabel metal2 14858 43938 14858 43938 0 S2MID[5]
rlabel metal2 15134 43632 15134 43632 0 S2MID[6]
rlabel metal2 15410 43938 15410 43938 0 S2MID[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18446 1180 18446 1180 0 S4BEG[10]
rlabel metal2 18722 534 18722 534 0 S4BEG[11]
rlabel metal2 19097 68 19097 68 0 S4BEG[12]
rlabel metal2 19274 1027 19274 1027 0 S4BEG[13]
rlabel metal2 19550 891 19550 891 0 S4BEG[14]
rlabel metal2 19925 68 19925 68 0 S4BEG[15]
rlabel metal2 15962 772 15962 772 0 S4BEG[1]
rlabel metal1 17526 1428 17526 1428 0 S4BEG[2]
rlabel metal2 16698 1343 16698 1343 0 S4BEG[3]
rlabel metal2 16843 68 16843 68 0 S4BEG[4]
rlabel metal2 17066 1350 17066 1350 0 S4BEG[5]
rlabel metal2 17395 68 17395 68 0 S4BEG[6]
rlabel metal2 17618 908 17618 908 0 S4BEG[7]
rlabel metal2 17894 772 17894 772 0 S4BEG[8]
rlabel metal2 18223 68 18223 68 0 S4BEG[9]
rlabel metal1 16606 42194 16606 42194 0 S4BEG_outbuf_0.A
rlabel via3 16491 1292 16491 1292 0 S4BEG_outbuf_0.X
rlabel metal1 16790 42296 16790 42296 0 S4BEG_outbuf_1.A
rlabel via2 16422 2397 16422 2397 0 S4BEG_outbuf_1.X
rlabel metal1 19366 40528 19366 40528 0 S4BEG_outbuf_10.A
rlabel metal2 19228 17238 19228 17238 0 S4BEG_outbuf_10.X
rlabel metal1 19458 40086 19458 40086 0 S4BEG_outbuf_11.A
rlabel metal2 18400 8262 18400 8262 0 S4BEG_outbuf_11.X
rlabel metal1 17250 42262 17250 42262 0 S4BEG_outbuf_2.A
rlabel metal1 17020 2482 17020 2482 0 S4BEG_outbuf_2.X
rlabel metal1 17664 42262 17664 42262 0 S4BEG_outbuf_3.A
rlabel metal3 17319 2652 17319 2652 0 S4BEG_outbuf_3.X
rlabel metal1 17986 42262 17986 42262 0 S4BEG_outbuf_4.A
rlabel metal1 24702 41582 24702 41582 0 S4BEG_outbuf_4.X
rlabel metal1 18262 42296 18262 42296 0 S4BEG_outbuf_5.A
rlabel via3 18515 2652 18515 2652 0 S4BEG_outbuf_5.X
rlabel metal2 18630 42398 18630 42398 0 S4BEG_outbuf_6.A
rlabel metal3 19527 2652 19527 2652 0 S4BEG_outbuf_6.X
rlabel metal1 18906 42262 18906 42262 0 S4BEG_outbuf_7.A
rlabel metal2 18492 37468 18492 37468 0 S4BEG_outbuf_7.X
rlabel metal1 18308 41582 18308 41582 0 S4BEG_outbuf_8.A
rlabel metal3 18193 41412 18193 41412 0 S4BEG_outbuf_8.X
rlabel metal1 19458 42262 19458 42262 0 S4BEG_outbuf_9.A
rlabel metal2 19274 7888 19274 7888 0 S4BEG_outbuf_9.X
rlabel metal2 15686 43904 15686 43904 0 S4END[0]
rlabel metal2 18446 44193 18446 44193 0 S4END[10]
rlabel metal2 18722 44125 18722 44125 0 S4END[11]
rlabel metal2 18998 44125 18998 44125 0 S4END[12]
rlabel metal1 19964 40426 19964 40426 0 S4END[13]
rlabel metal2 19550 43938 19550 43938 0 S4END[14]
rlabel metal2 19090 42279 19090 42279 0 S4END[15]
rlabel metal2 15962 43938 15962 43938 0 S4END[1]
rlabel metal2 16238 43938 16238 43938 0 S4END[2]
rlabel metal2 16514 43649 16514 43649 0 S4END[3]
rlabel metal2 16790 43938 16790 43938 0 S4END[4]
rlabel metal2 17066 43972 17066 43972 0 S4END[5]
rlabel metal2 17342 44261 17342 44261 0 S4END[6]
rlabel metal2 17618 43921 17618 43921 0 S4END[7]
rlabel metal2 17894 43989 17894 43989 0 S4END[8]
rlabel metal2 18170 44057 18170 44057 0 S4END[9]
rlabel metal1 19274 17578 19274 17578 0 UserCLK
rlabel metal2 20746 41939 20746 41939 0 UserCLKo
rlabel metal3 774 4964 774 4964 0 W1BEG[0]
rlabel metal2 2898 5389 2898 5389 0 W1BEG[1]
rlabel metal3 567 5508 567 5508 0 W1BEG[2]
rlabel metal3 728 5780 728 5780 0 W1BEG[3]
rlabel metal3 866 6052 866 6052 0 W2BEG[0]
rlabel metal3 728 6324 728 6324 0 W2BEG[1]
rlabel metal3 590 6596 590 6596 0 W2BEG[2]
rlabel metal3 682 6868 682 6868 0 W2BEG[3]
rlabel metal2 3542 6783 3542 6783 0 W2BEG[4]
rlabel metal3 958 7412 958 7412 0 W2BEG[5]
rlabel metal3 912 7684 912 7684 0 W2BEG[6]
rlabel metal2 3358 8143 3358 8143 0 W2BEG[7]
rlabel metal3 774 8228 774 8228 0 W2BEGb[0]
rlabel metal3 728 8500 728 8500 0 W2BEGb[1]
rlabel metal3 866 8772 866 8772 0 W2BEGb[2]
rlabel metal3 590 9044 590 9044 0 W2BEGb[3]
rlabel metal3 498 9316 498 9316 0 W2BEGb[4]
rlabel metal3 682 9588 682 9588 0 W2BEGb[5]
rlabel metal3 958 9860 958 9860 0 W2BEGb[6]
rlabel metal2 3082 10557 3082 10557 0 W2BEGb[7]
rlabel metal3 475 14756 475 14756 0 W6BEG[0]
rlabel metal3 958 17476 958 17476 0 W6BEG[10]
rlabel metal3 866 17748 866 17748 0 W6BEG[11]
rlabel metal3 659 15028 659 15028 0 W6BEG[1]
rlabel metal3 774 15300 774 15300 0 W6BEG[2]
rlabel metal2 3082 15181 3082 15181 0 W6BEG[3]
rlabel metal3 912 15844 912 15844 0 W6BEG[4]
rlabel metal2 3082 16269 3082 16269 0 W6BEG[5]
rlabel metal3 1418 16388 1418 16388 0 W6BEG[6]
rlabel metal2 2898 16167 2898 16167 0 W6BEG[7]
rlabel metal3 590 16932 590 16932 0 W6BEG[8]
rlabel metal2 3358 16983 3358 16983 0 W6BEG[9]
rlabel metal2 2898 9078 2898 9078 0 WW4BEG[0]
rlabel metal3 682 13124 682 13124 0 WW4BEG[10]
rlabel metal3 751 13396 751 13396 0 WW4BEG[11]
rlabel via2 3818 13685 3818 13685 0 WW4BEG[12]
rlabel metal3 774 13940 774 13940 0 WW4BEG[13]
rlabel metal3 958 14212 958 14212 0 WW4BEG[14]
rlabel metal2 2806 13991 2806 13991 0 WW4BEG[15]
rlabel metal2 4002 10829 4002 10829 0 WW4BEG[1]
rlabel metal3 912 10948 912 10948 0 WW4BEG[2]
rlabel metal2 3634 11271 3634 11271 0 WW4BEG[3]
rlabel metal1 1840 8058 1840 8058 0 WW4BEG[4]
rlabel metal2 3174 11509 3174 11509 0 WW4BEG[5]
rlabel metal3 774 12036 774 12036 0 WW4BEG[6]
rlabel metal2 3726 12189 3726 12189 0 WW4BEG[7]
rlabel metal3 406 12580 406 12580 0 WW4BEG[8]
rlabel metal3 1234 12852 1234 12852 0 WW4BEG[9]
rlabel metal1 23276 26554 23276 26554 0 data_inbuf_0.X
rlabel metal1 23782 27642 23782 27642 0 data_inbuf_1.X
rlabel metal1 21965 32266 21965 32266 0 data_inbuf_10.X
rlabel metal1 23598 32470 23598 32470 0 data_inbuf_11.X
rlabel metal1 23046 32946 23046 32946 0 data_inbuf_12.X
rlabel metal1 23552 33966 23552 33966 0 data_inbuf_13.X
rlabel metal1 23414 34646 23414 34646 0 data_inbuf_14.X
rlabel metal1 18998 34714 18998 34714 0 data_inbuf_15.X
rlabel metal1 22034 35632 22034 35632 0 data_inbuf_16.X
rlabel metal1 23322 35598 23322 35598 0 data_inbuf_17.X
rlabel metal1 21850 36108 21850 36108 0 data_inbuf_18.X
rlabel metal1 19826 36722 19826 36722 0 data_inbuf_19.X
rlabel metal1 23690 28016 23690 28016 0 data_inbuf_2.X
rlabel metal1 21114 36720 21114 36720 0 data_inbuf_20.X
rlabel metal1 23230 37094 23230 37094 0 data_inbuf_21.X
rlabel metal1 23000 37434 23000 37434 0 data_inbuf_22.X
rlabel metal1 22080 37434 22080 37434 0 data_inbuf_23.X
rlabel metal1 20286 38522 20286 38522 0 data_inbuf_24.X
rlabel metal1 23046 39338 23046 39338 0 data_inbuf_25.X
rlabel metal2 21114 39916 21114 39916 0 data_inbuf_26.X
rlabel metal1 20516 40494 20516 40494 0 data_inbuf_27.X
rlabel metal1 20194 41616 20194 41616 0 data_inbuf_28.X
rlabel metal1 23138 39984 23138 39984 0 data_inbuf_29.X
rlabel metal1 23690 28492 23690 28492 0 data_inbuf_3.X
rlabel metal2 21390 39780 21390 39780 0 data_inbuf_30.X
rlabel metal1 20512 40018 20512 40018 0 data_inbuf_31.X
rlabel metal1 23874 29172 23874 29172 0 data_inbuf_4.X
rlabel metal1 23736 29614 23736 29614 0 data_inbuf_5.X
rlabel metal1 23966 30192 23966 30192 0 data_inbuf_6.X
rlabel metal1 23690 30804 23690 30804 0 data_inbuf_7.X
rlabel metal1 23138 31280 23138 31280 0 data_inbuf_8.X
rlabel metal1 21390 31824 21390 31824 0 data_inbuf_9.X
rlabel metal1 24150 26928 24150 26928 0 data_outbuf_0.X
rlabel metal1 23506 26996 23506 26996 0 data_outbuf_1.X
rlabel metal1 23138 32402 23138 32402 0 data_outbuf_10.X
rlabel metal1 23874 32368 23874 32368 0 data_outbuf_11.X
rlabel metal1 23092 32742 23092 32742 0 data_outbuf_12.X
rlabel metal1 23368 33966 23368 33966 0 data_outbuf_13.X
rlabel metal1 23230 34476 23230 34476 0 data_outbuf_14.X
rlabel metal1 21022 35088 21022 35088 0 data_outbuf_15.X
rlabel metal1 22586 35734 22586 35734 0 data_outbuf_16.X
rlabel metal1 23092 35802 23092 35802 0 data_outbuf_17.X
rlabel metal1 21873 36006 21873 36006 0 data_outbuf_18.X
rlabel metal1 20838 36788 20838 36788 0 data_outbuf_19.X
rlabel viali 23414 28049 23414 28049 0 data_outbuf_2.X
rlabel metal1 21390 36890 21390 36890 0 data_outbuf_20.X
rlabel metal1 23782 39066 23782 39066 0 data_outbuf_21.X
rlabel metal1 23644 38522 23644 38522 0 data_outbuf_22.X
rlabel metal1 23414 38454 23414 38454 0 data_outbuf_23.X
rlabel metal2 20470 39168 20470 39168 0 data_outbuf_24.X
rlabel metal2 22862 39491 22862 39491 0 data_outbuf_25.X
rlabel metal1 20286 40086 20286 40086 0 data_outbuf_26.X
rlabel metal2 20286 40477 20286 40477 0 data_outbuf_27.X
rlabel metal2 21390 41633 21390 41633 0 data_outbuf_28.X
rlabel metal1 22034 40460 22034 40460 0 data_outbuf_29.X
rlabel metal1 23276 28526 23276 28526 0 data_outbuf_3.X
rlabel metal1 23414 40086 23414 40086 0 data_outbuf_30.X
rlabel metal1 22586 39950 22586 39950 0 data_outbuf_31.X
rlabel metal1 23598 29070 23598 29070 0 data_outbuf_4.X
rlabel metal1 23552 29614 23552 29614 0 data_outbuf_5.X
rlabel metal1 23828 30362 23828 30362 0 data_outbuf_6.X
rlabel metal1 23046 30736 23046 30736 0 data_outbuf_7.X
rlabel metal1 23598 31314 23598 31314 0 data_outbuf_8.X
rlabel metal1 21712 31790 21712 31790 0 data_outbuf_9.X
rlabel metal1 11822 17714 11822 17714 0 net1
rlabel metal1 7406 21522 7406 21522 0 net10
rlabel metal1 19182 19380 19182 19380 0 net100
rlabel metal1 2024 2550 2024 2550 0 net101
rlabel metal1 2070 2618 2070 2618 0 net102
rlabel metal3 10787 13668 10787 13668 0 net103
rlabel metal1 2254 3060 2254 3060 0 net104
rlabel metal1 4002 2074 4002 2074 0 net105
rlabel metal4 644 14688 644 14688 0 net106
rlabel metal2 368 12420 368 12420 0 net107
rlabel metal1 5152 2618 5152 2618 0 net108
rlabel metal2 3450 1088 3450 1088 0 net109
rlabel metal1 2576 29478 2576 29478 0 net11
rlabel metal1 5474 1802 5474 1802 0 net110
rlabel via3 5589 1292 5589 1292 0 net111
rlabel metal1 12696 3434 12696 3434 0 net112
rlabel metal1 2346 1734 2346 1734 0 net113
rlabel metal2 2070 7956 2070 7956 0 net114
rlabel metal2 2806 1088 2806 1088 0 net115
rlabel metal2 736 18428 736 18428 0 net116
rlabel metal1 2484 1530 2484 1530 0 net117
rlabel metal1 4554 2550 4554 2550 0 net118
rlabel metal1 3266 1224 3266 1224 0 net119
rlabel via2 9614 23715 9614 23715 0 net12
rlabel metal1 10902 3536 10902 3536 0 net120
rlabel metal1 5152 1190 5152 1190 0 net121
rlabel metal1 7590 1904 7590 1904 0 net122
rlabel metal1 8234 2006 8234 2006 0 net123
rlabel metal2 9154 2516 9154 2516 0 net124
rlabel metal2 8694 2193 8694 2193 0 net125
rlabel metal1 8556 1190 8556 1190 0 net126
rlabel metal1 8740 1326 8740 1326 0 net127
rlabel metal1 13110 24616 13110 24616 0 net128
rlabel metal2 6578 1241 6578 1241 0 net129
rlabel metal1 14168 18802 14168 18802 0 net13
rlabel metal2 12742 12886 12742 12886 0 net130
rlabel metal1 5566 2006 5566 2006 0 net131
rlabel metal1 6486 2040 6486 2040 0 net132
rlabel metal1 7268 1326 7268 1326 0 net133
rlabel metal1 6762 2006 6762 2006 0 net134
rlabel metal1 7130 1972 7130 1972 0 net135
rlabel metal1 8050 1258 8050 1258 0 net136
rlabel metal1 20930 6732 20930 6732 0 net137
rlabel metal1 20608 10030 20608 10030 0 net138
rlabel metal1 24518 7446 24518 7446 0 net139
rlabel metal1 1932 18394 1932 18394 0 net14
rlabel metal1 22540 8806 22540 8806 0 net140
rlabel metal1 18998 6766 18998 6766 0 net141
rlabel metal2 21666 9180 21666 9180 0 net142
rlabel metal1 21758 6970 21758 6970 0 net143
rlabel metal1 21574 6290 21574 6290 0 net144
rlabel metal1 19550 3128 19550 3128 0 net145
rlabel metal2 20378 5236 20378 5236 0 net146
rlabel metal1 18533 10642 18533 10642 0 net147
rlabel metal1 20603 12818 20603 12818 0 net148
rlabel metal1 17894 4012 17894 4012 0 net149
rlabel metal1 5566 21930 5566 21930 0 net15
rlabel metal2 21206 7072 21206 7072 0 net150
rlabel metal1 19642 2448 19642 2448 0 net151
rlabel metal1 17710 2924 17710 2924 0 net152
rlabel metal2 21666 19856 21666 19856 0 net153
rlabel metal2 3404 19822 3404 19822 0 net154
rlabel metal1 9200 19414 9200 19414 0 net155
rlabel metal1 14214 16422 14214 16422 0 net156
rlabel metal3 11408 11084 11408 11084 0 net157
rlabel metal3 6049 31212 6049 31212 0 net158
rlabel metal1 8878 38250 8878 38250 0 net159
rlabel metal2 1610 19635 1610 19635 0 net16
rlabel metal3 11477 24684 11477 24684 0 net160
rlabel via3 12581 42908 12581 42908 0 net161
rlabel metal2 12650 31824 12650 31824 0 net162
rlabel metal1 12834 42738 12834 42738 0 net163
rlabel metal3 14375 42908 14375 42908 0 net164
rlabel via3 13869 42908 13869 42908 0 net165
rlabel metal2 14950 42534 14950 42534 0 net166
rlabel metal2 13432 36516 13432 36516 0 net167
rlabel metal1 12098 23698 12098 23698 0 net168
rlabel via3 14973 42908 14973 42908 0 net169
rlabel metal2 1610 20927 1610 20927 0 net17
rlabel metal2 24426 42925 24426 42925 0 net170
rlabel metal2 14858 41400 14858 41400 0 net171
rlabel metal3 15088 18020 15088 18020 0 net172
rlabel metal2 15640 26894 15640 26894 0 net173
rlabel metal2 20838 42466 20838 42466 0 net174
rlabel metal1 18676 41786 18676 41786 0 net175
rlabel metal1 19596 41786 19596 41786 0 net176
rlabel metal1 20194 40698 20194 40698 0 net177
rlabel metal1 19412 41106 19412 41106 0 net178
rlabel metal1 19688 40494 19688 40494 0 net179
rlabel metal1 1932 20910 1932 20910 0 net18
rlabel metal1 4002 37842 4002 37842 0 net180
rlabel metal2 16882 42976 16882 42976 0 net181
rlabel metal1 15548 15130 15548 15130 0 net182
rlabel metal1 17158 42636 17158 42636 0 net183
rlabel metal1 17434 42704 17434 42704 0 net184
rlabel metal1 17756 42670 17756 42670 0 net185
rlabel metal1 18032 42670 18032 42670 0 net186
rlabel metal1 18354 42670 18354 42670 0 net187
rlabel metal1 21114 42772 21114 42772 0 net188
rlabel metal1 23920 8942 23920 8942 0 net189
rlabel metal1 1978 29478 1978 29478 0 net19
rlabel metal1 24104 7446 24104 7446 0 net190
rlabel metal1 22770 8874 22770 8874 0 net191
rlabel metal1 24150 11662 24150 11662 0 net192
rlabel metal2 22494 15300 22494 15300 0 net193
rlabel metal1 23690 16592 23690 16592 0 net194
rlabel metal1 24104 16218 24104 16218 0 net195
rlabel metal1 23138 17170 23138 17170 0 net196
rlabel metal2 20470 13634 20470 13634 0 net197
rlabel metal1 23460 14382 23460 14382 0 net198
rlabel metal1 23782 15096 23782 15096 0 net199
rlabel metal1 1702 35734 1702 35734 0 net2
rlabel metal2 4646 21471 4646 21471 0 net20
rlabel metal2 20838 19584 20838 19584 0 net200
rlabel metal2 21666 13333 21666 13333 0 net201
rlabel metal2 21390 30753 21390 30753 0 net202
rlabel metal1 24564 37706 24564 37706 0 net203
rlabel metal1 23920 12206 23920 12206 0 net204
rlabel metal1 24196 24786 24196 24786 0 net205
rlabel metal1 23230 25194 23230 25194 0 net206
rlabel metal2 18446 33864 18446 33864 0 net207
rlabel metal1 22218 26282 22218 26282 0 net208
rlabel metal1 24150 21624 24150 21624 0 net209
rlabel metal1 1656 28186 1656 28186 0 net21
rlabel metal1 23874 23086 23874 23086 0 net210
rlabel metal1 24150 23800 24150 23800 0 net211
rlabel metal2 21114 24956 21114 24956 0 net212
rlabel metal2 23690 20604 23690 20604 0 net213
rlabel metal1 23552 26758 23552 26758 0 net214
rlabel metal1 21942 31824 21942 31824 0 net215
rlabel metal1 23828 22066 23828 22066 0 net216
rlabel metal2 21344 21012 21344 21012 0 net217
rlabel metal2 23414 20298 23414 20298 0 net218
rlabel metal1 23782 19414 23782 19414 0 net219
rlabel metal1 6532 31382 6532 31382 0 net22
rlabel metal1 21574 24616 21574 24616 0 net220
rlabel metal1 24242 26996 24242 26996 0 net221
rlabel metal1 24242 32334 24242 32334 0 net222
rlabel metal1 23828 32538 23828 32538 0 net223
rlabel metal1 23920 33558 23920 33558 0 net224
rlabel metal1 23966 34000 23966 34000 0 net225
rlabel metal1 24150 34680 24150 34680 0 net226
rlabel metal1 23966 35020 23966 35020 0 net227
rlabel metal1 24150 35632 24150 35632 0 net228
rlabel metal1 23874 36176 23874 36176 0 net229
rlabel metal1 7406 31348 7406 31348 0 net23
rlabel metal2 22402 36516 22402 36516 0 net230
rlabel metal1 20654 36584 20654 36584 0 net231
rlabel metal1 23460 27098 23460 27098 0 net232
rlabel metal2 21666 37536 21666 37536 0 net233
rlabel metal2 23966 38794 23966 38794 0 net234
rlabel metal1 23782 38998 23782 38998 0 net235
rlabel metal2 23966 39610 23966 39610 0 net236
rlabel metal2 21482 39168 21482 39168 0 net237
rlabel metal2 19826 40256 19826 40256 0 net238
rlabel metal3 20332 39984 20332 39984 0 net239
rlabel metal1 2668 39338 2668 39338 0 net24
rlabel metal1 23782 40698 23782 40698 0 net240
rlabel metal2 23506 42636 23506 42636 0 net241
rlabel metal1 22218 42126 22218 42126 0 net242
rlabel metal1 24150 27982 24150 27982 0 net243
rlabel metal1 23368 39882 23368 39882 0 net244
rlabel metal1 22632 39814 22632 39814 0 net245
rlabel metal1 23966 28560 23966 28560 0 net246
rlabel metal1 24150 29104 24150 29104 0 net247
rlabel metal1 23966 29580 23966 29580 0 net248
rlabel metal1 24150 30328 24150 30328 0 net249
rlabel metal2 1610 28237 1610 28237 0 net25
rlabel metal1 23368 30634 23368 30634 0 net250
rlabel metal1 24242 31280 24242 31280 0 net251
rlabel metal1 21873 31926 21873 31926 0 net252
rlabel metal1 20102 41990 20102 41990 0 net253
rlabel metal2 22126 42092 22126 42092 0 net254
rlabel metal2 22126 40936 22126 40936 0 net255
rlabel metal1 23874 41446 23874 41446 0 net256
rlabel metal1 21390 40358 21390 40358 0 net257
rlabel metal1 21758 39814 21758 39814 0 net258
rlabel metal1 24012 42262 24012 42262 0 net259
rlabel via2 1794 21947 1794 21947 0 net26
rlabel metal1 22126 42568 22126 42568 0 net260
rlabel metal1 22218 39814 22218 39814 0 net261
rlabel metal1 23322 41650 23322 41650 0 net262
rlabel metal1 23276 42058 23276 42058 0 net263
rlabel metal1 20516 42058 20516 42058 0 net264
rlabel metal1 20194 40970 20194 40970 0 net265
rlabel metal1 21758 42330 21758 42330 0 net266
rlabel metal1 22724 42806 22724 42806 0 net267
rlabel metal1 22402 40970 22402 40970 0 net268
rlabel metal2 20838 40834 20838 40834 0 net269
rlabel via1 13858 26962 13858 26962 0 net27
rlabel metal1 22448 42602 22448 42602 0 net270
rlabel metal2 21390 42432 21390 42432 0 net271
rlabel metal1 21390 41242 21390 41242 0 net272
rlabel metal2 9154 42585 9154 42585 0 net273
rlabel metal1 3266 40698 3266 40698 0 net274
rlabel metal1 10258 42126 10258 42126 0 net275
rlabel metal2 15502 42432 15502 42432 0 net276
rlabel metal1 2346 41480 2346 41480 0 net277
rlabel metal1 1886 41514 1886 41514 0 net278
rlabel metal1 2162 42330 2162 42330 0 net279
rlabel metal1 2898 24820 2898 24820 0 net28
rlabel metal1 8464 41786 8464 41786 0 net280
rlabel metal1 3036 41242 3036 41242 0 net281
rlabel metal2 2806 41463 2806 41463 0 net282
rlabel metal2 2530 42262 2530 42262 0 net283
rlabel metal1 3358 42330 3358 42330 0 net284
rlabel metal1 2852 41786 2852 41786 0 net285
rlabel metal1 3542 41786 3542 41786 0 net286
rlabel metal2 4462 42194 4462 42194 0 net287
rlabel metal1 3266 41786 3266 41786 0 net288
rlabel metal1 4048 41786 4048 41786 0 net289
rlabel metal1 4416 29682 4416 29682 0 net29
rlabel metal1 4922 42670 4922 42670 0 net290
rlabel metal1 4830 42262 4830 42262 0 net291
rlabel metal1 5014 41786 5014 41786 0 net292
rlabel metal1 5520 41786 5520 41786 0 net293
rlabel metal1 8786 42330 8786 42330 0 net294
rlabel metal2 9982 42500 9982 42500 0 net295
rlabel metal2 10626 42976 10626 42976 0 net296
rlabel metal1 9246 42602 9246 42602 0 net297
rlabel metal1 10028 42874 10028 42874 0 net298
rlabel metal1 16100 42534 16100 42534 0 net299
rlabel metal1 1886 16422 1886 16422 0 net3
rlabel via1 17779 22610 17779 22610 0 net30
rlabel metal1 6118 41786 6118 41786 0 net300
rlabel metal1 5658 41446 5658 41446 0 net301
rlabel metal1 5888 41786 5888 41786 0 net302
rlabel metal1 6762 43384 6762 43384 0 net303
rlabel metal1 7268 41786 7268 41786 0 net304
rlabel metal2 7590 42228 7590 42228 0 net305
rlabel metal1 7866 41480 7866 41480 0 net306
rlabel metal2 8142 42500 8142 42500 0 net307
rlabel metal1 7820 41242 7820 41242 0 net308
rlabel metal1 9338 1224 9338 1224 0 net309
rlabel metal2 1886 26996 1886 26996 0 net31
rlabel metal1 9936 2006 9936 2006 0 net310
rlabel metal2 12558 1632 12558 1632 0 net311
rlabel metal1 15226 2312 15226 2312 0 net312
rlabel metal1 13478 1326 13478 1326 0 net313
rlabel metal1 14076 1258 14076 1258 0 net314
rlabel metal1 14352 1326 14352 1326 0 net315
rlabel metal1 14490 1972 14490 1972 0 net316
rlabel metal1 15042 1938 15042 1938 0 net317
rlabel metal1 15042 1326 15042 1326 0 net318
rlabel metal1 15180 1258 15180 1258 0 net319
rlabel metal1 5750 32776 5750 32776 0 net32
rlabel metal1 16146 1972 16146 1972 0 net320
rlabel metal1 13018 1326 13018 1326 0 net321
rlabel metal1 10304 1326 10304 1326 0 net322
rlabel metal1 12006 2040 12006 2040 0 net323
rlabel metal1 11316 1326 11316 1326 0 net324
rlabel metal1 12236 1326 12236 1326 0 net325
rlabel metal1 12650 2006 12650 2006 0 net326
rlabel metal2 11822 1530 11822 1530 0 net327
rlabel metal1 12696 1326 12696 1326 0 net328
rlabel metal2 16330 1700 16330 1700 0 net329
rlabel metal2 12650 25670 12650 25670 0 net33
rlabel metal1 18676 2414 18676 2414 0 net330
rlabel metal2 18768 3026 18768 3026 0 net331
rlabel metal1 17848 2550 17848 2550 0 net332
rlabel metal1 18998 4182 18998 4182 0 net333
rlabel metal1 20792 3502 20792 3502 0 net334
rlabel metal1 21666 3026 21666 3026 0 net335
rlabel metal2 16238 1768 16238 1768 0 net336
rlabel metal1 16974 1326 16974 1326 0 net337
rlabel metal1 17710 1326 17710 1326 0 net338
rlabel metal2 16790 2550 16790 2550 0 net339
rlabel metal1 9246 35054 9246 35054 0 net34
rlabel metal1 18170 2074 18170 2074 0 net340
rlabel metal1 17802 1938 17802 1938 0 net341
rlabel metal1 17848 2006 17848 2006 0 net342
rlabel metal1 18400 1326 18400 1326 0 net343
rlabel metal1 18308 2414 18308 2414 0 net344
rlabel metal1 20562 41614 20562 41614 0 net345
rlabel metal1 2438 3162 2438 3162 0 net346
rlabel metal1 3496 5610 3496 5610 0 net347
rlabel metal1 1702 3536 1702 3536 0 net348
rlabel metal2 3818 5508 3818 5508 0 net349
rlabel metal1 15548 30702 15548 30702 0 net35
rlabel metal1 2714 2924 2714 2924 0 net350
rlabel metal1 4002 6358 4002 6358 0 net351
rlabel metal1 3542 5678 3542 5678 0 net352
rlabel metal1 2254 6256 2254 6256 0 net353
rlabel metal2 2162 3808 2162 3808 0 net354
rlabel metal1 1702 5712 1702 5712 0 net355
rlabel metal1 1518 4216 1518 4216 0 net356
rlabel metal2 3174 5644 3174 5644 0 net357
rlabel metal2 2162 6086 2162 6086 0 net358
rlabel metal1 2392 7514 2392 7514 0 net359
rlabel metal1 12834 27030 12834 27030 0 net36
rlabel metal2 2254 7854 2254 7854 0 net360
rlabel metal1 2691 8534 2691 8534 0 net361
rlabel metal1 3772 6630 3772 6630 0 net362
rlabel metal1 3174 9044 3174 9044 0 net363
rlabel metal2 1518 6086 1518 6086 0 net364
rlabel metal1 2852 3638 2852 3638 0 net365
rlabel metal1 1518 12920 1518 12920 0 net366
rlabel metal2 2070 17816 2070 17816 0 net367
rlabel metal1 10534 14552 10534 14552 0 net368
rlabel metal1 2070 15402 2070 15402 0 net369
rlabel metal2 1978 26656 1978 26656 0 net37
rlabel via2 1794 36635 1794 36635 0 net370
rlabel metal1 3312 15062 3312 15062 0 net371
rlabel metal1 3358 13328 3358 13328 0 net372
rlabel metal1 1886 15130 1886 15130 0 net373
rlabel metal1 2438 16592 2438 16592 0 net374
rlabel metal1 3082 15402 3082 15402 0 net375
rlabel metal1 14582 16456 14582 16456 0 net376
rlabel metal1 3864 16490 3864 16490 0 net377
rlabel metal2 2070 8262 2070 8262 0 net378
rlabel metal1 1932 13226 1932 13226 0 net379
rlabel metal1 3266 28186 3266 28186 0 net38
rlabel metal1 3910 12240 3910 12240 0 net380
rlabel metal1 3956 9146 3956 9146 0 net381
rlabel metal1 2116 10982 2116 10982 0 net382
rlabel metal1 2622 7752 2622 7752 0 net383
rlabel metal1 10994 10744 10994 10744 0 net384
rlabel metal2 1978 12410 1978 12410 0 net385
rlabel metal1 1886 8942 1886 8942 0 net386
rlabel metal1 2093 9350 2093 9350 0 net387
rlabel metal2 2530 8670 2530 8670 0 net388
rlabel metal1 5244 11118 5244 11118 0 net389
rlabel metal1 16284 26894 16284 26894 0 net39
rlabel metal1 1748 8534 1748 8534 0 net390
rlabel metal1 4416 12206 4416 12206 0 net391
rlabel metal2 2622 10268 2622 10268 0 net392
rlabel metal2 2254 10914 2254 10914 0 net393
rlabel metal1 14536 16558 14536 16558 0 net394
rlabel metal1 16468 19278 16468 19278 0 net395
rlabel metal1 7406 19380 7406 19380 0 net396
rlabel metal1 5382 19754 5382 19754 0 net397
rlabel metal1 15594 20978 15594 20978 0 net398
rlabel metal1 16100 23698 16100 23698 0 net399
rlabel metal1 17434 18258 17434 18258 0 net4
rlabel metal2 5014 33660 5014 33660 0 net40
rlabel metal1 6762 21590 6762 21590 0 net400
rlabel metal1 6854 25908 6854 25908 0 net401
rlabel metal1 14950 22066 14950 22066 0 net402
rlabel metal1 13662 17714 13662 17714 0 net403
rlabel metal1 4186 33082 4186 33082 0 net404
rlabel metal2 12742 40256 12742 40256 0 net405
rlabel metal1 11684 18258 11684 18258 0 net406
rlabel metal1 3450 39508 3450 39508 0 net407
rlabel metal1 11086 40052 11086 40052 0 net408
rlabel metal1 18400 17782 18400 17782 0 net409
rlabel metal1 1932 25466 1932 25466 0 net41
rlabel metal1 16192 28526 16192 28526 0 net42
rlabel metal1 6852 24072 6852 24072 0 net43
rlabel metal1 3864 24922 3864 24922 0 net44
rlabel metal1 11270 33490 11270 33490 0 net45
rlabel metal1 14858 25330 14858 25330 0 net46
rlabel metal1 11592 26282 11592 26282 0 net47
rlabel metal2 3542 27302 3542 27302 0 net48
rlabel metal2 20838 14518 20838 14518 0 net49
rlabel metal1 15686 19788 15686 19788 0 net5
rlabel metal1 1885 34578 1885 34578 0 net50
rlabel metal1 19642 32198 19642 32198 0 net51
rlabel via1 2621 19822 2621 19822 0 net52
rlabel metal1 2115 18734 2115 18734 0 net53
rlabel metal1 16882 20842 16882 20842 0 net54
rlabel metal1 14903 34578 14903 34578 0 net55
rlabel metal1 1702 40120 1702 40120 0 net56
rlabel metal1 14719 35666 14719 35666 0 net57
rlabel metal1 20101 33966 20101 33966 0 net58
rlabel metal2 2024 32028 2024 32028 0 net59
rlabel metal1 3910 22202 3910 22202 0 net6
rlabel via2 1702 32827 1702 32827 0 net60
rlabel metal1 2024 1938 2024 1938 0 net61
rlabel metal1 2575 2414 2575 2414 0 net62
rlabel via1 14657 20434 14657 20434 0 net63
rlabel viali 14205 12848 14205 12848 0 net64
rlabel metal2 1702 21641 1702 21641 0 net65
rlabel via2 14950 13923 14950 13923 0 net66
rlabel metal1 19182 40086 19182 40086 0 net67
rlabel viali 2254 40023 2254 40023 0 net68
rlabel metal2 1012 16660 1012 16660 0 net69
rlabel metal1 2806 21658 2806 21658 0 net7
rlabel metal2 20194 15674 20194 15674 0 net70
rlabel metal2 17986 11475 17986 11475 0 net71
rlabel metal1 19550 20944 19550 20944 0 net72
rlabel metal2 19642 19958 19642 19958 0 net73
rlabel metal1 22080 28492 22080 28492 0 net74
rlabel metal2 12558 40834 12558 40834 0 net75
rlabel metal1 14811 28526 14811 28526 0 net76
rlabel metal2 15272 21692 15272 21692 0 net77
rlabel metal4 2484 34748 2484 34748 0 net78
rlabel metal1 8832 2482 8832 2482 0 net79
rlabel metal1 3726 21862 3726 21862 0 net8
rlabel metal2 20654 32411 20654 32411 0 net80
rlabel metal1 19964 1870 19964 1870 0 net81
rlabel metal2 21528 8364 21528 8364 0 net82
rlabel metal1 20102 1190 20102 1190 0 net83
rlabel metal2 25162 17204 25162 17204 0 net84
rlabel metal1 21436 5882 21436 5882 0 net85
rlabel metal2 20424 13396 20424 13396 0 net86
rlabel metal2 20102 7378 20102 7378 0 net87
rlabel metal3 22839 35972 22839 35972 0 net88
rlabel metal3 19895 2652 19895 2652 0 net89
rlabel metal1 1702 23562 1702 23562 0 net9
rlabel metal1 19826 1530 19826 1530 0 net90
rlabel metal2 21298 1020 21298 1020 0 net91
rlabel metal2 16330 40868 16330 40868 0 net92
rlabel metal1 21436 2006 21436 2006 0 net93
rlabel metal1 2208 29070 2208 29070 0 net94
rlabel metal1 20746 2380 20746 2380 0 net95
rlabel metal1 1518 18802 1518 18802 0 net96
rlabel metal1 14122 18258 14122 18258 0 net97
rlabel metal3 13547 17884 13547 17884 0 net98
rlabel metal1 19826 16660 19826 16660 0 net99
rlabel metal1 20194 42228 20194 42228 0 strobe_inbuf_0.X
rlabel metal1 20194 41242 20194 41242 0 strobe_inbuf_1.X
rlabel metal2 22218 13311 22218 13311 0 strobe_inbuf_10.X
rlabel metal1 24012 40630 24012 40630 0 strobe_inbuf_11.X
rlabel metal1 23552 35802 23552 35802 0 strobe_inbuf_12.X
rlabel metal2 23414 25092 23414 25092 0 strobe_inbuf_13.X
rlabel metal1 23920 21862 23920 21862 0 strobe_inbuf_14.X
rlabel metal1 23644 32878 23644 32878 0 strobe_inbuf_15.X
rlabel metal1 22632 37434 22632 37434 0 strobe_inbuf_16.X
rlabel metal1 22908 34170 22908 34170 0 strobe_inbuf_17.X
rlabel metal1 24012 36890 24012 36890 0 strobe_inbuf_18.X
rlabel metal1 23828 31994 23828 31994 0 strobe_inbuf_19.X
rlabel metal1 20562 36890 20562 36890 0 strobe_inbuf_2.X
rlabel metal1 20838 39066 20838 39066 0 strobe_inbuf_3.X
rlabel metal1 21850 41582 21850 41582 0 strobe_inbuf_4.X
rlabel metal1 21804 21658 21804 21658 0 strobe_inbuf_5.X
rlabel metal1 21620 39406 21620 39406 0 strobe_inbuf_6.X
rlabel metal1 20838 37978 20838 37978 0 strobe_inbuf_7.X
rlabel metal2 22402 40052 22402 40052 0 strobe_inbuf_8.X
rlabel metal2 20654 40681 20654 40681 0 strobe_inbuf_9.X
rlabel metal1 20470 42262 20470 42262 0 strobe_outbuf_0.X
rlabel metal2 20286 41956 20286 41956 0 strobe_outbuf_1.X
rlabel metal1 21758 39984 21758 39984 0 strobe_outbuf_10.X
rlabel metal1 21896 40494 21896 40494 0 strobe_outbuf_11.X
rlabel metal1 23506 36346 23506 36346 0 strobe_outbuf_12.X
rlabel metal1 24150 26010 24150 26010 0 strobe_outbuf_13.X
rlabel metal1 21804 40086 21804 40086 0 strobe_outbuf_14.X
rlabel metal1 23598 32742 23598 32742 0 strobe_outbuf_15.X
rlabel metal2 21114 39083 21114 39083 0 strobe_outbuf_16.X
rlabel metal1 22862 35258 22862 35258 0 strobe_outbuf_17.X
rlabel metal2 20746 38964 20746 38964 0 strobe_outbuf_18.X
rlabel metal1 24012 32198 24012 32198 0 strobe_outbuf_19.X
rlabel metal2 20562 39100 20562 39100 0 strobe_outbuf_2.X
rlabel metal1 20838 39610 20838 39610 0 strobe_outbuf_3.X
rlabel metal1 22080 41446 22080 41446 0 strobe_outbuf_4.X
rlabel metal2 22218 40358 22218 40358 0 strobe_outbuf_5.X
rlabel metal1 21298 39610 21298 39610 0 strobe_outbuf_6.X
rlabel metal1 18216 40630 18216 40630 0 strobe_outbuf_7.X
rlabel metal1 22402 40698 22402 40698 0 strobe_outbuf_8.X
rlabel metal2 22770 40868 22770 40868 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 44623
<< end >>
