magic
tech sky130A
magscale 1 2
timestamp 1732489752
<< viali >>
rect 2329 6409 2363 6443
rect 3433 6409 3467 6443
rect 4353 6409 4387 6443
rect 4905 6409 4939 6443
rect 5457 6409 5491 6443
rect 6469 6409 6503 6443
rect 7113 6409 7147 6443
rect 7573 6409 7607 6443
rect 8033 6409 8067 6443
rect 8585 6409 8619 6443
rect 9413 6409 9447 6443
rect 9873 6409 9907 6443
rect 10517 6409 10551 6443
rect 10885 6409 10919 6443
rect 11529 6409 11563 6443
rect 12633 6409 12667 6443
rect 14657 6409 14691 6443
rect 14933 6409 14967 6443
rect 16957 6409 16991 6443
rect 17233 6409 17267 6443
rect 19257 6409 19291 6443
rect 20361 6409 20395 6443
rect 20913 6409 20947 6443
rect 22201 6409 22235 6443
rect 22569 6409 22603 6443
rect 23673 6409 23707 6443
rect 1501 6341 1535 6375
rect 2421 6341 2455 6375
rect 5549 6341 5583 6375
rect 7205 6341 7239 6375
rect 8125 6341 8159 6375
rect 8677 6341 8711 6375
rect 1869 6273 1903 6307
rect 2973 6273 3007 6307
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 4445 6273 4479 6307
rect 4997 6273 5031 6307
rect 6101 6273 6135 6307
rect 6665 6273 6699 6307
rect 7389 6273 7423 6307
rect 9321 6273 9355 6307
rect 10149 6273 10183 6307
rect 10425 6273 10459 6307
rect 11069 6273 11103 6307
rect 11345 6273 11379 6307
rect 11713 6273 11747 6307
rect 11805 6273 11839 6307
rect 12265 6273 12299 6307
rect 12357 6273 12391 6307
rect 12825 6277 12859 6311
rect 13093 6273 13127 6307
rect 13369 6273 13403 6307
rect 13645 6273 13679 6307
rect 13921 6273 13955 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 14841 6273 14875 6307
rect 15117 6273 15151 6307
rect 15393 6273 15427 6307
rect 15669 6273 15703 6307
rect 15945 6273 15979 6307
rect 16221 6273 16255 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 17141 6273 17175 6307
rect 17417 6273 17451 6307
rect 17693 6273 17727 6307
rect 17969 6273 18003 6307
rect 18245 6273 18279 6307
rect 18521 6273 18555 6307
rect 18797 6273 18831 6307
rect 19073 6273 19107 6307
rect 19441 6273 19475 6307
rect 19717 6273 19751 6307
rect 19993 6273 20027 6307
rect 20269 6273 20303 6307
rect 20821 6273 20855 6307
rect 21465 6273 21499 6307
rect 21925 6273 21959 6307
rect 22477 6273 22511 6307
rect 23029 6273 23063 6307
rect 23581 6273 23615 6307
rect 2697 6205 2731 6239
rect 11161 6137 11195 6171
rect 13185 6137 13219 6171
rect 13461 6137 13495 6171
rect 14105 6137 14139 6171
rect 15485 6137 15519 6171
rect 16037 6137 16071 6171
rect 16313 6137 16347 6171
rect 16681 6137 16715 6171
rect 17509 6137 17543 6171
rect 18061 6137 18095 6171
rect 18337 6137 18371 6171
rect 19533 6137 19567 6171
rect 3985 6069 4019 6103
rect 6009 6069 6043 6103
rect 11989 6069 12023 6103
rect 12081 6069 12115 6103
rect 12541 6069 12575 6103
rect 12909 6069 12943 6103
rect 13737 6069 13771 6103
rect 14381 6069 14415 6103
rect 15209 6069 15243 6103
rect 15761 6069 15795 6103
rect 17785 6069 17819 6103
rect 18613 6069 18647 6103
rect 18889 6069 18923 6103
rect 19809 6069 19843 6103
rect 21649 6069 21683 6103
rect 23121 6069 23155 6103
rect 1777 5865 1811 5899
rect 2329 5865 2363 5899
rect 2697 5865 2731 5899
rect 3249 5865 3283 5899
rect 4077 5865 4111 5899
rect 4537 5865 4571 5899
rect 4905 5865 4939 5899
rect 6009 5865 6043 5899
rect 6561 5865 6595 5899
rect 7941 5865 7975 5899
rect 8401 5865 8435 5899
rect 9137 5865 9171 5899
rect 9413 5865 9447 5899
rect 12633 5865 12667 5899
rect 14657 5865 14691 5899
rect 15393 5865 15427 5899
rect 15669 5865 15703 5899
rect 16497 5865 16531 5899
rect 16957 5865 16991 5899
rect 17601 5865 17635 5899
rect 18429 5865 18463 5899
rect 19257 5865 19291 5899
rect 19533 5865 19567 5899
rect 21465 5865 21499 5899
rect 22569 5865 22603 5899
rect 23121 5865 23155 5899
rect 23673 5865 23707 5899
rect 5825 5797 5859 5831
rect 7205 5797 7239 5831
rect 9965 5797 9999 5831
rect 10241 5797 10275 5831
rect 11345 5797 11379 5831
rect 12173 5797 12207 5831
rect 15945 5797 15979 5831
rect 16221 5797 16255 5831
rect 17325 5797 17359 5831
rect 18705 5797 18739 5831
rect 19809 5797 19843 5831
rect 20545 5797 20579 5831
rect 21189 5797 21223 5831
rect 22201 5797 22235 5831
rect 1869 5661 1903 5695
rect 2973 5661 3007 5695
rect 3525 5661 3559 5695
rect 4721 5661 4755 5695
rect 5549 5661 5583 5695
rect 5641 5661 5675 5695
rect 9321 5661 9355 5695
rect 9597 5661 9631 5695
rect 9689 5661 9723 5695
rect 10149 5661 10183 5695
rect 10425 5661 10459 5695
rect 10701 5661 10735 5695
rect 10977 5661 11011 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 11805 5661 11839 5695
rect 12081 5661 12115 5695
rect 12357 5661 12391 5695
rect 12817 5661 12851 5695
rect 13185 5661 13219 5695
rect 13461 5661 13495 5695
rect 14565 5661 14599 5695
rect 14841 5661 14875 5695
rect 15577 5661 15611 5695
rect 15853 5661 15887 5695
rect 16129 5661 16163 5695
rect 16405 5661 16439 5695
rect 16681 5661 16715 5695
rect 16773 5661 16807 5695
rect 17233 5661 17267 5695
rect 17509 5661 17543 5695
rect 17785 5661 17819 5695
rect 18061 5661 18095 5695
rect 18337 5661 18371 5695
rect 18613 5661 18647 5695
rect 18889 5661 18923 5695
rect 19441 5661 19475 5695
rect 19717 5661 19751 5695
rect 19993 5661 20027 5695
rect 20269 5661 20303 5695
rect 20361 5661 20395 5695
rect 20821 5661 20855 5695
rect 21649 5661 21683 5695
rect 24225 5661 24259 5695
rect 2421 5593 2455 5627
rect 4353 5593 4387 5627
rect 5181 5593 5215 5627
rect 6285 5593 6319 5627
rect 6837 5593 6871 5627
rect 7389 5593 7423 5627
rect 7849 5593 7883 5627
rect 8677 5593 8711 5627
rect 21005 5593 21039 5627
rect 21925 5593 21959 5627
rect 22477 5593 22511 5627
rect 23029 5593 23063 5627
rect 23581 5593 23615 5627
rect 5365 5525 5399 5559
rect 9873 5525 9907 5559
rect 10517 5525 10551 5559
rect 10793 5525 10827 5559
rect 11069 5525 11103 5559
rect 11621 5525 11655 5559
rect 11897 5525 11931 5559
rect 13001 5525 13035 5559
rect 13277 5525 13311 5559
rect 14381 5525 14415 5559
rect 17049 5525 17083 5559
rect 17877 5525 17911 5559
rect 18153 5525 18187 5559
rect 20085 5525 20119 5559
rect 20637 5525 20671 5559
rect 24041 5525 24075 5559
rect 1869 5321 1903 5355
rect 3433 5321 3467 5355
rect 3709 5321 3743 5355
rect 4537 5321 4571 5355
rect 4905 5321 4939 5355
rect 5181 5321 5215 5355
rect 5549 5321 5583 5355
rect 5825 5321 5859 5355
rect 6377 5321 6411 5355
rect 6929 5321 6963 5355
rect 7297 5321 7331 5355
rect 7573 5321 7607 5355
rect 7849 5321 7883 5355
rect 8677 5321 8711 5355
rect 9137 5321 9171 5355
rect 10149 5321 10183 5355
rect 10241 5321 10275 5355
rect 18705 5321 18739 5355
rect 18981 5321 19015 5355
rect 19533 5321 19567 5355
rect 20913 5321 20947 5355
rect 21649 5321 21683 5355
rect 23857 5321 23891 5355
rect 2145 5253 2179 5287
rect 3065 5253 3099 5287
rect 4629 5253 4663 5287
rect 22109 5253 22143 5287
rect 23489 5253 23523 5287
rect 1961 5185 1995 5219
rect 2513 5185 2547 5219
rect 3617 5185 3651 5219
rect 3893 5185 3927 5219
rect 4169 5185 4203 5219
rect 5089 5185 5123 5219
rect 5365 5185 5399 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7113 5185 7147 5219
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 8033 5185 8067 5219
rect 8309 5185 8343 5219
rect 8585 5185 8619 5219
rect 8861 5185 8895 5219
rect 9321 5185 9355 5219
rect 9689 5185 9723 5219
rect 9965 5185 9999 5219
rect 10425 5185 10459 5219
rect 10977 5185 11011 5219
rect 11253 5185 11287 5219
rect 11713 5185 11747 5219
rect 18521 5185 18555 5219
rect 18797 5185 18831 5219
rect 19073 5185 19107 5219
rect 19349 5185 19383 5219
rect 19809 5185 19843 5219
rect 20269 5185 20303 5219
rect 20453 5185 20487 5219
rect 20729 5185 20763 5219
rect 21373 5185 21407 5219
rect 21465 5185 21499 5219
rect 22937 5185 22971 5219
rect 23765 5185 23799 5219
rect 2789 5117 2823 5151
rect 22385 5117 22419 5151
rect 22661 5117 22695 5151
rect 8401 5049 8435 5083
rect 9873 5049 9907 5083
rect 11529 5049 11563 5083
rect 19257 5049 19291 5083
rect 19993 5049 20027 5083
rect 20085 5049 20119 5083
rect 3985 4981 4019 5015
rect 6653 4981 6687 5015
rect 8125 4981 8159 5015
rect 10793 4981 10827 5015
rect 11069 4981 11103 5015
rect 20637 4981 20671 5015
rect 21189 4981 21223 5015
rect 23397 4981 23431 5015
rect 1501 4777 1535 4811
rect 2145 4777 2179 4811
rect 2605 4777 2639 4811
rect 3065 4777 3099 4811
rect 4629 4777 4663 4811
rect 19441 4777 19475 4811
rect 21741 4777 21775 4811
rect 22569 4777 22603 4811
rect 23121 4777 23155 4811
rect 23949 4777 23983 4811
rect 3157 4709 3191 4743
rect 2789 4573 2823 4607
rect 2881 4573 2915 4607
rect 3341 4573 3375 4607
rect 4813 4573 4847 4607
rect 16865 4573 16899 4607
rect 19257 4573 19291 4607
rect 21557 4573 21591 4607
rect 21833 4573 21867 4607
rect 22109 4573 22143 4607
rect 23489 4573 23523 4607
rect 1777 4505 1811 4539
rect 2053 4505 2087 4539
rect 22477 4505 22511 4539
rect 23029 4505 23063 4539
rect 23857 4505 23891 4539
rect 17049 4437 17083 4471
rect 22017 4437 22051 4471
rect 22293 4437 22327 4471
rect 23673 4437 23707 4471
rect 19441 4233 19475 4267
rect 22109 4233 22143 4267
rect 23121 4165 23155 4199
rect 1501 4097 1535 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 19257 4097 19291 4131
rect 20085 4097 20119 4131
rect 22293 4097 22327 4131
rect 22385 4097 22419 4131
rect 22661 4097 22695 4131
rect 23673 4097 23707 4131
rect 24317 4097 24351 4131
rect 23397 4029 23431 4063
rect 23949 4029 23983 4063
rect 2421 3961 2455 3995
rect 20269 3961 20303 3995
rect 1593 3893 1627 3927
rect 2145 3893 2179 3927
rect 22569 3893 22603 3927
rect 22845 3893 22879 3927
rect 24133 3893 24167 3927
rect 1501 3689 1535 3723
rect 1961 3689 1995 3723
rect 18797 3689 18831 3723
rect 19625 3689 19659 3723
rect 23305 3689 23339 3723
rect 24133 3689 24167 3723
rect 22937 3621 22971 3655
rect 1685 3485 1719 3519
rect 1777 3485 1811 3519
rect 18613 3485 18647 3519
rect 19441 3485 19475 3519
rect 22753 3485 22787 3519
rect 23121 3485 23155 3519
rect 23673 3485 23707 3519
rect 23857 3417 23891 3451
rect 23489 3349 23523 3383
rect 18245 3145 18279 3179
rect 19073 3145 19107 3179
rect 18061 3009 18095 3043
rect 18889 3009 18923 3043
rect 24041 3009 24075 3043
rect 24317 3009 24351 3043
rect 24133 2873 24167 2907
rect 23857 2805 23891 2839
rect 11989 2601 12023 2635
rect 13461 2601 13495 2635
rect 19993 2601 20027 2635
rect 24041 2601 24075 2635
rect 8585 2533 8619 2567
rect 15669 2533 15703 2567
rect 7113 2397 7147 2431
rect 8401 2397 8435 2431
rect 9597 2397 9631 2431
rect 10793 2397 10827 2431
rect 11805 2397 11839 2431
rect 12173 2397 12207 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 15485 2397 15519 2431
rect 19809 2397 19843 2431
rect 24225 2397 24259 2431
rect 7297 2261 7331 2295
rect 9781 2261 9815 2295
rect 10977 2261 11011 2295
rect 12357 2261 12391 2295
rect 14565 2261 14599 2295
rect 6745 2057 6779 2091
rect 8033 2057 8067 2091
rect 9229 2057 9263 2091
rect 10425 2057 10459 2091
rect 11713 2057 11747 2091
rect 11989 2057 12023 2091
rect 12817 2057 12851 2091
rect 14013 2057 14047 2091
rect 15117 2057 15151 2091
rect 18797 2057 18831 2091
rect 19441 2057 19475 2091
rect 24317 2057 24351 2091
rect 6561 1921 6595 1955
rect 7849 1921 7883 1955
rect 9045 1921 9079 1955
rect 10241 1921 10275 1955
rect 11529 1921 11563 1955
rect 11805 1921 11839 1955
rect 12633 1921 12667 1955
rect 13829 1921 13863 1955
rect 14933 1921 14967 1955
rect 18613 1921 18647 1955
rect 19257 1921 19291 1955
rect 24133 1921 24167 1955
rect 2421 1513 2455 1547
rect 6561 1513 6595 1547
rect 7481 1513 7515 1547
rect 8677 1513 8711 1547
rect 9873 1513 9907 1547
rect 11161 1513 11195 1547
rect 12265 1513 12299 1547
rect 14657 1513 14691 1547
rect 23489 1513 23523 1547
rect 6009 1445 6043 1479
rect 7205 1445 7239 1479
rect 1409 1309 1443 1343
rect 2237 1309 2271 1343
rect 3433 1309 3467 1343
rect 4629 1309 4663 1343
rect 5825 1309 5859 1343
rect 6377 1309 6411 1343
rect 7021 1309 7055 1343
rect 7297 1309 7331 1343
rect 8217 1309 8251 1343
rect 8493 1309 8527 1343
rect 9413 1309 9447 1343
rect 9689 1309 9723 1343
rect 10425 1309 10459 1343
rect 10701 1309 10735 1343
rect 10977 1309 11011 1343
rect 11805 1309 11839 1343
rect 12081 1309 12115 1343
rect 13001 1309 13035 1343
rect 13277 1309 13311 1343
rect 14197 1309 14231 1343
rect 14473 1309 14507 1343
rect 15393 1309 15427 1343
rect 16681 1309 16715 1343
rect 17785 1309 17819 1343
rect 18705 1309 18739 1343
rect 19257 1309 19291 1343
rect 20177 1309 20211 1343
rect 21373 1309 21407 1343
rect 22569 1309 22603 1343
rect 23305 1309 23339 1343
rect 23949 1309 23983 1343
rect 24041 1309 24075 1343
rect 1593 1173 1627 1207
rect 3617 1173 3651 1207
rect 4813 1173 4847 1207
rect 8401 1173 8435 1207
rect 9597 1173 9631 1207
rect 10609 1173 10643 1207
rect 10885 1173 10919 1207
rect 11989 1173 12023 1207
rect 13185 1173 13219 1207
rect 13461 1173 13495 1207
rect 14381 1173 14415 1207
rect 15577 1173 15611 1207
rect 16865 1173 16899 1207
rect 17969 1173 18003 1207
rect 18889 1173 18923 1207
rect 19441 1173 19475 1207
rect 20361 1173 20395 1207
rect 21557 1173 21591 1207
rect 22753 1173 22787 1207
rect 23765 1173 23799 1207
rect 24225 1173 24259 1207
<< metal1 >>
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 19426 7936 19432 7948
rect 9180 7908 19432 7936
rect 9180 7896 9186 7908
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 8018 7828 8024 7880
rect 8076 7868 8082 7880
rect 19334 7868 19340 7880
rect 8076 7840 19340 7868
rect 8076 7828 8082 7840
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 7742 7760 7748 7812
rect 7800 7800 7806 7812
rect 17954 7800 17960 7812
rect 7800 7772 17960 7800
rect 7800 7760 7806 7772
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 21910 7760 21916 7812
rect 21968 7800 21974 7812
rect 23474 7800 23480 7812
rect 21968 7772 23480 7800
rect 21968 7760 21974 7772
rect 23474 7760 23480 7772
rect 23532 7760 23538 7812
rect 18230 7732 18236 7744
rect 7668 7704 18236 7732
rect 7668 7608 7696 7704
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 8754 7624 8760 7676
rect 8812 7664 8818 7676
rect 17402 7664 17408 7676
rect 8812 7636 17408 7664
rect 8812 7624 8818 7636
rect 17402 7624 17408 7636
rect 17460 7624 17466 7676
rect 7650 7556 7656 7608
rect 7708 7556 7714 7608
rect 8110 7556 8116 7608
rect 8168 7596 8174 7608
rect 11146 7596 11152 7608
rect 8168 7568 11152 7596
rect 8168 7556 8174 7568
rect 11146 7556 11152 7568
rect 11204 7556 11210 7608
rect 10778 7528 10784 7540
rect 4724 7500 10784 7528
rect 4724 7404 4752 7500
rect 10778 7488 10784 7500
rect 10836 7488 10842 7540
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 11054 7460 11060 7472
rect 5960 7432 11060 7460
rect 5960 7420 5966 7432
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 21542 7460 21548 7472
rect 11940 7432 21548 7460
rect 11940 7420 11946 7432
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 8662 7392 8668 7404
rect 5040 7364 8668 7392
rect 5040 7352 5046 7364
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 10870 7324 10876 7336
rect 2924 7296 10876 7324
rect 2924 7284 2930 7296
rect 10870 7284 10876 7296
rect 10928 7284 10934 7336
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12342 7324 12348 7336
rect 11756 7296 12348 7324
rect 11756 7284 11762 7296
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12250 7256 12256 7268
rect 9692 7228 12256 7256
rect 9692 7200 9720 7228
rect 12250 7216 12256 7228
rect 12308 7216 12314 7268
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 8110 7188 8116 7200
rect 4580 7160 8116 7188
rect 4580 7148 4586 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9674 7148 9680 7200
rect 9732 7148 9738 7200
rect 12618 7188 12624 7200
rect 12360 7160 12624 7188
rect 4798 7080 4804 7132
rect 4856 7120 4862 7132
rect 12360 7120 12388 7160
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 17678 7148 17684 7200
rect 17736 7188 17742 7200
rect 18414 7188 18420 7200
rect 17736 7160 18420 7188
rect 17736 7148 17742 7160
rect 18414 7148 18420 7160
rect 18472 7148 18478 7200
rect 17494 7120 17500 7132
rect 4856 7092 12388 7120
rect 12452 7092 17500 7120
rect 4856 7080 4862 7092
rect 8294 7012 8300 7064
rect 8352 7052 8358 7064
rect 12452 7052 12480 7092
rect 17494 7080 17500 7092
rect 17552 7080 17558 7132
rect 20530 7052 20536 7064
rect 8352 7024 12480 7052
rect 19306 7024 20536 7052
rect 8352 7012 8358 7024
rect 8110 6944 8116 6996
rect 8168 6984 8174 6996
rect 12342 6984 12348 6996
rect 8168 6956 12348 6984
rect 8168 6944 8174 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 19306 6984 19334 7024
rect 20530 7012 20536 7024
rect 20588 7012 20594 7064
rect 14148 6956 19334 6984
rect 14148 6944 14154 6956
rect 3418 6876 3424 6928
rect 3476 6916 3482 6928
rect 9674 6916 9680 6928
rect 3476 6888 9680 6916
rect 3476 6876 3482 6888
rect 9674 6876 9680 6888
rect 9732 6876 9738 6928
rect 9766 6876 9772 6928
rect 9824 6916 9830 6928
rect 16942 6916 16948 6928
rect 9824 6888 16948 6916
rect 9824 6876 9830 6888
rect 16942 6876 16948 6888
rect 17000 6876 17006 6928
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 9214 6848 9220 6860
rect 4304 6820 9220 6848
rect 4304 6808 4310 6820
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 14734 6848 14740 6860
rect 9548 6820 14740 6848
rect 9548 6808 9554 6820
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15746 6848 15752 6860
rect 14884 6820 15752 6848
rect 14884 6808 14890 6820
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 15930 6808 15936 6860
rect 15988 6848 15994 6860
rect 16390 6848 16396 6860
rect 15988 6820 16396 6848
rect 15988 6808 15994 6820
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 18046 6848 18052 6860
rect 16816 6820 18052 6848
rect 16816 6808 16822 6820
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 14090 6780 14096 6792
rect 6236 6752 14096 6780
rect 6236 6740 6242 6752
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 19610 6780 19616 6792
rect 14476 6752 19616 6780
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 14476 6644 14504 6752
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 18138 6672 18144 6724
rect 18196 6712 18202 6724
rect 19702 6712 19708 6724
rect 18196 6684 19708 6712
rect 18196 6672 18202 6684
rect 19702 6672 19708 6684
rect 19760 6672 19766 6724
rect 8444 6616 14504 6644
rect 8444 6604 8450 6616
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 18322 6644 18328 6656
rect 17092 6616 18328 6644
rect 17092 6604 17098 6616
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 2317 6443 2375 6449
rect 2317 6409 2329 6443
rect 2363 6440 2375 6443
rect 2958 6440 2964 6452
rect 2363 6412 2964 6440
rect 2363 6409 2375 6412
rect 2317 6403 2375 6409
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 4062 6440 4068 6452
rect 3467 6412 4068 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4246 6400 4252 6452
rect 4304 6400 4310 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 4893 6443 4951 6449
rect 4893 6409 4905 6443
rect 4939 6440 4951 6443
rect 5258 6440 5264 6452
rect 4939 6412 5264 6440
rect 4939 6409 4951 6412
rect 4893 6403 4951 6409
rect 474 6332 480 6384
rect 532 6372 538 6384
rect 1489 6375 1547 6381
rect 1489 6372 1501 6375
rect 532 6344 1501 6372
rect 532 6332 538 6344
rect 1489 6341 1501 6344
rect 1535 6341 1547 6375
rect 1489 6335 1547 6341
rect 2409 6375 2467 6381
rect 2409 6341 2421 6375
rect 2455 6372 2467 6375
rect 2866 6372 2872 6384
rect 2455 6344 2872 6372
rect 2455 6341 2467 6344
rect 2409 6335 2467 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 4264 6372 4292 6400
rect 2976 6344 4292 6372
rect 4356 6372 4384 6403
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5445 6443 5503 6449
rect 5445 6409 5457 6443
rect 5491 6440 5503 6443
rect 5718 6440 5724 6452
rect 5491 6412 5724 6440
rect 5491 6409 5503 6412
rect 5445 6403 5503 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 6178 6440 6184 6452
rect 6012 6412 6184 6440
rect 5166 6372 5172 6384
rect 4356 6344 5172 6372
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6304 1915 6307
rect 2222 6304 2228 6316
rect 1903 6276 2228 6304
rect 1903 6273 1915 6276
rect 1857 6267 1915 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2976 6313 3004 6344
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 5537 6375 5595 6381
rect 5537 6341 5549 6375
rect 5583 6372 5595 6375
rect 6012 6372 6040 6412
rect 6178 6400 6184 6412
rect 6236 6400 6242 6452
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6457 6443 6515 6449
rect 6457 6440 6469 6443
rect 6328 6412 6469 6440
rect 6328 6400 6334 6412
rect 6457 6409 6469 6412
rect 6503 6409 6515 6443
rect 6457 6403 6515 6409
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7374 6440 7380 6452
rect 7147 6412 7380 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7558 6400 7564 6452
rect 7616 6400 7622 6452
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 8478 6440 8484 6452
rect 8067 6412 8484 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 8570 6400 8576 6452
rect 8628 6400 8634 6452
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 9766 6440 9772 6452
rect 9508 6412 9772 6440
rect 7193 6375 7251 6381
rect 5583 6344 6040 6372
rect 6104 6344 7144 6372
rect 5583 6341 5595 6344
rect 5537 6335 5595 6341
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 2685 6239 2743 6245
rect 2685 6205 2697 6239
rect 2731 6236 2743 6239
rect 3326 6236 3332 6248
rect 2731 6208 3332 6236
rect 2731 6205 2743 6208
rect 2685 6199 2743 6205
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 3804 6168 3832 6267
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5810 6304 5816 6316
rect 5031 6276 5816 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6104 6313 6132 6344
rect 7116 6316 7144 6344
rect 7193 6341 7205 6375
rect 7239 6372 7251 6375
rect 7466 6372 7472 6384
rect 7239 6344 7472 6372
rect 7239 6341 7251 6344
rect 7193 6335 7251 6341
rect 7466 6332 7472 6344
rect 7524 6332 7530 6384
rect 8113 6375 8171 6381
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8294 6372 8300 6384
rect 8159 6344 8300 6372
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 8386 6332 8392 6384
rect 8444 6332 8450 6384
rect 8665 6375 8723 6381
rect 8665 6341 8677 6375
rect 8711 6372 8723 6375
rect 9508 6372 9536 6412
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 8711 6344 9536 6372
rect 8711 6341 8723 6344
rect 8665 6335 8723 6341
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 10520 6372 10548 6403
rect 10870 6400 10876 6452
rect 10928 6400 10934 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11112 6412 11529 6440
rect 11112 6400 11118 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11517 6403 11575 6409
rect 11808 6412 12572 6440
rect 9640 6344 10548 6372
rect 9640 6332 9646 6344
rect 6089 6307 6147 6313
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6653 6307 6711 6313
rect 6653 6273 6665 6307
rect 6699 6304 6711 6307
rect 6699 6276 6914 6304
rect 6699 6273 6711 6276
rect 6653 6267 6711 6273
rect 6886 6236 6914 6276
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 8018 6304 8024 6316
rect 7616 6276 8024 6304
rect 7616 6264 7622 6276
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8404 6236 8432 6332
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6304 10195 6307
rect 10226 6304 10232 6316
rect 10183 6276 10232 6304
rect 10183 6273 10195 6276
rect 10137 6267 10195 6273
rect 10226 6264 10232 6276
rect 10284 6264 10290 6316
rect 10413 6307 10471 6313
rect 10413 6273 10425 6307
rect 10459 6304 10471 6307
rect 10502 6304 10508 6316
rect 10459 6276 10508 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 11333 6307 11391 6313
rect 11103 6276 11192 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 6886 6208 8432 6236
rect 3804 6140 6868 6168
rect 3973 6103 4031 6109
rect 3973 6069 3985 6103
rect 4019 6100 4031 6103
rect 4338 6100 4344 6112
rect 4019 6072 4344 6100
rect 4019 6069 4031 6072
rect 3973 6063 4031 6069
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 5997 6103 6055 6109
rect 5997 6069 6009 6103
rect 6043 6100 6055 6103
rect 6730 6100 6736 6112
rect 6043 6072 6736 6100
rect 6043 6069 6055 6072
rect 5997 6063 6055 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 6840 6100 6868 6140
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 11054 6168 11060 6180
rect 9640 6140 11060 6168
rect 9640 6128 9646 6140
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 11164 6177 11192 6276
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11348 6236 11376 6267
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 11808 6313 11836 6412
rect 12434 6372 12440 6384
rect 12268 6344 12440 6372
rect 12268 6313 12296 6344
rect 12434 6332 12440 6344
rect 12492 6332 12498 6384
rect 12544 6372 12572 6412
rect 12618 6400 12624 6452
rect 12676 6400 12682 6452
rect 12802 6440 12808 6452
rect 12728 6412 12808 6440
rect 12728 6372 12756 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 14645 6443 14703 6449
rect 14645 6440 14657 6443
rect 13044 6412 14657 6440
rect 13044 6400 13050 6412
rect 14645 6409 14657 6412
rect 14691 6409 14703 6443
rect 14645 6403 14703 6409
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6409 14979 6443
rect 14921 6403 14979 6409
rect 12544 6344 12756 6372
rect 14182 6332 14188 6384
rect 14240 6372 14246 6384
rect 14936 6372 14964 6403
rect 15102 6400 15108 6452
rect 15160 6440 15166 6452
rect 15160 6412 16252 6440
rect 15160 6400 15166 6412
rect 14240 6344 14412 6372
rect 14240 6332 14246 6344
rect 12813 6316 12871 6317
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 12618 6304 12624 6316
rect 12391 6276 12624 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 12802 6264 12808 6316
rect 12860 6271 12871 6316
rect 12860 6264 12866 6271
rect 13078 6264 13084 6316
rect 13136 6264 13142 6316
rect 13354 6264 13360 6316
rect 13412 6264 13418 6316
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14277 6307 14335 6313
rect 13955 6276 14136 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 12526 6236 12532 6248
rect 11348 6208 12532 6236
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12710 6196 12716 6248
rect 12768 6236 12774 6248
rect 12768 6208 13492 6236
rect 12768 6196 12774 6208
rect 11149 6171 11207 6177
rect 11149 6137 11161 6171
rect 11195 6137 11207 6171
rect 11149 6131 11207 6137
rect 11330 6128 11336 6180
rect 11388 6168 11394 6180
rect 13464 6177 13492 6208
rect 14108 6177 14136 6276
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 13173 6171 13231 6177
rect 13173 6168 13185 6171
rect 11388 6140 13185 6168
rect 11388 6128 11394 6140
rect 13173 6137 13185 6140
rect 13219 6137 13231 6171
rect 13173 6131 13231 6137
rect 13449 6171 13507 6177
rect 13449 6137 13461 6171
rect 13495 6137 13507 6171
rect 13449 6131 13507 6137
rect 14093 6171 14151 6177
rect 14093 6137 14105 6171
rect 14139 6137 14151 6171
rect 14292 6168 14320 6267
rect 14384 6236 14412 6344
rect 14568 6344 14964 6372
rect 15120 6344 15608 6372
rect 14568 6313 14596 6344
rect 15120 6313 15148 6344
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 15381 6307 15439 6313
rect 15381 6273 15393 6307
rect 15427 6273 15439 6307
rect 15381 6267 15439 6273
rect 14844 6236 14872 6267
rect 14384 6208 14872 6236
rect 15396 6168 15424 6267
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 14292 6140 15332 6168
rect 15396 6140 15485 6168
rect 14093 6131 14151 6137
rect 11698 6100 11704 6112
rect 6840 6072 11704 6100
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 11974 6060 11980 6112
rect 12032 6060 12038 6112
rect 12069 6103 12127 6109
rect 12069 6069 12081 6103
rect 12115 6100 12127 6103
rect 12158 6100 12164 6112
rect 12115 6072 12164 6100
rect 12115 6069 12127 6072
rect 12069 6063 12127 6069
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12526 6060 12532 6112
rect 12584 6060 12590 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12860 6072 12909 6100
rect 12860 6060 12866 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 13722 6060 13728 6112
rect 13780 6060 13786 6112
rect 14366 6060 14372 6112
rect 14424 6060 14430 6112
rect 15194 6060 15200 6112
rect 15252 6060 15258 6112
rect 15304 6100 15332 6140
rect 15473 6137 15485 6140
rect 15519 6137 15531 6171
rect 15580 6168 15608 6344
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16224 6313 16252 6412
rect 16942 6400 16948 6452
rect 17000 6400 17006 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15804 6276 15945 6304
rect 15804 6264 15810 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 16209 6307 16267 6313
rect 16209 6273 16221 6307
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 16850 6264 16856 6316
rect 16908 6264 16914 6316
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6304 17187 6307
rect 17236 6304 17264 6403
rect 17310 6400 17316 6452
rect 17368 6440 17374 6452
rect 19245 6443 19303 6449
rect 17368 6412 18828 6440
rect 17368 6400 17374 6412
rect 17420 6344 17908 6372
rect 17420 6313 17448 6344
rect 17175 6276 17264 6304
rect 17405 6307 17463 6313
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 17405 6273 17417 6307
rect 17451 6273 17463 6307
rect 17405 6267 17463 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17727 6276 17816 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 16025 6171 16083 6177
rect 16025 6168 16037 6171
rect 15580 6140 16037 6168
rect 15473 6131 15531 6137
rect 16025 6137 16037 6140
rect 16071 6137 16083 6171
rect 16025 6131 16083 6137
rect 16114 6128 16120 6180
rect 16172 6168 16178 6180
rect 16301 6171 16359 6177
rect 16301 6168 16313 6171
rect 16172 6140 16313 6168
rect 16172 6128 16178 6140
rect 16301 6137 16313 6140
rect 16347 6137 16359 6171
rect 16301 6131 16359 6137
rect 16666 6128 16672 6180
rect 16724 6128 16730 6180
rect 17494 6128 17500 6180
rect 17552 6128 17558 6180
rect 17788 6109 17816 6276
rect 17880 6168 17908 6344
rect 18414 6332 18420 6384
rect 18472 6372 18478 6384
rect 18472 6344 18644 6372
rect 18472 6332 18478 6344
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 17972 6236 18000 6267
rect 18046 6264 18052 6316
rect 18104 6304 18110 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18104 6276 18245 6304
rect 18104 6264 18110 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 18509 6307 18567 6313
rect 18509 6304 18521 6307
rect 18380 6276 18521 6304
rect 18380 6264 18386 6276
rect 18509 6273 18521 6276
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 18616 6236 18644 6344
rect 18800 6313 18828 6412
rect 19245 6409 19257 6443
rect 19291 6440 19303 6443
rect 19334 6440 19340 6452
rect 19291 6412 19340 6440
rect 19291 6409 19303 6412
rect 19245 6403 19303 6409
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 20070 6400 20076 6452
rect 20128 6440 20134 6452
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 20128 6412 20361 6440
rect 20128 6400 20134 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20901 6443 20959 6449
rect 20901 6440 20913 6443
rect 20496 6412 20913 6440
rect 20496 6400 20502 6412
rect 20901 6409 20913 6412
rect 20947 6409 20959 6443
rect 20901 6403 20959 6409
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 22189 6443 22247 6449
rect 22189 6440 22201 6443
rect 21324 6412 22201 6440
rect 21324 6400 21330 6412
rect 22189 6409 22201 6412
rect 22235 6409 22247 6443
rect 22189 6403 22247 6409
rect 22557 6443 22615 6449
rect 22557 6409 22569 6443
rect 22603 6409 22615 6443
rect 22557 6403 22615 6409
rect 18966 6332 18972 6384
rect 19024 6372 19030 6384
rect 19024 6344 19472 6372
rect 19024 6332 19030 6344
rect 19444 6313 19472 6344
rect 19518 6332 19524 6384
rect 19576 6372 19582 6384
rect 21082 6372 21088 6384
rect 19576 6344 21088 6372
rect 19576 6332 19582 6344
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 21358 6332 21364 6384
rect 21416 6372 21422 6384
rect 22572 6372 22600 6403
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23532 6412 23673 6440
rect 23532 6400 23538 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 23661 6403 23719 6409
rect 21416 6344 22600 6372
rect 21416 6332 21422 6344
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 19429 6307 19487 6313
rect 19429 6273 19441 6307
rect 19475 6273 19487 6307
rect 19429 6267 19487 6273
rect 19076 6236 19104 6267
rect 19702 6264 19708 6316
rect 19760 6264 19766 6316
rect 19886 6264 19892 6316
rect 19944 6304 19950 6316
rect 19981 6307 20039 6313
rect 19981 6304 19993 6307
rect 19944 6276 19993 6304
rect 19944 6264 19950 6276
rect 19981 6273 19993 6276
rect 20027 6273 20039 6307
rect 19981 6267 20039 6273
rect 20254 6264 20260 6316
rect 20312 6264 20318 6316
rect 20806 6264 20812 6316
rect 20864 6264 20870 6316
rect 21450 6264 21456 6316
rect 21508 6264 21514 6316
rect 21542 6264 21548 6316
rect 21600 6304 21606 6316
rect 21913 6307 21971 6313
rect 21913 6304 21925 6307
rect 21600 6276 21925 6304
rect 21600 6264 21606 6276
rect 21913 6273 21925 6276
rect 21959 6273 21971 6307
rect 21913 6267 21971 6273
rect 22462 6264 22468 6316
rect 22520 6264 22526 6316
rect 23014 6264 23020 6316
rect 23072 6264 23078 6316
rect 23569 6307 23627 6313
rect 23569 6273 23581 6307
rect 23615 6304 23627 6307
rect 24026 6304 24032 6316
rect 23615 6276 24032 6304
rect 23615 6273 23627 6276
rect 23569 6267 23627 6273
rect 24026 6264 24032 6276
rect 24084 6264 24090 6316
rect 17972 6208 18368 6236
rect 18616 6208 19104 6236
rect 18340 6177 18368 6208
rect 18049 6171 18107 6177
rect 18049 6168 18061 6171
rect 17880 6140 18061 6168
rect 18049 6137 18061 6140
rect 18095 6137 18107 6171
rect 18049 6131 18107 6137
rect 18325 6171 18383 6177
rect 18325 6137 18337 6171
rect 18371 6137 18383 6171
rect 18325 6131 18383 6137
rect 18414 6128 18420 6180
rect 18472 6168 18478 6180
rect 19521 6171 19579 6177
rect 19521 6168 19533 6171
rect 18472 6140 19533 6168
rect 18472 6128 18478 6140
rect 19521 6137 19533 6140
rect 19567 6137 19579 6171
rect 19521 6131 19579 6137
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 15304 6072 15761 6100
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 15749 6063 15807 6069
rect 17773 6103 17831 6109
rect 17773 6069 17785 6103
rect 17819 6069 17831 6103
rect 17773 6063 17831 6069
rect 18598 6060 18604 6112
rect 18656 6060 18662 6112
rect 18874 6060 18880 6112
rect 18932 6060 18938 6112
rect 19610 6060 19616 6112
rect 19668 6100 19674 6112
rect 19797 6103 19855 6109
rect 19797 6100 19809 6103
rect 19668 6072 19809 6100
rect 19668 6060 19674 6072
rect 19797 6069 19809 6072
rect 19843 6069 19855 6103
rect 19797 6063 19855 6069
rect 21634 6060 21640 6112
rect 21692 6060 21698 6112
rect 21818 6060 21824 6112
rect 21876 6100 21882 6112
rect 23109 6103 23167 6109
rect 23109 6100 23121 6103
rect 21876 6072 23121 6100
rect 21876 6060 21882 6072
rect 23109 6069 23121 6072
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5896 1823 5899
rect 2130 5896 2136 5908
rect 1811 5868 2136 5896
rect 1811 5865 1823 5868
rect 1765 5859 1823 5865
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 2314 5856 2320 5908
rect 2372 5856 2378 5908
rect 2682 5856 2688 5908
rect 2740 5856 2746 5908
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3844 5868 4077 5896
rect 3844 5856 3850 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4430 5856 4436 5908
rect 4488 5896 4494 5908
rect 4525 5899 4583 5905
rect 4525 5896 4537 5899
rect 4488 5868 4537 5896
rect 4488 5856 4494 5868
rect 4525 5865 4537 5868
rect 4571 5865 4583 5899
rect 4525 5859 4583 5865
rect 4798 5856 4804 5908
rect 4856 5856 4862 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 5994 5856 6000 5908
rect 6052 5856 6058 5908
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 7374 5896 7380 5908
rect 6886 5868 7380 5896
rect 4816 5828 4844 5856
rect 1872 5800 4844 5828
rect 5813 5831 5871 5837
rect 1872 5701 1900 5800
rect 5813 5797 5825 5831
rect 5859 5828 5871 5831
rect 6886 5828 6914 5868
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7926 5856 7932 5908
rect 7984 5856 7990 5908
rect 8110 5856 8116 5908
rect 8168 5856 8174 5908
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 8389 5899 8447 5905
rect 8389 5896 8401 5899
rect 8260 5868 8401 5896
rect 8260 5856 8266 5868
rect 8389 5865 8401 5868
rect 8435 5865 8447 5899
rect 8389 5859 8447 5865
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 9030 5856 9036 5908
rect 9088 5896 9094 5908
rect 9125 5899 9183 5905
rect 9125 5896 9137 5899
rect 9088 5868 9137 5896
rect 9088 5856 9094 5868
rect 9125 5865 9137 5868
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 9214 5856 9220 5908
rect 9272 5896 9278 5908
rect 9401 5899 9459 5905
rect 9401 5896 9413 5899
rect 9272 5868 9413 5896
rect 9272 5856 9278 5868
rect 9401 5865 9413 5868
rect 9447 5865 9459 5899
rect 9401 5859 9459 5865
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 12308 5868 12633 5896
rect 12308 5856 12314 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 12621 5859 12679 5865
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 14645 5899 14703 5905
rect 14645 5896 14657 5899
rect 13136 5868 14657 5896
rect 13136 5856 13142 5868
rect 14645 5865 14657 5868
rect 14691 5865 14703 5899
rect 14645 5859 14703 5865
rect 14734 5856 14740 5908
rect 14792 5896 14798 5908
rect 15381 5899 15439 5905
rect 15381 5896 15393 5899
rect 14792 5868 15393 5896
rect 14792 5856 14798 5868
rect 15381 5865 15393 5868
rect 15427 5865 15439 5899
rect 15381 5859 15439 5865
rect 15654 5856 15660 5908
rect 15712 5856 15718 5908
rect 15764 5868 16252 5896
rect 5859 5800 6914 5828
rect 5859 5797 5871 5800
rect 5813 5791 5871 5797
rect 7190 5788 7196 5840
rect 7248 5788 7254 5840
rect 8128 5760 8156 5856
rect 8680 5828 8708 5856
rect 9858 5828 9864 5840
rect 8680 5800 9864 5828
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5797 10011 5831
rect 9953 5791 10011 5797
rect 9490 5760 9496 5772
rect 2976 5732 5304 5760
rect 2976 5701 3004 5732
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 4522 5692 4528 5704
rect 3559 5664 4528 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 2409 5627 2467 5633
rect 2409 5593 2421 5627
rect 2455 5624 2467 5627
rect 3436 5624 3464 5652
rect 2455 5596 3464 5624
rect 4341 5627 4399 5633
rect 2455 5593 2467 5596
rect 2409 5587 2467 5593
rect 4341 5593 4353 5627
rect 4387 5593 4399 5627
rect 4341 5587 4399 5593
rect 4356 5556 4384 5587
rect 5166 5584 5172 5636
rect 5224 5584 5230 5636
rect 5276 5624 5304 5732
rect 5644 5732 8156 5760
rect 9324 5732 9496 5760
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 5644 5701 5672 5732
rect 9324 5701 9352 5732
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9968 5760 9996 5791
rect 10042 5788 10048 5840
rect 10100 5828 10106 5840
rect 10229 5831 10287 5837
rect 10229 5828 10241 5831
rect 10100 5800 10241 5828
rect 10100 5788 10106 5800
rect 10229 5797 10241 5800
rect 10275 5797 10287 5831
rect 10229 5791 10287 5797
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11333 5831 11391 5837
rect 11333 5828 11345 5831
rect 11112 5800 11345 5828
rect 11112 5788 11118 5800
rect 11333 5797 11345 5800
rect 11379 5797 11391 5831
rect 12161 5831 12219 5837
rect 12161 5828 12173 5831
rect 11333 5791 11391 5797
rect 11808 5800 12173 5828
rect 11808 5760 11836 5800
rect 12161 5797 12173 5800
rect 12207 5797 12219 5831
rect 15764 5828 15792 5868
rect 16224 5837 16252 5868
rect 16482 5856 16488 5908
rect 16540 5856 16546 5908
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 16945 5899 17003 5905
rect 16945 5896 16957 5899
rect 16908 5868 16957 5896
rect 16908 5856 16914 5868
rect 16945 5865 16957 5868
rect 16991 5865 17003 5899
rect 16945 5859 17003 5865
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17589 5899 17647 5905
rect 17589 5896 17601 5899
rect 17460 5868 17601 5896
rect 17460 5856 17466 5868
rect 17589 5865 17601 5868
rect 17635 5865 17647 5899
rect 17589 5859 17647 5865
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 18322 5896 18328 5908
rect 17828 5868 18328 5896
rect 17828 5856 17834 5868
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 18417 5899 18475 5905
rect 18417 5865 18429 5899
rect 18463 5896 18475 5899
rect 18782 5896 18788 5908
rect 18463 5868 18788 5896
rect 18463 5865 18475 5868
rect 18417 5859 18475 5865
rect 18782 5856 18788 5868
rect 18840 5856 18846 5908
rect 18874 5856 18880 5908
rect 18932 5856 18938 5908
rect 19245 5899 19303 5905
rect 19245 5865 19257 5899
rect 19291 5896 19303 5899
rect 19334 5896 19340 5908
rect 19291 5868 19340 5896
rect 19291 5865 19303 5868
rect 19245 5859 19303 5865
rect 19334 5856 19340 5868
rect 19392 5856 19398 5908
rect 19518 5856 19524 5908
rect 19576 5856 19582 5908
rect 19610 5856 19616 5908
rect 19668 5856 19674 5908
rect 21453 5899 21511 5905
rect 21453 5896 21465 5899
rect 20364 5868 21465 5896
rect 12161 5791 12219 5797
rect 13096 5800 15792 5828
rect 15933 5831 15991 5837
rect 9600 5732 9996 5760
rect 10060 5732 11836 5760
rect 9600 5701 9628 5732
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 9309 5695 9367 5701
rect 5629 5655 5687 5661
rect 5736 5664 9260 5692
rect 5736 5624 5764 5664
rect 5276 5596 5764 5624
rect 6270 5584 6276 5636
rect 6328 5584 6334 5636
rect 6825 5627 6883 5633
rect 6825 5593 6837 5627
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 4356 5528 5365 5556
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 6840 5556 6868 5587
rect 7374 5584 7380 5636
rect 7432 5584 7438 5636
rect 7834 5584 7840 5636
rect 7892 5584 7898 5636
rect 8662 5584 8668 5636
rect 8720 5584 8726 5636
rect 9122 5584 9128 5636
rect 9180 5584 9186 5636
rect 9232 5624 9260 5664
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5692 9735 5695
rect 9950 5692 9956 5704
rect 9723 5664 9956 5692
rect 9723 5661 9735 5664
rect 9677 5655 9735 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10060 5624 10088 5732
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12032 5732 12388 5760
rect 12032 5720 12038 5732
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 9232 5596 10088 5624
rect 10152 5624 10180 5655
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5692 10747 5695
rect 10870 5692 10876 5704
rect 10735 5664 10876 5692
rect 10735 5661 10747 5664
rect 10689 5655 10747 5661
rect 10870 5652 10876 5664
rect 10928 5652 10934 5704
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11054 5692 11060 5704
rect 11011 5664 11060 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5692 11299 5695
rect 11330 5692 11336 5704
rect 11287 5664 11336 5692
rect 11287 5661 11299 5664
rect 11241 5655 11299 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11514 5652 11520 5704
rect 11572 5652 11578 5704
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 12066 5652 12072 5704
rect 12124 5652 12130 5704
rect 12360 5701 12388 5732
rect 12526 5720 12532 5772
rect 12584 5720 12590 5772
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 13096 5760 13124 5800
rect 15933 5797 15945 5831
rect 15979 5797 15991 5831
rect 15933 5791 15991 5797
rect 16209 5831 16267 5837
rect 16209 5797 16221 5831
rect 16255 5797 16267 5831
rect 16209 5791 16267 5797
rect 15948 5760 15976 5791
rect 16298 5788 16304 5840
rect 16356 5828 16362 5840
rect 16356 5800 17080 5828
rect 16356 5788 16362 5800
rect 12768 5732 13124 5760
rect 15580 5732 15976 5760
rect 16132 5732 16896 5760
rect 12768 5720 12774 5732
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5661 12403 5695
rect 12544 5692 12572 5720
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12544 5664 12817 5692
rect 12345 5655 12403 5661
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 13078 5652 13084 5704
rect 13136 5688 13142 5704
rect 13173 5695 13231 5701
rect 13173 5688 13185 5695
rect 13136 5661 13185 5688
rect 13219 5661 13231 5695
rect 13136 5660 13231 5661
rect 13136 5652 13142 5660
rect 13173 5655 13231 5660
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14332 5664 14565 5692
rect 14332 5652 14338 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 15580 5701 15608 5732
rect 16132 5701 16160 5732
rect 15565 5695 15623 5701
rect 15565 5661 15577 5695
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5661 15899 5695
rect 15841 5655 15899 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16393 5695 16451 5701
rect 16393 5692 16405 5695
rect 16117 5655 16175 5661
rect 16224 5664 16405 5692
rect 10152 5596 13124 5624
rect 9140 5556 9168 5584
rect 6840 5528 9168 5556
rect 5353 5519 5411 5525
rect 9858 5516 9864 5568
rect 9916 5516 9922 5568
rect 9950 5516 9956 5568
rect 10008 5556 10014 5568
rect 10505 5559 10563 5565
rect 10505 5556 10517 5559
rect 10008 5528 10517 5556
rect 10008 5516 10014 5528
rect 10505 5525 10517 5528
rect 10551 5525 10563 5559
rect 10505 5519 10563 5525
rect 10778 5516 10784 5568
rect 10836 5516 10842 5568
rect 11054 5516 11060 5568
rect 11112 5516 11118 5568
rect 11606 5516 11612 5568
rect 11664 5516 11670 5568
rect 11698 5516 11704 5568
rect 11756 5556 11762 5568
rect 11885 5559 11943 5565
rect 11885 5556 11897 5559
rect 11756 5528 11897 5556
rect 11756 5516 11762 5528
rect 11885 5525 11897 5528
rect 11931 5525 11943 5559
rect 11885 5519 11943 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12989 5559 13047 5565
rect 12989 5556 13001 5559
rect 12032 5528 13001 5556
rect 12032 5516 12038 5528
rect 12989 5525 13001 5528
rect 13035 5525 13047 5559
rect 13096 5556 13124 5596
rect 15470 5584 15476 5636
rect 15528 5624 15534 5636
rect 15856 5624 15884 5655
rect 15528 5596 15884 5624
rect 15528 5584 15534 5596
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 13096 5528 13277 5556
rect 12989 5519 13047 5525
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13265 5519 13323 5525
rect 13998 5516 14004 5568
rect 14056 5556 14062 5568
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 14056 5528 14381 5556
rect 14056 5516 14062 5528
rect 14369 5525 14381 5528
rect 14415 5525 14427 5559
rect 14369 5519 14427 5525
rect 15654 5516 15660 5568
rect 15712 5556 15718 5568
rect 16224 5556 16252 5664
rect 16393 5661 16405 5664
rect 16439 5661 16451 5695
rect 16393 5655 16451 5661
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 16540 5664 16681 5692
rect 16540 5652 16546 5664
rect 16669 5661 16681 5664
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 16761 5695 16819 5701
rect 16761 5661 16773 5695
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 16298 5584 16304 5636
rect 16356 5624 16362 5636
rect 16776 5624 16804 5655
rect 16356 5596 16804 5624
rect 16868 5624 16896 5732
rect 17052 5692 17080 5800
rect 17310 5788 17316 5840
rect 17368 5788 17374 5840
rect 18598 5828 18604 5840
rect 17512 5800 18604 5828
rect 17512 5701 17540 5800
rect 18598 5788 18604 5800
rect 18656 5788 18662 5840
rect 18693 5831 18751 5837
rect 18693 5797 18705 5831
rect 18739 5797 18751 5831
rect 18693 5791 18751 5797
rect 18708 5760 18736 5791
rect 18892 5760 18920 5856
rect 18064 5732 18736 5760
rect 18800 5732 18920 5760
rect 18064 5701 18092 5732
rect 17221 5695 17279 5701
rect 17221 5692 17233 5695
rect 17052 5664 17233 5692
rect 17221 5661 17233 5664
rect 17267 5661 17279 5695
rect 17221 5655 17279 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5692 18383 5695
rect 18414 5692 18420 5704
rect 18371 5664 18420 5692
rect 18371 5661 18383 5664
rect 18325 5655 18383 5661
rect 17788 5624 17816 5655
rect 18414 5652 18420 5664
rect 18472 5652 18478 5704
rect 18598 5652 18604 5704
rect 18656 5652 18662 5704
rect 18800 5624 18828 5732
rect 18877 5695 18935 5701
rect 18877 5661 18889 5695
rect 18923 5661 18935 5695
rect 18877 5655 18935 5661
rect 19429 5695 19487 5701
rect 19429 5661 19441 5695
rect 19475 5692 19487 5695
rect 19628 5692 19656 5856
rect 19797 5831 19855 5837
rect 19797 5797 19809 5831
rect 19843 5797 19855 5831
rect 19797 5791 19855 5797
rect 19475 5664 19656 5692
rect 19705 5695 19763 5701
rect 19475 5661 19487 5664
rect 19429 5655 19487 5661
rect 19705 5661 19717 5695
rect 19751 5692 19763 5695
rect 19812 5692 19840 5791
rect 20364 5760 20392 5868
rect 21453 5865 21465 5868
rect 21499 5865 21511 5899
rect 21453 5859 21511 5865
rect 21634 5856 21640 5908
rect 21692 5896 21698 5908
rect 21692 5868 22094 5896
rect 21692 5856 21698 5868
rect 20533 5831 20591 5837
rect 20533 5797 20545 5831
rect 20579 5797 20591 5831
rect 20533 5791 20591 5797
rect 20272 5732 20392 5760
rect 19751 5664 19840 5692
rect 19751 5661 19763 5664
rect 19705 5655 19763 5661
rect 16868 5596 17080 5624
rect 17788 5596 18828 5624
rect 16356 5584 16362 5596
rect 17052 5565 17080 5596
rect 15712 5528 16252 5556
rect 17037 5559 17095 5565
rect 15712 5516 15718 5528
rect 17037 5525 17049 5559
rect 17083 5525 17095 5559
rect 17037 5519 17095 5525
rect 17862 5516 17868 5568
rect 17920 5516 17926 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18141 5559 18199 5565
rect 18141 5556 18153 5559
rect 18012 5528 18153 5556
rect 18012 5516 18018 5528
rect 18141 5525 18153 5528
rect 18187 5525 18199 5559
rect 18141 5519 18199 5525
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 18892 5556 18920 5655
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 20272 5701 20300 5732
rect 20257 5695 20315 5701
rect 20257 5661 20269 5695
rect 20303 5661 20315 5695
rect 20257 5655 20315 5661
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5661 20407 5695
rect 20548 5692 20576 5791
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21177 5831 21235 5837
rect 21177 5828 21189 5831
rect 20680 5800 21189 5828
rect 20680 5788 20686 5800
rect 21177 5797 21189 5800
rect 21223 5797 21235 5831
rect 21177 5791 21235 5797
rect 20809 5695 20867 5701
rect 20809 5692 20821 5695
rect 20548 5664 20821 5692
rect 20349 5655 20407 5661
rect 20809 5661 20821 5664
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 20364 5624 20392 5655
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21637 5695 21695 5701
rect 21637 5692 21649 5695
rect 21140 5664 21649 5692
rect 21140 5652 21146 5664
rect 21637 5661 21649 5664
rect 21683 5661 21695 5695
rect 22066 5692 22094 5868
rect 22278 5856 22284 5908
rect 22336 5896 22342 5908
rect 22557 5899 22615 5905
rect 22557 5896 22569 5899
rect 22336 5868 22569 5896
rect 22336 5856 22342 5868
rect 22557 5865 22569 5868
rect 22603 5865 22615 5899
rect 22557 5859 22615 5865
rect 22830 5856 22836 5908
rect 22888 5896 22894 5908
rect 23109 5899 23167 5905
rect 23109 5896 23121 5899
rect 22888 5868 23121 5896
rect 22888 5856 22894 5868
rect 23109 5865 23121 5868
rect 23155 5865 23167 5899
rect 23109 5859 23167 5865
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 23661 5899 23719 5905
rect 23661 5896 23673 5899
rect 23532 5868 23673 5896
rect 23532 5856 23538 5868
rect 23661 5865 23673 5868
rect 23707 5865 23719 5899
rect 23661 5859 23719 5865
rect 25590 5856 25596 5908
rect 25648 5856 25654 5908
rect 22189 5831 22247 5837
rect 22189 5797 22201 5831
rect 22235 5828 22247 5831
rect 25608 5828 25636 5856
rect 22235 5800 25636 5828
rect 22235 5797 22247 5800
rect 22189 5791 22247 5797
rect 24213 5695 24271 5701
rect 24213 5692 24225 5695
rect 22066 5664 24225 5692
rect 21637 5655 21695 5661
rect 24213 5661 24225 5664
rect 24259 5661 24271 5695
rect 24213 5655 24271 5661
rect 20898 5624 20904 5636
rect 20364 5596 20904 5624
rect 20898 5584 20904 5596
rect 20956 5584 20962 5636
rect 20990 5584 20996 5636
rect 21048 5584 21054 5636
rect 21910 5584 21916 5636
rect 21968 5584 21974 5636
rect 22462 5584 22468 5636
rect 22520 5584 22526 5636
rect 23014 5584 23020 5636
rect 23072 5584 23078 5636
rect 23569 5627 23627 5633
rect 23569 5593 23581 5627
rect 23615 5624 23627 5627
rect 23934 5624 23940 5636
rect 23615 5596 23940 5624
rect 23615 5593 23627 5596
rect 23569 5587 23627 5593
rect 23934 5584 23940 5596
rect 23992 5584 23998 5636
rect 18380 5528 18920 5556
rect 18380 5516 18386 5528
rect 20070 5516 20076 5568
rect 20128 5516 20134 5568
rect 20622 5516 20628 5568
rect 20680 5516 20686 5568
rect 24026 5516 24032 5568
rect 24084 5516 24090 5568
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 1854 5312 1860 5364
rect 1912 5312 1918 5364
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 3602 5352 3608 5364
rect 3467 5324 3608 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 3697 5355 3755 5361
rect 3697 5321 3709 5355
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 2133 5287 2191 5293
rect 2133 5284 2145 5287
rect 1636 5256 2145 5284
rect 1636 5244 1642 5256
rect 2133 5253 2145 5256
rect 2179 5253 2191 5287
rect 2133 5247 2191 5253
rect 3053 5287 3111 5293
rect 3053 5253 3065 5287
rect 3099 5284 3111 5287
rect 3712 5284 3740 5315
rect 4338 5312 4344 5364
rect 4396 5312 4402 5364
rect 4522 5312 4528 5364
rect 4580 5312 4586 5364
rect 4893 5355 4951 5361
rect 4893 5321 4905 5355
rect 4939 5321 4951 5355
rect 4893 5315 4951 5321
rect 3099 5256 3740 5284
rect 4356 5284 4384 5312
rect 4617 5287 4675 5293
rect 4356 5256 4568 5284
rect 3099 5253 3111 5256
rect 3053 5247 3111 5253
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 2498 5176 2504 5228
rect 2556 5176 2562 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 290 5108 296 5160
rect 348 5148 354 5160
rect 2777 5151 2835 5157
rect 2777 5148 2789 5151
rect 348 5120 2789 5148
rect 348 5108 354 5120
rect 2777 5117 2789 5120
rect 2823 5117 2835 5151
rect 3620 5148 3648 5179
rect 3694 5176 3700 5228
rect 3752 5216 3758 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3752 5188 3893 5216
rect 3752 5176 3758 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5216 4215 5219
rect 4430 5216 4436 5228
rect 4203 5188 4436 5216
rect 4203 5185 4215 5188
rect 4157 5179 4215 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4540 5216 4568 5256
rect 4617 5253 4629 5287
rect 4663 5284 4675 5287
rect 4908 5284 4936 5315
rect 5166 5312 5172 5364
rect 5224 5312 5230 5364
rect 5537 5355 5595 5361
rect 5537 5321 5549 5355
rect 5583 5321 5595 5355
rect 5537 5315 5595 5321
rect 4663 5256 4936 5284
rect 4663 5253 4675 5256
rect 4617 5247 4675 5253
rect 5077 5219 5135 5225
rect 5077 5216 5089 5219
rect 4540 5188 5089 5216
rect 5077 5185 5089 5188
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 5552 5216 5580 5315
rect 5810 5312 5816 5364
rect 5868 5312 5874 5364
rect 6365 5355 6423 5361
rect 6365 5321 6377 5355
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 7285 5355 7343 5361
rect 6963 5324 7052 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 5399 5188 5580 5216
rect 5721 5219 5779 5225
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6380 5216 6408 5315
rect 7024 5284 7052 5324
rect 7285 5321 7297 5355
rect 7331 5352 7343 5355
rect 7374 5352 7380 5364
rect 7331 5324 7380 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 7561 5355 7619 5361
rect 7561 5352 7573 5355
rect 7524 5324 7573 5352
rect 7524 5312 7530 5324
rect 7561 5321 7573 5324
rect 7607 5321 7619 5355
rect 7561 5315 7619 5321
rect 7834 5312 7840 5364
rect 7892 5312 7898 5364
rect 8570 5352 8576 5364
rect 8036 5324 8576 5352
rect 6043 5188 6408 5216
rect 6472 5256 6684 5284
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 5258 5148 5264 5160
rect 3620 5120 5264 5148
rect 2777 5111 2835 5117
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5534 5108 5540 5160
rect 5592 5108 5598 5160
rect 5736 5148 5764 5179
rect 6472 5148 6500 5256
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 5736 5120 6500 5148
rect 5552 5080 5580 5108
rect 6564 5080 6592 5179
rect 6656 5148 6684 5256
rect 6840 5256 6960 5284
rect 7024 5256 7328 5284
rect 6840 5225 6868 5256
rect 6825 5219 6883 5225
rect 6825 5185 6837 5219
rect 6871 5185 6883 5219
rect 6932 5220 6960 5256
rect 7300 5228 7328 5256
rect 6932 5192 7052 5220
rect 6825 5179 6883 5185
rect 7024 5160 7052 5192
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7190 5216 7196 5228
rect 7147 5188 7196 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7469 5219 7527 5225
rect 7469 5185 7481 5219
rect 7515 5216 7527 5219
rect 7650 5216 7656 5228
rect 7515 5188 7656 5216
rect 7515 5185 7527 5188
rect 7469 5179 7527 5185
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 8036 5225 8064 5324
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 8662 5312 8668 5364
rect 8720 5312 8726 5364
rect 9125 5355 9183 5361
rect 9125 5321 9137 5355
rect 9171 5352 9183 5355
rect 9306 5352 9312 5364
rect 9171 5324 9312 5352
rect 9171 5321 9183 5324
rect 9125 5315 9183 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 10134 5312 10140 5364
rect 10192 5312 10198 5364
rect 10229 5355 10287 5361
rect 10229 5321 10241 5355
rect 10275 5321 10287 5355
rect 10229 5315 10287 5321
rect 9766 5284 9772 5296
rect 8588 5256 9772 5284
rect 8588 5225 8616 5256
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8573 5219 8631 5225
rect 8343 5188 8432 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 6914 5148 6920 5160
rect 6656 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7006 5108 7012 5160
rect 7064 5108 7070 5160
rect 7392 5120 8340 5148
rect 7392 5080 7420 5120
rect 5552 5052 6132 5080
rect 6564 5052 7420 5080
rect 7484 5052 8156 5080
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3568 4984 3985 5012
rect 3568 4972 3574 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 6104 5012 6132 5052
rect 6641 5015 6699 5021
rect 6641 5012 6653 5015
rect 6104 4984 6653 5012
rect 3973 4975 4031 4981
rect 6641 4981 6653 4984
rect 6687 4981 6699 5015
rect 6641 4975 6699 4981
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7484 5012 7512 5052
rect 8128 5021 8156 5052
rect 6788 4984 7512 5012
rect 8113 5015 8171 5021
rect 6788 4972 6794 4984
rect 8113 4981 8125 5015
rect 8159 4981 8171 5015
rect 8312 5012 8340 5120
rect 8404 5089 8432 5188
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8849 5219 8907 5225
rect 8849 5185 8861 5219
rect 8895 5185 8907 5219
rect 8849 5179 8907 5185
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 8389 5083 8447 5089
rect 8389 5049 8401 5083
rect 8435 5049 8447 5083
rect 8864 5080 8892 5179
rect 9324 5148 9352 5179
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9640 5188 9689 5216
rect 9640 5176 9646 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9876 5216 9904 5312
rect 10244 5228 10272 5315
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 17862 5352 17868 5364
rect 12400 5324 17868 5352
rect 12400 5312 12406 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18598 5312 18604 5364
rect 18656 5352 18662 5364
rect 18693 5355 18751 5361
rect 18693 5352 18705 5355
rect 18656 5324 18705 5352
rect 18656 5312 18662 5324
rect 18693 5321 18705 5324
rect 18739 5321 18751 5355
rect 18693 5315 18751 5321
rect 18969 5355 19027 5361
rect 18969 5321 18981 5355
rect 19015 5352 19027 5355
rect 19242 5352 19248 5364
rect 19015 5324 19248 5352
rect 19015 5321 19027 5324
rect 18969 5315 19027 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19521 5355 19579 5361
rect 19521 5321 19533 5355
rect 19567 5352 19579 5355
rect 19978 5352 19984 5364
rect 19567 5324 19984 5352
rect 19567 5321 19579 5324
rect 19521 5315 19579 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20070 5312 20076 5364
rect 20128 5312 20134 5364
rect 20901 5355 20959 5361
rect 20901 5321 20913 5355
rect 20947 5352 20959 5355
rect 21450 5352 21456 5364
rect 20947 5324 21456 5352
rect 20947 5321 20959 5324
rect 20901 5315 20959 5321
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21910 5352 21916 5364
rect 21683 5324 21916 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 23566 5312 23572 5364
rect 23624 5352 23630 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 23624 5324 23857 5352
rect 23624 5312 23630 5324
rect 23845 5321 23857 5324
rect 23891 5321 23903 5355
rect 23845 5315 23903 5321
rect 10336 5256 10640 5284
rect 9953 5219 10011 5225
rect 9953 5216 9965 5219
rect 9876 5188 9965 5216
rect 9677 5179 9735 5185
rect 9953 5185 9965 5188
rect 9999 5185 10011 5219
rect 9953 5179 10011 5185
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10336 5148 10364 5256
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 9324 5120 10364 5148
rect 10502 5108 10508 5160
rect 10560 5108 10566 5160
rect 10612 5148 10640 5256
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10744 5188 10977 5216
rect 10744 5176 10750 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 11072 5216 11100 5312
rect 18414 5244 18420 5296
rect 18472 5284 18478 5296
rect 18472 5256 18828 5284
rect 18472 5244 18478 5256
rect 11241 5219 11299 5225
rect 11241 5216 11253 5219
rect 11072 5188 11253 5216
rect 10965 5179 11023 5185
rect 11241 5185 11253 5188
rect 11287 5185 11299 5219
rect 11241 5179 11299 5185
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11480 5188 11713 5216
rect 11480 5176 11486 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 18506 5176 18512 5228
rect 18564 5176 18570 5228
rect 18800 5225 18828 5256
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 19058 5176 19064 5228
rect 19116 5176 19122 5228
rect 19334 5176 19340 5228
rect 19392 5176 19398 5228
rect 19794 5176 19800 5228
rect 19852 5176 19858 5228
rect 20088 5216 20116 5312
rect 20162 5244 20168 5296
rect 20220 5284 20226 5296
rect 22097 5287 22155 5293
rect 22097 5284 22109 5287
rect 20220 5256 21404 5284
rect 20220 5244 20226 5256
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 20088 5188 20269 5216
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 20441 5219 20499 5225
rect 20441 5185 20453 5219
rect 20487 5185 20499 5219
rect 20441 5179 20499 5185
rect 16666 5148 16672 5160
rect 10612 5120 16672 5148
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 20456 5148 20484 5179
rect 20714 5176 20720 5228
rect 20772 5176 20778 5228
rect 21376 5225 21404 5256
rect 21652 5256 22109 5284
rect 21652 5228 21680 5256
rect 22097 5253 22109 5256
rect 22143 5253 22155 5287
rect 22097 5247 22155 5253
rect 23477 5287 23535 5293
rect 23477 5253 23489 5287
rect 23523 5284 23535 5287
rect 24026 5284 24032 5296
rect 23523 5256 24032 5284
rect 23523 5253 23535 5256
rect 23477 5247 23535 5253
rect 24026 5244 24032 5256
rect 24084 5244 24090 5296
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 21450 5176 21456 5228
rect 21508 5176 21514 5228
rect 21634 5176 21640 5228
rect 21692 5176 21698 5228
rect 22922 5176 22928 5228
rect 22980 5176 22986 5228
rect 23750 5176 23756 5228
rect 23808 5176 23814 5228
rect 19996 5120 20484 5148
rect 22373 5151 22431 5157
rect 9674 5080 9680 5092
rect 8864 5052 9680 5080
rect 8389 5043 8447 5049
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 9861 5083 9919 5089
rect 9861 5049 9873 5083
rect 9907 5080 9919 5083
rect 10520 5080 10548 5108
rect 11517 5083 11575 5089
rect 11517 5080 11529 5083
rect 9907 5052 10548 5080
rect 10612 5052 11529 5080
rect 9907 5049 9919 5052
rect 9861 5043 9919 5049
rect 10612 5012 10640 5052
rect 11517 5049 11529 5052
rect 11563 5049 11575 5083
rect 11517 5043 11575 5049
rect 19245 5083 19303 5089
rect 19245 5049 19257 5083
rect 19291 5080 19303 5083
rect 19886 5080 19892 5092
rect 19291 5052 19892 5080
rect 19291 5049 19303 5052
rect 19245 5043 19303 5049
rect 19886 5040 19892 5052
rect 19944 5040 19950 5092
rect 19996 5089 20024 5120
rect 22373 5117 22385 5151
rect 22419 5148 22431 5151
rect 22649 5151 22707 5157
rect 22419 5120 22600 5148
rect 22419 5117 22431 5120
rect 22373 5111 22431 5117
rect 19981 5083 20039 5089
rect 19981 5049 19993 5083
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 20070 5040 20076 5092
rect 20128 5040 20134 5092
rect 22572 5080 22600 5120
rect 22649 5117 22661 5151
rect 22695 5148 22707 5151
rect 25038 5148 25044 5160
rect 22695 5120 25044 5148
rect 22695 5117 22707 5120
rect 22649 5111 22707 5117
rect 25038 5108 25044 5120
rect 25096 5108 25102 5160
rect 23842 5080 23848 5092
rect 20640 5052 21404 5080
rect 22572 5052 23848 5080
rect 8312 4984 10640 5012
rect 8113 4975 8171 4981
rect 10778 4972 10784 5024
rect 10836 4972 10842 5024
rect 11057 5015 11115 5021
rect 11057 4981 11069 5015
rect 11103 5012 11115 5015
rect 11146 5012 11152 5024
rect 11103 4984 11152 5012
rect 11103 4981 11115 4984
rect 11057 4975 11115 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 20254 5012 20260 5024
rect 18564 4984 20260 5012
rect 18564 4972 18570 4984
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 20640 5021 20668 5052
rect 20625 5015 20683 5021
rect 20625 4981 20637 5015
rect 20671 4981 20683 5015
rect 20625 4975 20683 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 20956 4984 21189 5012
rect 20956 4972 20962 4984
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 21376 5012 21404 5052
rect 23842 5040 23848 5052
rect 23900 5040 23906 5092
rect 22462 5012 22468 5024
rect 21376 4984 22468 5012
rect 21177 4975 21235 4981
rect 22462 4972 22468 4984
rect 22520 4972 22526 5024
rect 23385 5015 23443 5021
rect 23385 4981 23397 5015
rect 23431 5012 23443 5015
rect 24302 5012 24308 5024
rect 23431 4984 24308 5012
rect 23431 4981 23443 4984
rect 23385 4975 23443 4981
rect 24302 4972 24308 4984
rect 24360 4972 24366 5024
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1360 4780 1501 4808
rect 1360 4768 1366 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4777 2191 4811
rect 2133 4771 2191 4777
rect 750 4700 756 4752
rect 808 4740 814 4752
rect 2148 4740 2176 4771
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2593 4811 2651 4817
rect 2593 4808 2605 4811
rect 2280 4780 2605 4808
rect 2280 4768 2286 4780
rect 2593 4777 2605 4780
rect 2639 4777 2651 4811
rect 2593 4771 2651 4777
rect 3053 4811 3111 4817
rect 3053 4777 3065 4811
rect 3099 4808 3111 4811
rect 3694 4808 3700 4820
rect 3099 4780 3700 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4488 4780 4629 4808
rect 4488 4768 4494 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 6730 4808 6736 4820
rect 5316 4780 6736 4808
rect 5316 4768 5322 4780
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 12158 4808 12164 4820
rect 7064 4780 12164 4808
rect 7064 4768 7070 4780
rect 12158 4768 12164 4780
rect 12216 4768 12222 4820
rect 19429 4811 19487 4817
rect 19429 4777 19441 4811
rect 19475 4808 19487 4811
rect 19794 4808 19800 4820
rect 19475 4780 19800 4808
rect 19475 4777 19487 4780
rect 19429 4771 19487 4777
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 21729 4811 21787 4817
rect 21729 4777 21741 4811
rect 21775 4808 21787 4811
rect 22370 4808 22376 4820
rect 21775 4780 22376 4808
rect 21775 4777 21787 4780
rect 21729 4771 21787 4777
rect 22370 4768 22376 4780
rect 22428 4768 22434 4820
rect 22554 4768 22560 4820
rect 22612 4768 22618 4820
rect 23109 4811 23167 4817
rect 23109 4777 23121 4811
rect 23155 4777 23167 4811
rect 23109 4771 23167 4777
rect 808 4712 2176 4740
rect 3145 4743 3203 4749
rect 808 4700 814 4712
rect 3145 4709 3157 4743
rect 3191 4709 3203 4743
rect 3145 4703 3203 4709
rect 1946 4632 1952 4684
rect 2004 4632 2010 4684
rect 3160 4672 3188 4703
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 11606 4740 11612 4752
rect 6972 4712 11612 4740
rect 6972 4700 6978 4712
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 15562 4700 15568 4752
rect 15620 4740 15626 4752
rect 15620 4712 22140 4740
rect 15620 4700 15626 4712
rect 9766 4672 9772 4684
rect 2792 4644 3188 4672
rect 3252 4644 9772 4672
rect 1762 4496 1768 4548
rect 1820 4496 1826 4548
rect 1964 4468 1992 4632
rect 2792 4613 2820 4644
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4604 2927 4607
rect 3252 4604 3280 4644
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 10778 4632 10784 4684
rect 10836 4632 10842 4684
rect 2915 4576 3280 4604
rect 3329 4607 3387 4613
rect 2915 4573 2927 4576
rect 2869 4567 2927 4573
rect 3329 4573 3341 4607
rect 3375 4573 3387 4607
rect 3329 4567 3387 4573
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5902 4604 5908 4616
rect 4847 4576 5908 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 2038 4496 2044 4548
rect 2096 4496 2102 4548
rect 3344 4536 3372 4567
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 10796 4536 10824 4632
rect 16850 4564 16856 4616
rect 16908 4564 16914 4616
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 21542 4564 21548 4616
rect 21600 4564 21606 4616
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 22112 4613 22140 4712
rect 22186 4700 22192 4752
rect 22244 4740 22250 4752
rect 23124 4740 23152 4771
rect 23658 4768 23664 4820
rect 23716 4808 23722 4820
rect 23937 4811 23995 4817
rect 23937 4808 23949 4811
rect 23716 4780 23949 4808
rect 23716 4768 23722 4780
rect 23937 4777 23949 4780
rect 23983 4777 23995 4811
rect 23937 4771 23995 4777
rect 22244 4712 23152 4740
rect 22244 4700 22250 4712
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4573 22155 4607
rect 22097 4567 22155 4573
rect 23474 4564 23480 4616
rect 23532 4564 23538 4616
rect 3344 4508 10824 4536
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 22465 4539 22523 4545
rect 22465 4536 22477 4539
rect 13504 4508 22477 4536
rect 13504 4496 13510 4508
rect 22465 4505 22477 4508
rect 22511 4505 22523 4539
rect 22465 4499 22523 4505
rect 23014 4496 23020 4548
rect 23072 4496 23078 4548
rect 23842 4496 23848 4548
rect 23900 4496 23906 4548
rect 13722 4468 13728 4480
rect 1964 4440 13728 4468
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 17037 4471 17095 4477
rect 17037 4437 17049 4471
rect 17083 4468 17095 4471
rect 18598 4468 18604 4480
rect 17083 4440 18604 4468
rect 17083 4437 17095 4440
rect 17037 4431 17095 4437
rect 18598 4428 18604 4440
rect 18656 4428 18662 4480
rect 22005 4471 22063 4477
rect 22005 4437 22017 4471
rect 22051 4468 22063 4471
rect 22186 4468 22192 4480
rect 22051 4440 22192 4468
rect 22051 4437 22063 4440
rect 22005 4431 22063 4437
rect 22186 4428 22192 4440
rect 22244 4428 22250 4480
rect 22278 4428 22284 4480
rect 22336 4428 22342 4480
rect 23658 4428 23664 4480
rect 23716 4428 23722 4480
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 19429 4267 19487 4273
rect 19429 4233 19441 4267
rect 19475 4233 19487 4267
rect 19429 4227 19487 4233
rect 19444 4196 19472 4227
rect 21542 4224 21548 4276
rect 21600 4264 21606 4276
rect 22097 4267 22155 4273
rect 22097 4264 22109 4267
rect 21600 4236 22109 4264
rect 21600 4224 21606 4236
rect 22097 4233 22109 4236
rect 22143 4233 22155 4267
rect 22097 4227 22155 4233
rect 22278 4224 22284 4276
rect 22336 4224 22342 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 22428 4236 23612 4264
rect 22428 4224 22434 4236
rect 21634 4196 21640 4208
rect 19444 4168 21640 4196
rect 21634 4156 21640 4168
rect 21692 4156 21698 4208
rect 22296 4196 22324 4224
rect 22296 4168 22416 4196
rect 1486 4088 1492 4140
rect 1544 4088 1550 4140
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 10226 4128 10232 4140
rect 2639 4100 10232 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2332 4060 2360 4091
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 19242 4088 19248 4140
rect 19300 4088 19306 4140
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22388 4137 22416 4168
rect 22462 4156 22468 4208
rect 22520 4196 22526 4208
rect 23109 4199 23167 4205
rect 23109 4196 23121 4199
rect 22520 4168 23121 4196
rect 22520 4156 22526 4168
rect 23109 4165 23121 4168
rect 23155 4165 23167 4199
rect 23109 4159 23167 4165
rect 22281 4131 22339 4137
rect 22281 4128 22293 4131
rect 22244 4100 22293 4128
rect 22244 4088 22250 4100
rect 22281 4097 22293 4100
rect 22327 4097 22339 4131
rect 22281 4091 22339 4097
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 22649 4131 22707 4137
rect 22649 4097 22661 4131
rect 22695 4097 22707 4131
rect 23584 4128 23612 4236
rect 23658 4224 23664 4276
rect 23716 4224 23722 4276
rect 23676 4196 23704 4224
rect 23676 4168 24348 4196
rect 23661 4131 23719 4137
rect 23661 4128 23673 4131
rect 23584 4100 23673 4128
rect 22649 4091 22707 4097
rect 23661 4097 23673 4100
rect 23707 4097 23719 4131
rect 24210 4128 24216 4140
rect 23661 4091 23719 4097
rect 23768 4100 24216 4128
rect 4982 4060 4988 4072
rect 2332 4032 4988 4060
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 18598 4020 18604 4072
rect 18656 4060 18662 4072
rect 22664 4060 22692 4091
rect 18656 4032 22692 4060
rect 23385 4063 23443 4069
rect 18656 4020 18662 4032
rect 23385 4029 23397 4063
rect 23431 4060 23443 4063
rect 23768 4060 23796 4100
rect 24210 4088 24216 4100
rect 24268 4088 24274 4140
rect 24320 4137 24348 4168
rect 24305 4131 24363 4137
rect 24305 4097 24317 4131
rect 24351 4097 24363 4131
rect 24305 4091 24363 4097
rect 24578 4088 24584 4140
rect 24636 4088 24642 4140
rect 23431 4032 23796 4060
rect 23937 4063 23995 4069
rect 23431 4029 23443 4032
rect 23385 4023 23443 4029
rect 23937 4029 23949 4063
rect 23983 4060 23995 4063
rect 24596 4060 24624 4088
rect 23983 4032 24624 4060
rect 23983 4029 23995 4032
rect 23937 4023 23995 4029
rect 1854 3952 1860 4004
rect 1912 3992 1918 4004
rect 2409 3995 2467 4001
rect 2409 3992 2421 3995
rect 1912 3964 2421 3992
rect 1912 3952 1918 3964
rect 2409 3961 2421 3964
rect 2455 3961 2467 3995
rect 2409 3955 2467 3961
rect 20257 3995 20315 4001
rect 20257 3961 20269 3995
rect 20303 3992 20315 3995
rect 20990 3992 20996 4004
rect 20303 3964 20996 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 20990 3952 20996 3964
rect 21048 3952 21054 4004
rect 1026 3884 1032 3936
rect 1084 3924 1090 3936
rect 1581 3927 1639 3933
rect 1581 3924 1593 3927
rect 1084 3896 1593 3924
rect 1084 3884 1090 3896
rect 1581 3893 1593 3896
rect 1627 3893 1639 3927
rect 1581 3887 1639 3893
rect 2130 3884 2136 3936
rect 2188 3884 2194 3936
rect 22554 3884 22560 3936
rect 22612 3884 22618 3936
rect 22830 3884 22836 3936
rect 22888 3884 22894 3936
rect 24118 3884 24124 3936
rect 24176 3884 24182 3936
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 1486 3680 1492 3732
rect 1544 3680 1550 3732
rect 1854 3680 1860 3732
rect 1912 3680 1918 3732
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2038 3720 2044 3732
rect 1995 3692 2044 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2038 3680 2044 3692
rect 2096 3680 2102 3732
rect 2130 3680 2136 3732
rect 2188 3680 2194 3732
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 19242 3720 19248 3732
rect 18831 3692 19248 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19613 3723 19671 3729
rect 19613 3689 19625 3723
rect 19659 3720 19671 3723
rect 20070 3720 20076 3732
rect 19659 3692 20076 3720
rect 19659 3689 19671 3692
rect 19613 3683 19671 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 22554 3680 22560 3732
rect 22612 3680 22618 3732
rect 22830 3680 22836 3732
rect 22888 3680 22894 3732
rect 23293 3723 23351 3729
rect 23293 3689 23305 3723
rect 23339 3720 23351 3723
rect 23842 3720 23848 3732
rect 23339 3692 23848 3720
rect 23339 3689 23351 3692
rect 23293 3683 23351 3689
rect 23842 3680 23848 3692
rect 23900 3680 23906 3732
rect 24121 3723 24179 3729
rect 24121 3689 24133 3723
rect 24167 3720 24179 3723
rect 25314 3720 25320 3732
rect 24167 3692 25320 3720
rect 24167 3689 24179 3692
rect 24121 3683 24179 3689
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 1872 3584 1900 3680
rect 1688 3556 1900 3584
rect 1688 3525 1716 3556
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 2148 3516 2176 3680
rect 1811 3488 2176 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 18598 3476 18604 3528
rect 18656 3476 18662 3528
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 21450 3476 21456 3528
rect 21508 3476 21514 3528
rect 22572 3516 22600 3680
rect 22741 3519 22799 3525
rect 22741 3516 22753 3519
rect 22572 3488 22753 3516
rect 22741 3485 22753 3488
rect 22787 3485 22799 3519
rect 22848 3516 22876 3680
rect 22925 3655 22983 3661
rect 22925 3621 22937 3655
rect 22971 3652 22983 3655
rect 23750 3652 23756 3664
rect 22971 3624 23756 3652
rect 22971 3621 22983 3624
rect 22925 3615 22983 3621
rect 23750 3612 23756 3624
rect 23808 3612 23814 3664
rect 23109 3519 23167 3525
rect 23109 3516 23121 3519
rect 22848 3488 23121 3516
rect 22741 3479 22799 3485
rect 23109 3485 23121 3488
rect 23155 3485 23167 3519
rect 23109 3479 23167 3485
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 21468 3380 21496 3476
rect 23842 3408 23848 3460
rect 23900 3408 23906 3460
rect 23477 3383 23535 3389
rect 23477 3380 23489 3383
rect 21468 3352 23489 3380
rect 23477 3349 23489 3352
rect 23523 3349 23535 3383
rect 23477 3343 23535 3349
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18598 3176 18604 3188
rect 18279 3148 18604 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19061 3179 19119 3185
rect 19061 3145 19073 3179
rect 19107 3176 19119 3179
rect 19426 3176 19432 3188
rect 19107 3148 19432 3176
rect 19107 3145 19119 3148
rect 19061 3139 19119 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 23658 3136 23664 3188
rect 23716 3136 23722 3188
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 3602 3000 3608 3052
rect 3660 3040 3666 3052
rect 3660 3012 6914 3040
rect 3660 3000 3666 3012
rect 6886 2972 6914 3012
rect 18046 3000 18052 3052
rect 18104 3000 18110 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 18892 2972 18920 3003
rect 6886 2944 18920 2972
rect 22922 2932 22928 2984
rect 22980 2932 22986 2984
rect 22940 2836 22968 2932
rect 23676 2904 23704 3136
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3040 24087 3043
rect 24136 3040 24164 3136
rect 24075 3012 24164 3040
rect 24075 3009 24087 3012
rect 24029 3003 24087 3009
rect 24302 3000 24308 3052
rect 24360 3000 24366 3052
rect 24121 2907 24179 2913
rect 24121 2904 24133 2907
rect 23676 2876 24133 2904
rect 24121 2873 24133 2876
rect 24167 2873 24179 2907
rect 24121 2867 24179 2873
rect 23845 2839 23903 2845
rect 23845 2836 23857 2839
rect 22940 2808 23857 2836
rect 23845 2805 23857 2808
rect 23891 2805 23903 2839
rect 23845 2799 23903 2805
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 11882 2592 11888 2644
rect 11940 2632 11946 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11940 2604 11989 2632
rect 11940 2592 11946 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 11977 2595 12035 2601
rect 13446 2592 13452 2644
rect 13504 2592 13510 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20806 2632 20812 2644
rect 20027 2604 20812 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 23842 2592 23848 2644
rect 23900 2632 23906 2644
rect 24029 2635 24087 2641
rect 24029 2632 24041 2635
rect 23900 2604 24041 2632
rect 23900 2592 23906 2604
rect 24029 2601 24041 2604
rect 24075 2601 24087 2635
rect 24029 2595 24087 2601
rect 8570 2524 8576 2576
rect 8628 2524 8634 2576
rect 15657 2567 15715 2573
rect 15657 2533 15669 2567
rect 15703 2564 15715 2567
rect 23934 2564 23940 2576
rect 15703 2536 23940 2564
rect 15703 2533 15715 2536
rect 15657 2527 15715 2533
rect 23934 2524 23940 2536
rect 23992 2524 23998 2576
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6788 2400 7113 2428
rect 6788 2388 6794 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 10778 2388 10784 2440
rect 10836 2388 10842 2440
rect 11790 2388 11796 2440
rect 11848 2388 11854 2440
rect 12158 2388 12164 2440
rect 12216 2388 12222 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 14366 2388 14372 2440
rect 14424 2388 14430 2440
rect 15470 2388 15476 2440
rect 15528 2388 15534 2440
rect 19794 2388 19800 2440
rect 19852 2388 19858 2440
rect 24210 2388 24216 2440
rect 24268 2388 24274 2440
rect 24026 2360 24032 2372
rect 9784 2332 24032 2360
rect 7282 2252 7288 2304
rect 7340 2252 7346 2304
rect 9784 2301 9812 2332
rect 24026 2320 24032 2332
rect 24084 2320 24090 2372
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10962 2252 10968 2304
rect 11020 2252 11026 2304
rect 12342 2252 12348 2304
rect 12400 2252 12406 2304
rect 14550 2252 14556 2304
rect 14608 2252 14614 2304
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 6730 2048 6736 2100
rect 6788 2048 6794 2100
rect 8021 2091 8079 2097
rect 8021 2057 8033 2091
rect 8067 2088 8079 2091
rect 8386 2088 8392 2100
rect 8067 2060 8392 2088
rect 8067 2057 8079 2060
rect 8021 2051 8079 2057
rect 8386 2048 8392 2060
rect 8444 2048 8450 2100
rect 9217 2091 9275 2097
rect 9217 2057 9229 2091
rect 9263 2088 9275 2091
rect 9582 2088 9588 2100
rect 9263 2060 9588 2088
rect 9263 2057 9275 2060
rect 9217 2051 9275 2057
rect 9582 2048 9588 2060
rect 9640 2048 9646 2100
rect 10413 2091 10471 2097
rect 10413 2057 10425 2091
rect 10459 2088 10471 2091
rect 10778 2088 10784 2100
rect 10459 2060 10784 2088
rect 10459 2057 10471 2060
rect 10413 2051 10471 2057
rect 10778 2048 10784 2060
rect 10836 2048 10842 2100
rect 11701 2091 11759 2097
rect 11701 2057 11713 2091
rect 11747 2057 11759 2091
rect 11701 2051 11759 2057
rect 11716 2020 11744 2051
rect 11790 2048 11796 2100
rect 11848 2088 11854 2100
rect 11977 2091 12035 2097
rect 11977 2088 11989 2091
rect 11848 2060 11989 2088
rect 11848 2048 11854 2060
rect 11977 2057 11989 2060
rect 12023 2057 12035 2091
rect 11977 2051 12035 2057
rect 12158 2048 12164 2100
rect 12216 2048 12222 2100
rect 12805 2091 12863 2097
rect 12805 2057 12817 2091
rect 12851 2088 12863 2091
rect 13262 2088 13268 2100
rect 12851 2060 13268 2088
rect 12851 2057 12863 2060
rect 12805 2051 12863 2057
rect 13262 2048 13268 2060
rect 13320 2048 13326 2100
rect 14001 2091 14059 2097
rect 14001 2057 14013 2091
rect 14047 2088 14059 2091
rect 14366 2088 14372 2100
rect 14047 2060 14372 2088
rect 14047 2057 14059 2060
rect 14001 2051 14059 2057
rect 14366 2048 14372 2060
rect 14424 2048 14430 2100
rect 15105 2091 15163 2097
rect 15105 2057 15117 2091
rect 15151 2088 15163 2091
rect 15470 2088 15476 2100
rect 15151 2060 15476 2088
rect 15151 2057 15163 2060
rect 15105 2051 15163 2057
rect 15470 2048 15476 2060
rect 15528 2048 15534 2100
rect 18785 2091 18843 2097
rect 18785 2057 18797 2091
rect 18831 2057 18843 2091
rect 18785 2051 18843 2057
rect 19429 2091 19487 2097
rect 19429 2057 19441 2091
rect 19475 2088 19487 2091
rect 19794 2088 19800 2100
rect 19475 2060 19800 2088
rect 19475 2057 19487 2060
rect 19429 2051 19487 2057
rect 12176 2020 12204 2048
rect 11716 1992 12204 2020
rect 6546 1912 6552 1964
rect 6604 1912 6610 1964
rect 7834 1912 7840 1964
rect 7892 1912 7898 1964
rect 9030 1912 9036 1964
rect 9088 1912 9094 1964
rect 10226 1912 10232 1964
rect 10284 1912 10290 1964
rect 11514 1912 11520 1964
rect 11572 1912 11578 1964
rect 11606 1912 11612 1964
rect 11664 1952 11670 1964
rect 11793 1955 11851 1961
rect 11793 1952 11805 1955
rect 11664 1924 11805 1952
rect 11664 1912 11670 1924
rect 11793 1921 11805 1924
rect 11839 1921 11851 1955
rect 11793 1915 11851 1921
rect 12618 1912 12624 1964
rect 12676 1912 12682 1964
rect 13814 1912 13820 1964
rect 13872 1912 13878 1964
rect 14918 1912 14924 1964
rect 14976 1912 14982 1964
rect 18601 1955 18659 1961
rect 18601 1952 18613 1955
rect 16546 1924 18613 1952
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 16546 1884 16574 1924
rect 18601 1921 18613 1924
rect 18647 1921 18659 1955
rect 18800 1952 18828 2051
rect 19794 2048 19800 2060
rect 19852 2048 19858 2100
rect 24210 2048 24216 2100
rect 24268 2088 24274 2100
rect 24305 2091 24363 2097
rect 24305 2088 24317 2091
rect 24268 2060 24317 2088
rect 24268 2048 24274 2060
rect 24305 2057 24317 2060
rect 24351 2057 24363 2091
rect 24305 2051 24363 2057
rect 19245 1955 19303 1961
rect 19245 1952 19257 1955
rect 18800 1924 19257 1952
rect 18601 1915 18659 1921
rect 19245 1921 19257 1924
rect 19291 1921 19303 1955
rect 19245 1915 19303 1921
rect 24118 1912 24124 1964
rect 24176 1912 24182 1964
rect 2464 1856 16574 1884
rect 2464 1844 2470 1856
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 2406 1504 2412 1556
rect 2464 1504 2470 1556
rect 6546 1504 6552 1556
rect 6604 1504 6610 1556
rect 7469 1547 7527 1553
rect 7469 1513 7481 1547
rect 7515 1544 7527 1547
rect 7834 1544 7840 1556
rect 7515 1516 7840 1544
rect 7515 1513 7527 1516
rect 7469 1507 7527 1513
rect 7834 1504 7840 1516
rect 7892 1504 7898 1556
rect 8665 1547 8723 1553
rect 8665 1513 8677 1547
rect 8711 1544 8723 1547
rect 9030 1544 9036 1556
rect 8711 1516 9036 1544
rect 8711 1513 8723 1516
rect 8665 1507 8723 1513
rect 9030 1504 9036 1516
rect 9088 1504 9094 1556
rect 9861 1547 9919 1553
rect 9861 1513 9873 1547
rect 9907 1544 9919 1547
rect 10226 1544 10232 1556
rect 9907 1516 10232 1544
rect 9907 1513 9919 1516
rect 9861 1507 9919 1513
rect 10226 1504 10232 1516
rect 10284 1504 10290 1556
rect 11149 1547 11207 1553
rect 11149 1513 11161 1547
rect 11195 1544 11207 1547
rect 11514 1544 11520 1556
rect 11195 1516 11520 1544
rect 11195 1513 11207 1516
rect 11149 1507 11207 1513
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 12253 1547 12311 1553
rect 12253 1513 12265 1547
rect 12299 1544 12311 1547
rect 12618 1544 12624 1556
rect 12299 1516 12624 1544
rect 12299 1513 12311 1516
rect 12253 1507 12311 1513
rect 12618 1504 12624 1516
rect 12676 1504 12682 1556
rect 14645 1547 14703 1553
rect 14645 1513 14657 1547
rect 14691 1544 14703 1547
rect 14918 1544 14924 1556
rect 14691 1516 14924 1544
rect 14691 1513 14703 1516
rect 14645 1507 14703 1513
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
rect 23477 1547 23535 1553
rect 23477 1513 23489 1547
rect 23523 1544 23535 1547
rect 24118 1544 24124 1556
rect 23523 1516 24124 1544
rect 23523 1513 23535 1516
rect 23477 1507 23535 1513
rect 24118 1504 24124 1516
rect 24176 1504 24182 1556
rect 5997 1479 6055 1485
rect 5997 1445 6009 1479
rect 6043 1445 6055 1479
rect 5997 1439 6055 1445
rect 7193 1479 7251 1485
rect 7193 1445 7205 1479
rect 7239 1445 7251 1479
rect 7193 1439 7251 1445
rect 934 1300 940 1352
rect 992 1340 998 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 992 1312 1409 1340
rect 992 1300 998 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 2222 1300 2228 1352
rect 2280 1300 2286 1352
rect 3418 1300 3424 1352
rect 3476 1300 3482 1352
rect 4614 1300 4620 1352
rect 4672 1300 4678 1352
rect 5810 1300 5816 1352
rect 5868 1300 5874 1352
rect 6012 1340 6040 1439
rect 6365 1343 6423 1349
rect 6365 1340 6377 1343
rect 6012 1312 6377 1340
rect 6365 1309 6377 1312
rect 6411 1309 6423 1343
rect 6365 1303 6423 1309
rect 7006 1300 7012 1352
rect 7064 1300 7070 1352
rect 7208 1340 7236 1439
rect 7285 1343 7343 1349
rect 7285 1340 7297 1343
rect 7208 1312 7297 1340
rect 7285 1309 7297 1312
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 8404 1312 8493 1340
rect 1596 1244 8340 1272
rect 1596 1213 1624 1244
rect 8312 1216 8340 1244
rect 1581 1207 1639 1213
rect 1581 1173 1593 1207
rect 1627 1173 1639 1207
rect 1581 1167 1639 1173
rect 3602 1164 3608 1216
rect 3660 1164 3666 1216
rect 4798 1164 4804 1216
rect 4856 1164 4862 1216
rect 8294 1164 8300 1216
rect 8352 1164 8358 1216
rect 8404 1213 8432 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8481 1303 8539 1309
rect 9398 1300 9404 1352
rect 9456 1300 9462 1352
rect 9677 1343 9735 1349
rect 9677 1340 9689 1343
rect 9600 1312 9689 1340
rect 9600 1213 9628 1312
rect 9677 1309 9689 1312
rect 9723 1309 9735 1343
rect 9677 1303 9735 1309
rect 10410 1300 10416 1352
rect 10468 1300 10474 1352
rect 10686 1300 10692 1352
rect 10744 1300 10750 1352
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 10980 1272 11008 1303
rect 11606 1300 11612 1352
rect 11664 1300 11670 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 12069 1343 12127 1349
rect 12069 1340 12081 1343
rect 11992 1312 12081 1340
rect 10612 1244 11008 1272
rect 10612 1213 10640 1244
rect 8389 1207 8447 1213
rect 8389 1173 8401 1207
rect 8435 1173 8447 1207
rect 8389 1167 8447 1173
rect 9585 1207 9643 1213
rect 9585 1173 9597 1207
rect 9631 1173 9643 1207
rect 9585 1167 9643 1173
rect 10597 1207 10655 1213
rect 10597 1173 10609 1207
rect 10643 1173 10655 1207
rect 10597 1167 10655 1173
rect 10873 1207 10931 1213
rect 10873 1173 10885 1207
rect 10919 1204 10931 1207
rect 11624 1204 11652 1300
rect 11992 1213 12020 1312
rect 12069 1309 12081 1312
rect 12115 1309 12127 1343
rect 12069 1303 12127 1309
rect 12710 1300 12716 1352
rect 12768 1340 12774 1352
rect 12989 1343 13047 1349
rect 12989 1340 13001 1343
rect 12768 1312 13001 1340
rect 12768 1300 12774 1312
rect 12989 1309 13001 1312
rect 13035 1309 13047 1343
rect 13265 1343 13323 1349
rect 13265 1340 13277 1343
rect 12989 1303 13047 1309
rect 13188 1312 13277 1340
rect 13188 1213 13216 1312
rect 13265 1309 13277 1312
rect 13311 1309 13323 1343
rect 13265 1303 13323 1309
rect 13814 1300 13820 1352
rect 13872 1300 13878 1352
rect 14182 1300 14188 1352
rect 14240 1300 14246 1352
rect 14461 1343 14519 1349
rect 14461 1340 14473 1343
rect 14384 1312 14473 1340
rect 10919 1176 11652 1204
rect 11977 1207 12035 1213
rect 10919 1173 10931 1176
rect 10873 1167 10931 1173
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 13173 1207 13231 1213
rect 13173 1173 13185 1207
rect 13219 1173 13231 1207
rect 13173 1167 13231 1173
rect 13449 1207 13507 1213
rect 13449 1173 13461 1207
rect 13495 1204 13507 1207
rect 13832 1204 13860 1300
rect 14384 1213 14412 1312
rect 14461 1309 14473 1312
rect 14507 1309 14519 1343
rect 14461 1303 14519 1309
rect 15378 1300 15384 1352
rect 15436 1300 15442 1352
rect 15562 1300 15568 1352
rect 15620 1300 15626 1352
rect 16666 1300 16672 1352
rect 16724 1300 16730 1352
rect 16850 1300 16856 1352
rect 16908 1300 16914 1352
rect 17770 1300 17776 1352
rect 17828 1300 17834 1352
rect 18046 1300 18052 1352
rect 18104 1300 18110 1352
rect 18138 1300 18144 1352
rect 18196 1340 18202 1352
rect 18693 1343 18751 1349
rect 18693 1340 18705 1343
rect 18196 1312 18705 1340
rect 18196 1300 18202 1312
rect 18693 1309 18705 1312
rect 18739 1309 18751 1343
rect 18693 1303 18751 1309
rect 19150 1300 19156 1352
rect 19208 1300 19214 1352
rect 19242 1300 19248 1352
rect 19300 1300 19306 1352
rect 20162 1300 20168 1352
rect 20220 1300 20226 1352
rect 20714 1300 20720 1352
rect 20772 1300 20778 1352
rect 21358 1300 21364 1352
rect 21416 1300 21422 1352
rect 21634 1300 21640 1352
rect 21692 1300 21698 1352
rect 22554 1300 22560 1352
rect 22612 1300 22618 1352
rect 23293 1343 23351 1349
rect 23293 1309 23305 1343
rect 23339 1340 23351 1343
rect 23339 1312 23796 1340
rect 23339 1309 23351 1312
rect 23293 1303 23351 1309
rect 15580 1213 15608 1300
rect 16868 1213 16896 1300
rect 13495 1176 13860 1204
rect 14369 1207 14427 1213
rect 13495 1173 13507 1176
rect 13449 1167 13507 1173
rect 14369 1173 14381 1207
rect 14415 1173 14427 1207
rect 14369 1167 14427 1173
rect 15565 1207 15623 1213
rect 15565 1173 15577 1207
rect 15611 1173 15623 1207
rect 15565 1167 15623 1173
rect 16853 1207 16911 1213
rect 16853 1173 16865 1207
rect 16899 1173 16911 1207
rect 16853 1167 16911 1173
rect 17957 1207 18015 1213
rect 17957 1173 17969 1207
rect 18003 1204 18015 1207
rect 18064 1204 18092 1300
rect 18506 1232 18512 1284
rect 18564 1232 18570 1284
rect 18003 1176 18092 1204
rect 18524 1204 18552 1232
rect 18877 1207 18935 1213
rect 18877 1204 18889 1207
rect 18524 1176 18889 1204
rect 18003 1173 18015 1176
rect 17957 1167 18015 1173
rect 18877 1173 18889 1176
rect 18923 1173 18935 1207
rect 19168 1204 19196 1300
rect 19429 1207 19487 1213
rect 19429 1204 19441 1207
rect 19168 1176 19441 1204
rect 18877 1167 18935 1173
rect 19429 1173 19441 1176
rect 19475 1173 19487 1207
rect 19429 1167 19487 1173
rect 20349 1207 20407 1213
rect 20349 1173 20361 1207
rect 20395 1204 20407 1207
rect 20732 1204 20760 1300
rect 20395 1176 20760 1204
rect 21545 1207 21603 1213
rect 20395 1173 20407 1176
rect 20349 1167 20407 1173
rect 21545 1173 21557 1207
rect 21591 1204 21603 1207
rect 21652 1204 21680 1300
rect 23474 1232 23480 1284
rect 23532 1232 23538 1284
rect 21591 1176 21680 1204
rect 22741 1207 22799 1213
rect 21591 1173 21603 1176
rect 21545 1167 21603 1173
rect 22741 1173 22753 1207
rect 22787 1204 22799 1207
rect 23492 1204 23520 1232
rect 23768 1213 23796 1312
rect 23934 1300 23940 1352
rect 23992 1300 23998 1352
rect 24029 1343 24087 1349
rect 24029 1309 24041 1343
rect 24075 1340 24087 1343
rect 24486 1340 24492 1352
rect 24075 1312 24492 1340
rect 24075 1309 24087 1312
rect 24029 1303 24087 1309
rect 24486 1300 24492 1312
rect 24544 1300 24550 1352
rect 24302 1232 24308 1284
rect 24360 1232 24366 1284
rect 22787 1176 23520 1204
rect 23753 1207 23811 1213
rect 22787 1173 22799 1176
rect 22741 1167 22799 1173
rect 23753 1173 23765 1207
rect 23799 1173 23811 1207
rect 23753 1167 23811 1173
rect 24213 1207 24271 1213
rect 24213 1173 24225 1207
rect 24259 1204 24271 1207
rect 24320 1204 24348 1232
rect 24259 1176 24348 1204
rect 24259 1173 24271 1176
rect 24213 1167 24271 1173
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 4798 960 4804 1012
rect 4856 1000 4862 1012
rect 10686 1000 10692 1012
rect 4856 972 10692 1000
rect 4856 960 4862 972
rect 10686 960 10692 972
rect 10744 960 10750 1012
rect 18138 1000 18144 1012
rect 16546 972 18144 1000
rect 8294 892 8300 944
rect 8352 932 8358 944
rect 16546 932 16574 972
rect 18138 960 18144 972
rect 18196 960 18202 1012
rect 8352 904 16574 932
rect 8352 892 8358 904
<< via1 >>
rect 9128 7896 9180 7948
rect 19432 7896 19484 7948
rect 8024 7828 8076 7880
rect 19340 7828 19392 7880
rect 7748 7760 7800 7812
rect 17960 7760 18012 7812
rect 21916 7760 21968 7812
rect 23480 7760 23532 7812
rect 18236 7692 18288 7744
rect 8760 7624 8812 7676
rect 17408 7624 17460 7676
rect 7656 7556 7708 7608
rect 8116 7556 8168 7608
rect 11152 7556 11204 7608
rect 10784 7488 10836 7540
rect 5908 7420 5960 7472
rect 11060 7420 11112 7472
rect 11888 7420 11940 7472
rect 21548 7420 21600 7472
rect 4712 7352 4764 7404
rect 4988 7352 5040 7404
rect 8668 7352 8720 7404
rect 2872 7284 2924 7336
rect 10876 7284 10928 7336
rect 11704 7284 11756 7336
rect 12348 7284 12400 7336
rect 12256 7216 12308 7268
rect 4528 7148 4580 7200
rect 8116 7148 8168 7200
rect 9680 7148 9732 7200
rect 4804 7080 4856 7132
rect 12624 7148 12676 7200
rect 17684 7148 17736 7200
rect 18420 7148 18472 7200
rect 8300 7012 8352 7064
rect 17500 7080 17552 7132
rect 8116 6944 8168 6996
rect 12348 6944 12400 6996
rect 14096 6944 14148 6996
rect 20536 7012 20588 7064
rect 3424 6876 3476 6928
rect 9680 6876 9732 6928
rect 9772 6876 9824 6928
rect 16948 6876 17000 6928
rect 4252 6808 4304 6860
rect 9220 6808 9272 6860
rect 9496 6808 9548 6860
rect 14740 6808 14792 6860
rect 14832 6808 14884 6860
rect 15752 6808 15804 6860
rect 15936 6808 15988 6860
rect 16396 6808 16448 6860
rect 16764 6808 16816 6860
rect 18052 6808 18104 6860
rect 6184 6740 6236 6792
rect 14096 6740 14148 6792
rect 8392 6604 8444 6656
rect 19616 6740 19668 6792
rect 18144 6672 18196 6724
rect 19708 6672 19760 6724
rect 17040 6604 17092 6656
rect 18328 6604 18380 6656
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 2964 6400 3016 6452
rect 4068 6400 4120 6452
rect 4252 6400 4304 6452
rect 480 6332 532 6384
rect 2872 6332 2924 6384
rect 5264 6400 5316 6452
rect 5724 6400 5776 6452
rect 2228 6264 2280 6316
rect 5172 6332 5224 6384
rect 6184 6400 6236 6452
rect 6276 6400 6328 6452
rect 7380 6400 7432 6452
rect 7564 6443 7616 6452
rect 7564 6409 7573 6443
rect 7573 6409 7607 6443
rect 7607 6409 7616 6443
rect 7564 6400 7616 6409
rect 8484 6400 8536 6452
rect 8576 6443 8628 6452
rect 8576 6409 8585 6443
rect 8585 6409 8619 6443
rect 8619 6409 8628 6443
rect 8576 6400 8628 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 3332 6196 3384 6248
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 5816 6264 5868 6316
rect 7472 6332 7524 6384
rect 8300 6332 8352 6384
rect 8392 6332 8444 6384
rect 9772 6400 9824 6452
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 9588 6332 9640 6384
rect 10876 6443 10928 6452
rect 10876 6409 10885 6443
rect 10885 6409 10919 6443
rect 10919 6409 10928 6443
rect 10876 6400 10928 6409
rect 11060 6400 11112 6452
rect 7104 6264 7156 6316
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 7564 6264 7616 6316
rect 8024 6264 8076 6316
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 10232 6264 10284 6316
rect 10508 6264 10560 6316
rect 4344 6060 4396 6112
rect 6736 6060 6788 6112
rect 9588 6128 9640 6180
rect 11060 6128 11112 6180
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12440 6332 12492 6384
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 12808 6400 12860 6452
rect 12992 6400 13044 6452
rect 14188 6332 14240 6384
rect 15108 6400 15160 6452
rect 12624 6264 12676 6316
rect 12808 6311 12860 6316
rect 12808 6277 12825 6311
rect 12825 6277 12859 6311
rect 12859 6277 12860 6311
rect 12808 6264 12860 6277
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 12532 6196 12584 6248
rect 12716 6196 12768 6248
rect 11336 6128 11388 6180
rect 11704 6060 11756 6112
rect 11980 6103 12032 6112
rect 11980 6069 11989 6103
rect 11989 6069 12023 6103
rect 12023 6069 12032 6103
rect 11980 6060 12032 6069
rect 12164 6060 12216 6112
rect 12532 6103 12584 6112
rect 12532 6069 12541 6103
rect 12541 6069 12575 6103
rect 12575 6069 12584 6103
rect 12532 6060 12584 6069
rect 12808 6060 12860 6112
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 13728 6060 13780 6069
rect 14372 6103 14424 6112
rect 14372 6069 14381 6103
rect 14381 6069 14415 6103
rect 14415 6069 14424 6103
rect 14372 6060 14424 6069
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15200 6060 15252 6069
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 15752 6264 15804 6316
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17316 6400 17368 6452
rect 16120 6128 16172 6180
rect 16672 6171 16724 6180
rect 16672 6137 16681 6171
rect 16681 6137 16715 6171
rect 16715 6137 16724 6171
rect 16672 6128 16724 6137
rect 17500 6171 17552 6180
rect 17500 6137 17509 6171
rect 17509 6137 17543 6171
rect 17543 6137 17552 6171
rect 17500 6128 17552 6137
rect 18420 6332 18472 6384
rect 18052 6264 18104 6316
rect 18328 6264 18380 6316
rect 19340 6400 19392 6452
rect 20076 6400 20128 6452
rect 20444 6400 20496 6452
rect 21272 6400 21324 6452
rect 18972 6332 19024 6384
rect 19524 6332 19576 6384
rect 21088 6332 21140 6384
rect 21364 6332 21416 6384
rect 23480 6400 23532 6452
rect 19708 6307 19760 6316
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 19892 6264 19944 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20812 6307 20864 6316
rect 20812 6273 20821 6307
rect 20821 6273 20855 6307
rect 20855 6273 20864 6307
rect 20812 6264 20864 6273
rect 21456 6307 21508 6316
rect 21456 6273 21465 6307
rect 21465 6273 21499 6307
rect 21499 6273 21508 6307
rect 21456 6264 21508 6273
rect 21548 6264 21600 6316
rect 22468 6307 22520 6316
rect 22468 6273 22477 6307
rect 22477 6273 22511 6307
rect 22511 6273 22520 6307
rect 22468 6264 22520 6273
rect 23020 6307 23072 6316
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 24032 6264 24084 6316
rect 18420 6128 18472 6180
rect 18604 6103 18656 6112
rect 18604 6069 18613 6103
rect 18613 6069 18647 6103
rect 18647 6069 18656 6103
rect 18604 6060 18656 6069
rect 18880 6103 18932 6112
rect 18880 6069 18889 6103
rect 18889 6069 18923 6103
rect 18923 6069 18932 6103
rect 18880 6060 18932 6069
rect 19616 6060 19668 6112
rect 21640 6103 21692 6112
rect 21640 6069 21649 6103
rect 21649 6069 21683 6103
rect 21683 6069 21692 6103
rect 21640 6060 21692 6069
rect 21824 6060 21876 6112
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 2136 5856 2188 5908
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 2688 5899 2740 5908
rect 2688 5865 2697 5899
rect 2697 5865 2731 5899
rect 2731 5865 2740 5899
rect 2688 5856 2740 5865
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3792 5856 3844 5908
rect 4436 5856 4488 5908
rect 4804 5856 4856 5908
rect 4896 5899 4948 5908
rect 4896 5865 4905 5899
rect 4905 5865 4939 5899
rect 4939 5865 4948 5899
rect 4896 5856 4948 5865
rect 6000 5899 6052 5908
rect 6000 5865 6009 5899
rect 6009 5865 6043 5899
rect 6043 5865 6052 5899
rect 6000 5856 6052 5865
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7380 5856 7432 5908
rect 7932 5899 7984 5908
rect 7932 5865 7941 5899
rect 7941 5865 7975 5899
rect 7975 5865 7984 5899
rect 7932 5856 7984 5865
rect 8116 5856 8168 5908
rect 8208 5856 8260 5908
rect 8668 5856 8720 5908
rect 9036 5856 9088 5908
rect 9220 5856 9272 5908
rect 12256 5856 12308 5908
rect 13084 5856 13136 5908
rect 14740 5856 14792 5908
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 7196 5831 7248 5840
rect 7196 5797 7205 5831
rect 7205 5797 7239 5831
rect 7239 5797 7248 5831
rect 7196 5788 7248 5797
rect 9864 5788 9916 5840
rect 3424 5652 3476 5704
rect 4528 5652 4580 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 5172 5627 5224 5636
rect 5172 5593 5181 5627
rect 5181 5593 5215 5627
rect 5215 5593 5224 5627
rect 5172 5584 5224 5593
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 9496 5720 9548 5772
rect 10048 5788 10100 5840
rect 11060 5788 11112 5840
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 16856 5856 16908 5908
rect 17408 5856 17460 5908
rect 17776 5856 17828 5908
rect 18328 5856 18380 5908
rect 18788 5856 18840 5908
rect 18880 5856 18932 5908
rect 19340 5856 19392 5908
rect 19524 5899 19576 5908
rect 19524 5865 19533 5899
rect 19533 5865 19567 5899
rect 19567 5865 19576 5899
rect 19524 5856 19576 5865
rect 19616 5856 19668 5908
rect 6276 5627 6328 5636
rect 6276 5593 6285 5627
rect 6285 5593 6319 5627
rect 6319 5593 6328 5627
rect 6276 5584 6328 5593
rect 7380 5627 7432 5636
rect 7380 5593 7389 5627
rect 7389 5593 7423 5627
rect 7423 5593 7432 5627
rect 7380 5584 7432 5593
rect 7840 5627 7892 5636
rect 7840 5593 7849 5627
rect 7849 5593 7883 5627
rect 7883 5593 7892 5627
rect 7840 5584 7892 5593
rect 8668 5627 8720 5636
rect 8668 5593 8677 5627
rect 8677 5593 8711 5627
rect 8711 5593 8720 5627
rect 8668 5584 8720 5593
rect 9128 5584 9180 5636
rect 9956 5652 10008 5704
rect 11980 5720 12032 5772
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10876 5652 10928 5704
rect 11060 5652 11112 5704
rect 11336 5652 11388 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12532 5720 12584 5772
rect 12716 5720 12768 5772
rect 16304 5788 16356 5840
rect 13084 5652 13136 5704
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14280 5652 14332 5704
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 9864 5559 9916 5568
rect 9864 5525 9873 5559
rect 9873 5525 9907 5559
rect 9907 5525 9916 5559
rect 9864 5516 9916 5525
rect 9956 5516 10008 5568
rect 10784 5559 10836 5568
rect 10784 5525 10793 5559
rect 10793 5525 10827 5559
rect 10827 5525 10836 5559
rect 10784 5516 10836 5525
rect 11060 5559 11112 5568
rect 11060 5525 11069 5559
rect 11069 5525 11103 5559
rect 11103 5525 11112 5559
rect 11060 5516 11112 5525
rect 11612 5559 11664 5568
rect 11612 5525 11621 5559
rect 11621 5525 11655 5559
rect 11655 5525 11664 5559
rect 11612 5516 11664 5525
rect 11704 5516 11756 5568
rect 11980 5516 12032 5568
rect 15476 5584 15528 5636
rect 14004 5516 14056 5568
rect 15660 5516 15712 5568
rect 16488 5652 16540 5704
rect 16304 5584 16356 5636
rect 17316 5831 17368 5840
rect 17316 5797 17325 5831
rect 17325 5797 17359 5831
rect 17359 5797 17368 5831
rect 17316 5788 17368 5797
rect 18604 5788 18656 5840
rect 18420 5652 18472 5704
rect 18604 5695 18656 5704
rect 18604 5661 18613 5695
rect 18613 5661 18647 5695
rect 18647 5661 18656 5695
rect 18604 5652 18656 5661
rect 21640 5856 21692 5908
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 17868 5516 17920 5525
rect 17960 5516 18012 5568
rect 18328 5516 18380 5568
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 20628 5788 20680 5840
rect 21088 5652 21140 5704
rect 22284 5856 22336 5908
rect 22836 5856 22888 5908
rect 23480 5856 23532 5908
rect 25596 5856 25648 5908
rect 20904 5584 20956 5636
rect 20996 5627 21048 5636
rect 20996 5593 21005 5627
rect 21005 5593 21039 5627
rect 21039 5593 21048 5627
rect 20996 5584 21048 5593
rect 21916 5627 21968 5636
rect 21916 5593 21925 5627
rect 21925 5593 21959 5627
rect 21959 5593 21968 5627
rect 21916 5584 21968 5593
rect 22468 5627 22520 5636
rect 22468 5593 22477 5627
rect 22477 5593 22511 5627
rect 22511 5593 22520 5627
rect 22468 5584 22520 5593
rect 23020 5627 23072 5636
rect 23020 5593 23029 5627
rect 23029 5593 23063 5627
rect 23063 5593 23072 5627
rect 23020 5584 23072 5593
rect 23940 5584 23992 5636
rect 20076 5559 20128 5568
rect 20076 5525 20085 5559
rect 20085 5525 20119 5559
rect 20119 5525 20128 5559
rect 20076 5516 20128 5525
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 24032 5559 24084 5568
rect 24032 5525 24041 5559
rect 24041 5525 24075 5559
rect 24075 5525 24084 5559
rect 24032 5516 24084 5525
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 3608 5312 3660 5364
rect 1584 5244 1636 5296
rect 4344 5312 4396 5364
rect 4528 5355 4580 5364
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 296 5108 348 5160
rect 3700 5176 3752 5228
rect 4436 5176 4488 5228
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 5816 5355 5868 5364
rect 5816 5321 5825 5355
rect 5825 5321 5859 5355
rect 5859 5321 5868 5355
rect 5816 5312 5868 5321
rect 7380 5312 7432 5364
rect 7472 5312 7524 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 5264 5108 5316 5160
rect 5540 5108 5592 5160
rect 7196 5176 7248 5228
rect 7288 5176 7340 5228
rect 7656 5176 7708 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 8576 5312 8628 5364
rect 8668 5355 8720 5364
rect 8668 5321 8677 5355
rect 8677 5321 8711 5355
rect 8711 5321 8720 5355
rect 8668 5312 8720 5321
rect 9312 5312 9364 5364
rect 9864 5312 9916 5364
rect 10140 5355 10192 5364
rect 10140 5321 10149 5355
rect 10149 5321 10183 5355
rect 10183 5321 10192 5355
rect 10140 5312 10192 5321
rect 9772 5244 9824 5296
rect 6920 5108 6972 5160
rect 7012 5108 7064 5160
rect 3516 4972 3568 5024
rect 6736 4972 6788 5024
rect 9588 5176 9640 5228
rect 11060 5312 11112 5364
rect 12348 5312 12400 5364
rect 17868 5312 17920 5364
rect 18604 5312 18656 5364
rect 19248 5312 19300 5364
rect 19984 5312 20036 5364
rect 20076 5312 20128 5364
rect 21456 5312 21508 5364
rect 21916 5312 21968 5364
rect 23572 5312 23624 5364
rect 10232 5176 10284 5228
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 10508 5108 10560 5160
rect 10692 5176 10744 5228
rect 18420 5244 18472 5296
rect 11428 5176 11480 5228
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 19064 5219 19116 5228
rect 19064 5185 19073 5219
rect 19073 5185 19107 5219
rect 19107 5185 19116 5219
rect 19064 5176 19116 5185
rect 19340 5219 19392 5228
rect 19340 5185 19349 5219
rect 19349 5185 19383 5219
rect 19383 5185 19392 5219
rect 19340 5176 19392 5185
rect 19800 5219 19852 5228
rect 19800 5185 19809 5219
rect 19809 5185 19843 5219
rect 19843 5185 19852 5219
rect 19800 5176 19852 5185
rect 20168 5244 20220 5296
rect 16672 5108 16724 5160
rect 20720 5219 20772 5228
rect 20720 5185 20729 5219
rect 20729 5185 20763 5219
rect 20763 5185 20772 5219
rect 20720 5176 20772 5185
rect 24032 5244 24084 5296
rect 21456 5219 21508 5228
rect 21456 5185 21465 5219
rect 21465 5185 21499 5219
rect 21499 5185 21508 5219
rect 21456 5176 21508 5185
rect 21640 5176 21692 5228
rect 22928 5219 22980 5228
rect 22928 5185 22937 5219
rect 22937 5185 22971 5219
rect 22971 5185 22980 5219
rect 22928 5176 22980 5185
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 9680 5040 9732 5092
rect 19892 5040 19944 5092
rect 20076 5083 20128 5092
rect 20076 5049 20085 5083
rect 20085 5049 20119 5083
rect 20119 5049 20128 5083
rect 20076 5040 20128 5049
rect 25044 5108 25096 5160
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 11152 4972 11204 5024
rect 18512 4972 18564 5024
rect 20260 4972 20312 5024
rect 20904 4972 20956 5024
rect 23848 5040 23900 5092
rect 22468 4972 22520 5024
rect 24308 4972 24360 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 1308 4768 1360 4820
rect 756 4700 808 4752
rect 2228 4768 2280 4820
rect 3700 4768 3752 4820
rect 4436 4768 4488 4820
rect 5264 4768 5316 4820
rect 6736 4768 6788 4820
rect 7012 4768 7064 4820
rect 12164 4768 12216 4820
rect 19800 4768 19852 4820
rect 22376 4768 22428 4820
rect 22560 4811 22612 4820
rect 22560 4777 22569 4811
rect 22569 4777 22603 4811
rect 22603 4777 22612 4811
rect 22560 4768 22612 4777
rect 1952 4632 2004 4684
rect 6920 4700 6972 4752
rect 11612 4700 11664 4752
rect 15568 4700 15620 4752
rect 1768 4539 1820 4548
rect 1768 4505 1777 4539
rect 1777 4505 1811 4539
rect 1811 4505 1820 4539
rect 1768 4496 1820 4505
rect 9772 4632 9824 4684
rect 10784 4632 10836 4684
rect 2044 4539 2096 4548
rect 2044 4505 2053 4539
rect 2053 4505 2087 4539
rect 2087 4505 2096 4539
rect 2044 4496 2096 4505
rect 5908 4564 5960 4616
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 22192 4700 22244 4752
rect 23664 4768 23716 4820
rect 23480 4607 23532 4616
rect 23480 4573 23489 4607
rect 23489 4573 23523 4607
rect 23523 4573 23532 4607
rect 23480 4564 23532 4573
rect 13452 4496 13504 4548
rect 23020 4539 23072 4548
rect 23020 4505 23029 4539
rect 23029 4505 23063 4539
rect 23063 4505 23072 4539
rect 23020 4496 23072 4505
rect 23848 4539 23900 4548
rect 23848 4505 23857 4539
rect 23857 4505 23891 4539
rect 23891 4505 23900 4539
rect 23848 4496 23900 4505
rect 13728 4428 13780 4480
rect 18604 4428 18656 4480
rect 22192 4428 22244 4480
rect 22284 4471 22336 4480
rect 22284 4437 22293 4471
rect 22293 4437 22327 4471
rect 22327 4437 22336 4471
rect 22284 4428 22336 4437
rect 23664 4471 23716 4480
rect 23664 4437 23673 4471
rect 23673 4437 23707 4471
rect 23707 4437 23716 4471
rect 23664 4428 23716 4437
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 21548 4224 21600 4276
rect 22284 4224 22336 4276
rect 22376 4224 22428 4276
rect 21640 4156 21692 4208
rect 1492 4131 1544 4140
rect 1492 4097 1501 4131
rect 1501 4097 1535 4131
rect 1535 4097 1544 4131
rect 1492 4088 1544 4097
rect 10232 4088 10284 4140
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 22192 4088 22244 4140
rect 22468 4156 22520 4208
rect 23664 4224 23716 4276
rect 4988 4020 5040 4072
rect 18604 4020 18656 4072
rect 24216 4088 24268 4140
rect 24584 4088 24636 4140
rect 1860 3952 1912 4004
rect 20996 3952 21048 4004
rect 1032 3884 1084 3936
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 22560 3927 22612 3936
rect 22560 3893 22569 3927
rect 22569 3893 22603 3927
rect 22603 3893 22612 3927
rect 22560 3884 22612 3893
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 24124 3927 24176 3936
rect 24124 3893 24133 3927
rect 24133 3893 24167 3927
rect 24167 3893 24176 3927
rect 24124 3884 24176 3893
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 1492 3723 1544 3732
rect 1492 3689 1501 3723
rect 1501 3689 1535 3723
rect 1535 3689 1544 3723
rect 1492 3680 1544 3689
rect 1860 3680 1912 3732
rect 2044 3680 2096 3732
rect 2136 3680 2188 3732
rect 19248 3680 19300 3732
rect 20076 3680 20128 3732
rect 22560 3680 22612 3732
rect 22836 3680 22888 3732
rect 23848 3680 23900 3732
rect 25320 3680 25372 3732
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 21456 3476 21508 3528
rect 23756 3612 23808 3664
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 23848 3451 23900 3460
rect 23848 3417 23857 3451
rect 23857 3417 23891 3451
rect 23891 3417 23900 3451
rect 23848 3408 23900 3417
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 18604 3136 18656 3188
rect 19432 3136 19484 3188
rect 23664 3136 23716 3188
rect 24124 3136 24176 3188
rect 3608 3000 3660 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 22928 2932 22980 2984
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 11888 2592 11940 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 20812 2592 20864 2644
rect 23848 2592 23900 2644
rect 8576 2567 8628 2576
rect 8576 2533 8585 2567
rect 8585 2533 8619 2567
rect 8619 2533 8628 2567
rect 8576 2524 8628 2533
rect 23940 2524 23992 2576
rect 6736 2388 6788 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9588 2431 9640 2440
rect 9588 2397 9597 2431
rect 9597 2397 9631 2431
rect 9631 2397 9640 2431
rect 9588 2388 9640 2397
rect 10784 2431 10836 2440
rect 10784 2397 10793 2431
rect 10793 2397 10827 2431
rect 10827 2397 10836 2431
rect 10784 2388 10836 2397
rect 11796 2431 11848 2440
rect 11796 2397 11805 2431
rect 11805 2397 11839 2431
rect 11839 2397 11848 2431
rect 11796 2388 11848 2397
rect 12164 2431 12216 2440
rect 12164 2397 12173 2431
rect 12173 2397 12207 2431
rect 12207 2397 12216 2431
rect 12164 2388 12216 2397
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 24216 2431 24268 2440
rect 24216 2397 24225 2431
rect 24225 2397 24259 2431
rect 24259 2397 24268 2431
rect 24216 2388 24268 2397
rect 7288 2295 7340 2304
rect 7288 2261 7297 2295
rect 7297 2261 7331 2295
rect 7331 2261 7340 2295
rect 7288 2252 7340 2261
rect 24032 2320 24084 2372
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 12348 2295 12400 2304
rect 12348 2261 12357 2295
rect 12357 2261 12391 2295
rect 12391 2261 12400 2295
rect 12348 2252 12400 2261
rect 14556 2295 14608 2304
rect 14556 2261 14565 2295
rect 14565 2261 14599 2295
rect 14599 2261 14608 2295
rect 14556 2252 14608 2261
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 6736 2091 6788 2100
rect 6736 2057 6745 2091
rect 6745 2057 6779 2091
rect 6779 2057 6788 2091
rect 6736 2048 6788 2057
rect 8392 2048 8444 2100
rect 9588 2048 9640 2100
rect 10784 2048 10836 2100
rect 11796 2048 11848 2100
rect 12164 2048 12216 2100
rect 13268 2048 13320 2100
rect 14372 2048 14424 2100
rect 15476 2048 15528 2100
rect 6552 1955 6604 1964
rect 6552 1921 6561 1955
rect 6561 1921 6595 1955
rect 6595 1921 6604 1955
rect 6552 1912 6604 1921
rect 7840 1955 7892 1964
rect 7840 1921 7849 1955
rect 7849 1921 7883 1955
rect 7883 1921 7892 1955
rect 7840 1912 7892 1921
rect 9036 1955 9088 1964
rect 9036 1921 9045 1955
rect 9045 1921 9079 1955
rect 9079 1921 9088 1955
rect 9036 1912 9088 1921
rect 10232 1955 10284 1964
rect 10232 1921 10241 1955
rect 10241 1921 10275 1955
rect 10275 1921 10284 1955
rect 10232 1912 10284 1921
rect 11520 1955 11572 1964
rect 11520 1921 11529 1955
rect 11529 1921 11563 1955
rect 11563 1921 11572 1955
rect 11520 1912 11572 1921
rect 11612 1912 11664 1964
rect 12624 1955 12676 1964
rect 12624 1921 12633 1955
rect 12633 1921 12667 1955
rect 12667 1921 12676 1955
rect 12624 1912 12676 1921
rect 13820 1955 13872 1964
rect 13820 1921 13829 1955
rect 13829 1921 13863 1955
rect 13863 1921 13872 1955
rect 13820 1912 13872 1921
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 14924 1912 14976 1921
rect 2412 1844 2464 1896
rect 19800 2048 19852 2100
rect 24216 2048 24268 2100
rect 24124 1955 24176 1964
rect 24124 1921 24133 1955
rect 24133 1921 24167 1955
rect 24167 1921 24176 1955
rect 24124 1912 24176 1921
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 2412 1547 2464 1556
rect 2412 1513 2421 1547
rect 2421 1513 2455 1547
rect 2455 1513 2464 1547
rect 2412 1504 2464 1513
rect 6552 1547 6604 1556
rect 6552 1513 6561 1547
rect 6561 1513 6595 1547
rect 6595 1513 6604 1547
rect 6552 1504 6604 1513
rect 7840 1504 7892 1556
rect 9036 1504 9088 1556
rect 10232 1504 10284 1556
rect 11520 1504 11572 1556
rect 12624 1504 12676 1556
rect 14924 1504 14976 1556
rect 24124 1504 24176 1556
rect 940 1300 992 1352
rect 2228 1343 2280 1352
rect 2228 1309 2237 1343
rect 2237 1309 2271 1343
rect 2271 1309 2280 1343
rect 2228 1300 2280 1309
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 7012 1343 7064 1352
rect 7012 1309 7021 1343
rect 7021 1309 7055 1343
rect 7055 1309 7064 1343
rect 7012 1300 7064 1309
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 3608 1207 3660 1216
rect 3608 1173 3617 1207
rect 3617 1173 3651 1207
rect 3651 1173 3660 1207
rect 3608 1164 3660 1173
rect 4804 1207 4856 1216
rect 4804 1173 4813 1207
rect 4813 1173 4847 1207
rect 4847 1173 4856 1207
rect 4804 1164 4856 1173
rect 8300 1164 8352 1216
rect 9404 1343 9456 1352
rect 9404 1309 9413 1343
rect 9413 1309 9447 1343
rect 9447 1309 9456 1343
rect 9404 1300 9456 1309
rect 10416 1343 10468 1352
rect 10416 1309 10425 1343
rect 10425 1309 10459 1343
rect 10459 1309 10468 1343
rect 10416 1300 10468 1309
rect 10692 1343 10744 1352
rect 10692 1309 10701 1343
rect 10701 1309 10735 1343
rect 10735 1309 10744 1343
rect 10692 1300 10744 1309
rect 11612 1300 11664 1352
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 12716 1300 12768 1352
rect 13820 1300 13872 1352
rect 14188 1343 14240 1352
rect 14188 1309 14197 1343
rect 14197 1309 14231 1343
rect 14231 1309 14240 1343
rect 14188 1300 14240 1309
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 15568 1300 15620 1352
rect 16672 1343 16724 1352
rect 16672 1309 16681 1343
rect 16681 1309 16715 1343
rect 16715 1309 16724 1343
rect 16672 1300 16724 1309
rect 16856 1300 16908 1352
rect 17776 1343 17828 1352
rect 17776 1309 17785 1343
rect 17785 1309 17819 1343
rect 17819 1309 17828 1343
rect 17776 1300 17828 1309
rect 18052 1300 18104 1352
rect 18144 1300 18196 1352
rect 19156 1300 19208 1352
rect 19248 1343 19300 1352
rect 19248 1309 19257 1343
rect 19257 1309 19291 1343
rect 19291 1309 19300 1343
rect 19248 1300 19300 1309
rect 20168 1343 20220 1352
rect 20168 1309 20177 1343
rect 20177 1309 20211 1343
rect 20211 1309 20220 1343
rect 20168 1300 20220 1309
rect 20720 1300 20772 1352
rect 21364 1343 21416 1352
rect 21364 1309 21373 1343
rect 21373 1309 21407 1343
rect 21407 1309 21416 1343
rect 21364 1300 21416 1309
rect 21640 1300 21692 1352
rect 22560 1343 22612 1352
rect 22560 1309 22569 1343
rect 22569 1309 22603 1343
rect 22603 1309 22612 1343
rect 22560 1300 22612 1309
rect 18512 1232 18564 1284
rect 23480 1232 23532 1284
rect 23940 1343 23992 1352
rect 23940 1309 23949 1343
rect 23949 1309 23983 1343
rect 23983 1309 23992 1343
rect 23940 1300 23992 1309
rect 24492 1300 24544 1352
rect 24308 1232 24360 1284
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 4804 960 4856 1012
rect 10692 960 10744 1012
rect 8300 892 8352 944
rect 18144 960 18196 1012
<< metal2 >>
rect 202 7840 258 8000
rect 478 7840 534 8000
rect 754 7840 810 8000
rect 1030 7840 1086 8000
rect 1306 7840 1362 8000
rect 1582 7840 1638 8000
rect 1858 7840 1914 8000
rect 2134 7840 2190 8000
rect 2410 7970 2466 8000
rect 2332 7942 2466 7970
rect 216 6474 244 7840
rect 216 6446 336 6474
rect 308 5166 336 6446
rect 492 6390 520 7840
rect 480 6384 532 6390
rect 480 6326 532 6332
rect 296 5160 348 5166
rect 296 5102 348 5108
rect 768 4758 796 7840
rect 756 4752 808 4758
rect 756 4694 808 4700
rect 1044 3942 1072 7840
rect 1320 4826 1348 7840
rect 1596 5302 1624 7840
rect 1872 5370 1900 7840
rect 2148 5914 2176 7840
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1860 5364 1912 5370
rect 1860 5306 1912 5312
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1964 4690 1992 5170
rect 2240 4826 2268 6258
rect 2332 5914 2360 7942
rect 2410 7840 2466 7942
rect 2686 7840 2742 8000
rect 2962 7840 3018 8000
rect 3238 7840 3294 8000
rect 3514 7970 3570 8000
rect 3344 7942 3570 7970
rect 2700 5914 2728 7840
rect 2872 7336 2924 7342
rect 2872 7278 2924 7284
rect 2884 6390 2912 7278
rect 2976 6458 3004 7840
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 3252 5914 3280 7840
rect 3344 6254 3372 7942
rect 3514 7840 3570 7942
rect 3790 7840 3846 8000
rect 4066 7970 4122 8000
rect 4342 7970 4398 8000
rect 3896 7942 4122 7970
rect 3804 7800 3832 7840
rect 3712 7772 3832 7800
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3436 5710 3464 6870
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 2502 5264 2558 5273
rect 2502 5199 2504 5208
rect 2556 5199 2558 5208
rect 2504 5170 2556 5176
rect 3528 5030 3556 6258
rect 3608 5364 3660 5370
rect 3712 5352 3740 7772
rect 3896 7698 3924 7942
rect 4066 7840 4122 7942
rect 4172 7942 4398 7970
rect 3804 7670 3924 7698
rect 3804 5914 3832 7670
rect 4172 6474 4200 7942
rect 4342 7840 4398 7942
rect 4618 7840 4674 8000
rect 4894 7840 4950 8000
rect 5170 7840 5226 8000
rect 5446 7970 5502 8000
rect 5276 7942 5502 7970
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4080 6458 4200 6474
rect 4264 6458 4292 6802
rect 4068 6452 4200 6458
rect 4120 6446 4200 6452
rect 4252 6452 4304 6458
rect 4068 6394 4120 6400
rect 4252 6394 4304 6400
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 4356 5370 4384 6054
rect 4448 5914 4476 6258
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4540 5710 4568 7142
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 3660 5324 3740 5352
rect 4344 5364 4396 5370
rect 3608 5306 3660 5312
rect 4344 5306 4396 5312
rect 4528 5364 4580 5370
rect 4632 5352 4660 7840
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4724 5710 4752 7346
rect 4804 7132 4856 7138
rect 4804 7074 4856 7080
rect 4816 5914 4844 7074
rect 4908 5914 4936 7840
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4580 5324 4660 5352
rect 4528 5306 4580 5312
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3712 4826 3740 5170
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 4448 4826 4476 5170
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1766 4584 1822 4593
rect 1766 4519 1768 4528
rect 1820 4519 1822 4528
rect 2044 4548 2096 4554
rect 1768 4490 1820 4496
rect 2044 4490 2096 4496
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1032 3936 1084 3942
rect 1032 3878 1084 3884
rect 1504 3738 1532 4082
rect 1860 4004 1912 4010
rect 1860 3946 1912 3952
rect 1872 3738 1900 3946
rect 2056 3738 2084 4490
rect 5000 4078 5028 7346
rect 5184 6390 5212 7840
rect 5276 6458 5304 7942
rect 5446 7840 5502 7942
rect 5722 7840 5778 8000
rect 5998 7840 6054 8000
rect 6274 7840 6330 8000
rect 6550 7840 6606 8000
rect 6826 7840 6882 8000
rect 7102 7840 7158 8000
rect 7378 7840 7434 8000
rect 7654 7970 7710 8000
rect 7576 7942 7710 7970
rect 5736 6458 5764 7840
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5172 5636 5224 5642
rect 5172 5578 5224 5584
rect 5184 5370 5212 5578
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5552 5166 5580 5646
rect 5828 5370 5856 6258
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 5276 4826 5304 5102
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5920 4622 5948 7414
rect 6012 5914 6040 7840
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6196 6458 6224 6734
rect 6288 6458 6316 7840
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6564 5914 6592 7840
rect 6840 6746 6868 7840
rect 6748 6718 6868 6746
rect 7116 6746 7144 7840
rect 7116 6718 7328 6746
rect 6748 6118 6776 6718
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 7116 5658 7144 6258
rect 7196 5840 7248 5846
rect 7300 5794 7328 6718
rect 7392 6458 7420 7840
rect 7576 6458 7604 7942
rect 7654 7840 7710 7942
rect 7930 7840 7986 8000
rect 8024 7880 8076 7886
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7656 7608 7708 7614
rect 7656 7550 7708 7556
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5914 7420 6258
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7248 5788 7328 5794
rect 7196 5782 7328 5788
rect 7208 5766 7328 5782
rect 6276 5636 6328 5642
rect 7116 5630 7328 5658
rect 6276 5578 6328 5584
rect 6288 5137 6316 5578
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 7300 5234 7328 5630
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7392 5370 7420 5578
rect 7484 5370 7512 6326
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6920 5160 6972 5166
rect 6274 5128 6330 5137
rect 6920 5102 6972 5108
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7208 5114 7236 5170
rect 7576 5114 7604 6258
rect 7668 5234 7696 7550
rect 7760 5234 7788 7754
rect 7944 5914 7972 7840
rect 8206 7840 8262 8000
rect 8482 7840 8538 8000
rect 8758 7970 8814 8000
rect 8588 7942 8814 7970
rect 8024 7822 8076 7828
rect 8036 6322 8064 7822
rect 8116 7608 8168 7614
rect 8116 7550 8168 7556
rect 8128 7206 8156 7550
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8116 6996 8168 7002
rect 8116 6938 8168 6944
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8128 5914 8156 6938
rect 8220 5914 8248 7840
rect 8300 7064 8352 7070
rect 8300 7006 8352 7012
rect 8312 6390 8340 7006
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6390 8432 6598
rect 8496 6458 8524 7840
rect 8588 6458 8616 7942
rect 8758 7840 8814 7942
rect 9034 7840 9090 8000
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8760 7676 8812 7682
rect 8760 7618 8812 7624
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8392 6384 8444 6390
rect 8392 6326 8444 6332
rect 8680 5914 8708 7346
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8772 5794 8800 7618
rect 9048 5914 9076 7840
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 8588 5766 8800 5794
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5370 7880 5578
rect 8588 5370 8616 5766
rect 9140 5642 9168 7890
rect 9310 7840 9366 8000
rect 9586 7840 9642 8000
rect 9862 7840 9918 8000
rect 10138 7840 10194 8000
rect 10414 7840 10470 8000
rect 10690 7840 10746 8000
rect 10966 7840 11022 8000
rect 11242 7840 11298 8000
rect 11518 7840 11574 8000
rect 11794 7840 11850 8000
rect 12070 7840 12126 8000
rect 12346 7840 12402 8000
rect 12622 7970 12678 8000
rect 12452 7942 12678 7970
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9232 5914 9260 6802
rect 9324 6440 9352 7840
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9404 6452 9456 6458
rect 9324 6412 9404 6440
rect 9404 6394 9456 6400
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 8680 5370 8708 5578
rect 9324 5370 9352 6258
rect 9508 5778 9536 6802
rect 9600 6390 9628 7840
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6934 9720 7142
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9784 6458 9812 6870
rect 9876 6458 9904 7840
rect 10152 7426 10180 7840
rect 10152 7398 10364 7426
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9600 5234 9628 6122
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 9864 5840 9916 5846
rect 9678 5808 9734 5817
rect 10048 5840 10100 5846
rect 9916 5788 10048 5794
rect 9864 5782 10100 5788
rect 9876 5766 10088 5782
rect 9678 5743 9734 5752
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 6274 5063 6330 5072
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4826 6776 4966
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6932 4758 6960 5102
rect 7024 4826 7052 5102
rect 7208 5086 7604 5114
rect 9692 5098 9720 5743
rect 9956 5704 10008 5710
rect 10138 5672 10194 5681
rect 10008 5652 10138 5658
rect 9956 5646 10138 5652
rect 9968 5630 10138 5646
rect 10138 5607 10194 5616
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9956 5568 10008 5574
rect 10244 5522 10272 6258
rect 9956 5510 10008 5516
rect 9770 5400 9826 5409
rect 9876 5370 9904 5510
rect 9770 5335 9826 5344
rect 9864 5364 9916 5370
rect 9784 5302 9812 5335
rect 9864 5306 9916 5312
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9968 5012 9996 5510
rect 10152 5494 10272 5522
rect 10336 5522 10364 7398
rect 10428 5710 10456 7840
rect 10704 6610 10732 7840
rect 10784 7540 10836 7546
rect 10784 7482 10836 7488
rect 10612 6582 10732 6610
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10336 5494 10456 5522
rect 10152 5370 10180 5494
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10428 5234 10456 5494
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 9784 4984 9996 5012
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 9784 4690 9812 4984
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 10244 4146 10272 5170
rect 10520 5166 10548 6258
rect 10612 5522 10640 6582
rect 10796 5574 10824 7482
rect 10876 7336 10928 7342
rect 10876 7278 10928 7284
rect 10888 6458 10916 7278
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10876 5704 10928 5710
rect 10980 5692 11008 7840
rect 11152 7608 11204 7614
rect 11152 7550 11204 7556
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 6458 11100 7414
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 11058 6216 11114 6225
rect 11058 6151 11060 6160
rect 11112 6151 11114 6160
rect 11060 6122 11112 6128
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5710 11100 5782
rect 10928 5664 11008 5692
rect 11060 5704 11112 5710
rect 10876 5646 10928 5652
rect 11060 5646 11112 5652
rect 10784 5568 10836 5574
rect 10612 5494 10732 5522
rect 10784 5510 10836 5516
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10704 5234 10732 5494
rect 11072 5370 11100 5510
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 11164 5030 11192 7550
rect 11256 6610 11284 7840
rect 11256 6582 11468 6610
rect 11336 6180 11388 6186
rect 11336 6122 11388 6128
rect 11348 5710 11376 6122
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11440 5234 11468 6582
rect 11532 5710 11560 7840
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11716 6322 11744 7278
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 11716 5574 11744 6054
rect 11808 5710 11836 7840
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11612 5568 11664 5574
rect 11612 5510 11664 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 10796 4690 10824 4966
rect 11624 4758 11652 5510
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3738 2176 3878
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 3608 3052 3660 3058
rect 3608 2994 3660 3000
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2424 1562 2452 1838
rect 2412 1556 2464 1562
rect 2412 1498 2464 1504
rect 940 1352 992 1358
rect 940 1294 992 1300
rect 2228 1352 2280 1358
rect 3424 1352 3476 1358
rect 2228 1294 2280 1300
rect 3344 1312 3424 1340
rect 952 160 980 1294
rect 938 0 994 160
rect 2134 82 2190 160
rect 2240 82 2268 1294
rect 3344 160 3372 1312
rect 3424 1294 3476 1300
rect 3620 1222 3648 2994
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 11900 2650 11928 7414
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11992 5778 12020 6054
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12084 5710 12112 7840
rect 12360 7342 12388 7840
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5409 12020 5510
rect 11978 5400 12034 5409
rect 11978 5335 12034 5344
rect 12176 4826 12204 6054
rect 12268 5914 12296 7210
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12360 5370 12388 6938
rect 12452 6390 12480 7942
rect 12622 7840 12678 7942
rect 12898 7970 12954 8000
rect 12898 7942 13124 7970
rect 12898 7840 12954 7942
rect 13096 7562 13124 7942
rect 13174 7840 13230 8000
rect 13450 7840 13506 8000
rect 13726 7970 13782 8000
rect 13648 7942 13782 7970
rect 13188 7800 13216 7840
rect 13188 7772 13308 7800
rect 13096 7534 13216 7562
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6458 12664 7142
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12808 6452 12860 6458
rect 12992 6452 13044 6458
rect 12860 6412 12992 6440
rect 12808 6394 12860 6400
rect 12992 6394 13044 6400
rect 12440 6384 12492 6390
rect 12440 6326 12492 6332
rect 12622 6352 12678 6361
rect 12622 6287 12624 6296
rect 12676 6287 12678 6296
rect 12808 6316 12860 6322
rect 12624 6258 12676 6264
rect 12808 6258 12860 6264
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 12532 6248 12584 6254
rect 12716 6248 12768 6254
rect 12584 6196 12716 6202
rect 12532 6190 12768 6196
rect 12544 6174 12756 6190
rect 12820 6118 12848 6258
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12544 5778 12572 6054
rect 13096 5914 13124 6258
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5681 12756 5714
rect 13084 5704 13136 5710
rect 12714 5672 12770 5681
rect 13188 5692 13216 7534
rect 13136 5664 13216 5692
rect 13280 5692 13308 7772
rect 13360 6316 13412 6322
rect 13464 6304 13492 7840
rect 13648 6322 13676 7942
rect 13726 7840 13782 7942
rect 14002 7970 14058 8000
rect 14002 7942 14228 7970
rect 14002 7840 14058 7942
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14108 6798 14136 6938
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14200 6390 14228 7942
rect 14278 7840 14334 8000
rect 14554 7840 14610 8000
rect 14830 7840 14886 8000
rect 15106 7840 15162 8000
rect 15382 7840 15438 8000
rect 15658 7840 15714 8000
rect 15934 7840 15990 8000
rect 16210 7840 16266 8000
rect 16486 7840 16542 8000
rect 16762 7840 16818 8000
rect 17038 7840 17094 8000
rect 17314 7840 17370 8000
rect 17590 7840 17646 8000
rect 17866 7970 17922 8000
rect 17788 7942 17922 7970
rect 14188 6384 14240 6390
rect 14002 6352 14058 6361
rect 13412 6276 13492 6304
rect 13636 6316 13688 6322
rect 13360 6258 13412 6264
rect 14188 6326 14240 6332
rect 14002 6287 14058 6296
rect 13636 6258 13688 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13452 5704 13504 5710
rect 13280 5664 13452 5692
rect 13084 5646 13136 5652
rect 13452 5646 13504 5652
rect 12714 5607 12770 5616
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12164 4820 12216 4826
rect 12164 4762 12216 4768
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 13464 2650 13492 4490
rect 13740 4486 13768 6054
rect 14016 5574 14044 6287
rect 14292 5710 14320 7840
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14384 5273 14412 6054
rect 14568 5692 14596 7840
rect 14844 6866 14872 7840
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14752 5914 14780 6802
rect 15120 6458 15148 7840
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 14832 5704 14884 5710
rect 14568 5664 14832 5692
rect 14832 5646 14884 5652
rect 14370 5264 14426 5273
rect 14370 5199 14426 5208
rect 15212 4593 15240 6054
rect 15396 5624 15424 7840
rect 15672 6882 15700 7840
rect 15580 6854 15700 6882
rect 15948 6866 15976 7840
rect 15752 6860 15804 6866
rect 15476 5636 15528 5642
rect 15396 5596 15476 5624
rect 15476 5578 15528 5584
rect 15580 5556 15608 6854
rect 15752 6802 15804 6808
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15764 6322 15792 6802
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15672 5914 15700 6258
rect 16118 6216 16174 6225
rect 16118 6151 16120 6160
rect 16172 6151 16174 6160
rect 16120 6122 16172 6128
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 16224 5624 16252 7840
rect 16500 7018 16528 7840
rect 16316 6990 16528 7018
rect 16316 5846 16344 6990
rect 16776 6866 16804 7840
rect 16948 6928 17000 6934
rect 16948 6870 17000 6876
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16408 5692 16436 6802
rect 16960 6458 16988 6870
rect 17052 6662 17080 7840
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17328 6458 17356 7840
rect 17408 7676 17460 7682
rect 17408 7618 17460 7624
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16500 5914 16528 6258
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16488 5704 16540 5710
rect 16408 5664 16488 5692
rect 16488 5646 16540 5652
rect 16304 5636 16356 5642
rect 16224 5596 16304 5624
rect 16304 5578 16356 5584
rect 15660 5568 15712 5574
rect 15580 5528 15660 5556
rect 15660 5510 15712 5516
rect 16684 5166 16712 6122
rect 16868 5914 16896 6258
rect 17420 5914 17448 7618
rect 17604 7290 17632 7840
rect 17604 7262 17724 7290
rect 17696 7206 17724 7262
rect 17684 7200 17736 7206
rect 17684 7142 17736 7148
rect 17500 7132 17552 7138
rect 17500 7074 17552 7080
rect 17512 6186 17540 7074
rect 17500 6180 17552 6186
rect 17500 6122 17552 6128
rect 17788 5914 17816 7942
rect 17866 7840 17922 7942
rect 18142 7840 18198 8000
rect 18418 7970 18474 8000
rect 18418 7942 18552 7970
rect 18418 7840 18474 7942
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17316 5840 17368 5846
rect 17314 5808 17316 5817
rect 17368 5808 17370 5817
rect 17314 5743 17370 5752
rect 17972 5574 18000 7754
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18064 6322 18092 6802
rect 18156 6730 18184 7840
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18248 6361 18276 7686
rect 18420 7200 18472 7206
rect 18420 7142 18472 7148
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18234 6352 18290 6361
rect 18052 6316 18104 6322
rect 18340 6322 18368 6598
rect 18432 6390 18460 7142
rect 18420 6384 18472 6390
rect 18420 6326 18472 6332
rect 18234 6287 18290 6296
rect 18328 6316 18380 6322
rect 18052 6258 18104 6264
rect 18328 6258 18380 6264
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 18340 5574 18368 5850
rect 18432 5710 18460 6122
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 18418 5536 18474 5545
rect 17880 5370 17908 5510
rect 18418 5471 18474 5480
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 18432 5302 18460 5471
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18524 5234 18552 7942
rect 18694 7840 18750 8000
rect 18970 7970 19026 8000
rect 18970 7942 19196 7970
rect 18970 7840 19026 7942
rect 18708 6644 18736 7840
rect 18616 6616 18736 6644
rect 18616 6440 18644 6616
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 18616 6412 18736 6440
rect 18604 6112 18656 6118
rect 18604 6054 18656 6060
rect 18616 5846 18644 6054
rect 18604 5840 18656 5846
rect 18604 5782 18656 5788
rect 18604 5704 18656 5710
rect 18708 5681 18736 6412
rect 18972 6384 19024 6390
rect 18786 6352 18842 6361
rect 18972 6326 19024 6332
rect 18786 6287 18842 6296
rect 18800 5914 18828 6287
rect 18880 6112 18932 6118
rect 18880 6054 18932 6060
rect 18892 5914 18920 6054
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 5681 19012 6326
rect 18604 5646 18656 5652
rect 18694 5672 18750 5681
rect 18616 5370 18644 5646
rect 18694 5607 18750 5616
rect 18970 5672 19026 5681
rect 18970 5607 19026 5616
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 19168 5250 19196 7942
rect 19246 7840 19302 8000
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19340 7880 19392 7886
rect 19260 5522 19288 7840
rect 19340 7822 19392 7828
rect 19352 6458 19380 7822
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19444 6338 19472 7890
rect 19522 7840 19578 8000
rect 19798 7840 19854 8000
rect 20074 7840 20130 8000
rect 20350 7840 20406 8000
rect 20626 7840 20682 8000
rect 20902 7970 20958 8000
rect 21178 7970 21234 8000
rect 20902 7942 21128 7970
rect 20902 7840 20958 7942
rect 19536 6390 19564 7840
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19352 6310 19472 6338
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19352 5914 19380 6310
rect 19628 6202 19656 6734
rect 19708 6724 19760 6730
rect 19708 6666 19760 6672
rect 19720 6322 19748 6666
rect 19812 6610 19840 7840
rect 19812 6582 20024 6610
rect 19996 6338 20024 6582
rect 20088 6458 20116 7840
rect 20364 7018 20392 7840
rect 20536 7064 20588 7070
rect 20364 6990 20484 7018
rect 20536 7006 20588 7012
rect 20456 6458 20484 6990
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19892 6316 19944 6322
rect 19996 6310 20208 6338
rect 19892 6258 19944 6264
rect 19536 6174 19656 6202
rect 19536 5914 19564 6174
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5914 19656 6054
rect 19340 5908 19392 5914
rect 19340 5850 19392 5856
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19260 5494 19380 5522
rect 19246 5400 19302 5409
rect 19246 5335 19248 5344
rect 19300 5335 19302 5344
rect 19248 5306 19300 5312
rect 19076 5234 19196 5250
rect 19352 5234 19380 5494
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 19064 5228 19196 5234
rect 19116 5222 19196 5228
rect 19340 5228 19392 5234
rect 19064 5170 19116 5176
rect 19340 5170 19392 5176
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 18512 5024 18564 5030
rect 18512 4966 18564 4972
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15198 4584 15254 4593
rect 15198 4519 15254 4528
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 8576 2576 8628 2582
rect 8574 2544 8576 2553
rect 8628 2544 8630 2553
rect 8574 2479 8630 2488
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 10784 2440 10836 2446
rect 10784 2382 10836 2388
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 12164 2440 12216 2446
rect 13268 2440 13320 2446
rect 12164 2382 12216 2388
rect 12346 2408 12402 2417
rect 6748 2106 6776 2382
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 7300 2009 7328 2246
rect 8404 2106 8432 2382
rect 9600 2106 9628 2382
rect 10796 2106 10824 2382
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 10784 2100 10836 2106
rect 10784 2042 10836 2048
rect 7286 2000 7342 2009
rect 6552 1964 6604 1970
rect 7286 1935 7342 1944
rect 7840 1964 7892 1970
rect 6552 1906 6604 1912
rect 7840 1906 7892 1912
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 6564 1562 6592 1906
rect 7852 1562 7880 1906
rect 9048 1562 9076 1906
rect 9851 1660 10159 1669
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 10244 1562 10272 1906
rect 10980 1873 11008 2246
rect 11808 2106 11836 2382
rect 12176 2106 12204 2382
rect 13268 2382 13320 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 12346 2343 12402 2352
rect 12360 2310 12388 2343
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 13280 2106 13308 2382
rect 14384 2106 14412 2382
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 11796 2100 11848 2106
rect 11796 2042 11848 2048
rect 12164 2100 12216 2106
rect 12164 2042 12216 2048
rect 13268 2100 13320 2106
rect 13268 2042 13320 2048
rect 14372 2100 14424 2106
rect 14372 2042 14424 2048
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 10966 1864 11022 1873
rect 10966 1799 11022 1808
rect 11532 1562 11560 1906
rect 6552 1556 6604 1562
rect 6552 1498 6604 1504
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 10232 1556 10284 1562
rect 10232 1498 10284 1504
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11624 1358 11652 1906
rect 12636 1562 12664 1906
rect 12624 1556 12676 1562
rect 12624 1498 12676 1504
rect 13832 1358 13860 1906
rect 14568 1465 14596 2246
rect 15488 2106 15516 2382
rect 15476 2100 15528 2106
rect 15476 2042 15528 2048
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 14936 1562 14964 1906
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 14554 1456 14610 1465
rect 14554 1391 14610 1400
rect 15580 1358 15608 4694
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16868 1358 16896 4558
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18064 1358 18092 2994
rect 4620 1352 4672 1358
rect 5816 1352 5868 1358
rect 4620 1294 4672 1300
rect 5736 1312 5816 1340
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 2134 54 2268 82
rect 2134 0 2190 54
rect 3330 0 3386 160
rect 4526 82 4582 160
rect 4632 82 4660 1294
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4816 1018 4844 1158
rect 4804 1012 4856 1018
rect 4804 954 4856 960
rect 5736 160 5764 1312
rect 5816 1294 5868 1300
rect 7012 1352 7064 1358
rect 8208 1352 8260 1358
rect 7064 1312 7328 1340
rect 7012 1294 7064 1300
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 4526 54 4660 82
rect 4526 0 4582 54
rect 5722 0 5778 160
rect 6918 82 6974 160
rect 7300 82 7328 1312
rect 8128 1312 8208 1340
rect 8128 160 8156 1312
rect 9404 1352 9456 1358
rect 8208 1294 8260 1300
rect 9324 1312 9404 1340
rect 8300 1216 8352 1222
rect 8300 1158 8352 1164
rect 8312 950 8340 1158
rect 8300 944 8352 950
rect 8300 886 8352 892
rect 9324 160 9352 1312
rect 9404 1294 9456 1300
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 11612 1352 11664 1358
rect 11796 1352 11848 1358
rect 11612 1294 11664 1300
rect 11716 1312 11796 1340
rect 6918 54 7328 82
rect 6918 0 6974 54
rect 8114 0 8170 160
rect 9310 0 9366 160
rect 10428 82 10456 1294
rect 10704 1018 10732 1294
rect 10692 1012 10744 1018
rect 10692 954 10744 960
rect 11716 160 11744 1312
rect 11796 1294 11848 1300
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 13820 1352 13872 1358
rect 13820 1294 13872 1300
rect 14188 1352 14240 1358
rect 14188 1294 14240 1300
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15568 1352 15620 1358
rect 16672 1352 16724 1358
rect 15568 1294 15620 1300
rect 16500 1312 16672 1340
rect 10506 82 10562 160
rect 10428 54 10562 82
rect 10506 0 10562 54
rect 11702 0 11758 160
rect 12728 82 12756 1294
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12898 82 12954 160
rect 12728 54 12954 82
rect 12898 0 12954 54
rect 14094 82 14150 160
rect 14200 82 14228 1294
rect 14094 54 14228 82
rect 15290 82 15346 160
rect 15396 82 15424 1294
rect 16500 160 16528 1312
rect 16672 1294 16724 1300
rect 16856 1352 16908 1358
rect 17776 1352 17828 1358
rect 16856 1294 16908 1300
rect 17696 1312 17776 1340
rect 17696 160 17724 1312
rect 17776 1294 17828 1300
rect 18052 1352 18104 1358
rect 18052 1294 18104 1300
rect 18144 1352 18196 1358
rect 18144 1294 18196 1300
rect 18156 1018 18184 1294
rect 18524 1290 18552 4966
rect 19812 4826 19840 5170
rect 19904 5098 19932 6258
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19996 5370 20024 5646
rect 20076 5568 20128 5574
rect 20076 5510 20128 5516
rect 20088 5370 20116 5510
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20180 5302 20208 6310
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20168 5296 20220 5302
rect 20168 5238 20220 5244
rect 20074 5128 20130 5137
rect 19892 5092 19944 5098
rect 20074 5063 20076 5072
rect 19892 5034 19944 5040
rect 20128 5063 20130 5072
rect 20076 5034 20128 5040
rect 20272 5030 20300 6258
rect 20548 5556 20576 7006
rect 20640 5846 20668 7840
rect 21100 7698 21128 7942
rect 21178 7942 21404 7970
rect 21178 7840 21234 7942
rect 21100 7670 21312 7698
rect 21284 6458 21312 7670
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21376 6390 21404 7942
rect 21454 7840 21510 8000
rect 21730 7970 21786 8000
rect 21730 7942 21956 7970
rect 21730 7840 21786 7942
rect 21468 7800 21496 7840
rect 21928 7818 21956 7942
rect 22006 7840 22062 8000
rect 22282 7840 22338 8000
rect 22558 7840 22614 8000
rect 22834 7840 22890 8000
rect 23110 7840 23166 8000
rect 23386 7840 23442 8000
rect 23662 7840 23718 8000
rect 23938 7970 23994 8000
rect 23860 7942 23994 7970
rect 21916 7812 21968 7818
rect 21468 7772 21864 7800
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20628 5568 20680 5574
rect 20548 5528 20628 5556
rect 20628 5510 20680 5516
rect 20720 5228 20772 5234
rect 20720 5170 20772 5176
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18616 4078 18644 4422
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 19260 4264 19288 4558
rect 19168 4236 19288 4264
rect 18604 4072 18656 4078
rect 18604 4014 18656 4020
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18616 3194 18644 3470
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 19168 1358 19196 4236
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19260 3738 19288 4082
rect 20088 3738 20116 4082
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19812 2106 19840 2382
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 20732 1358 20760 5170
rect 20824 2650 20852 6258
rect 21100 5710 21128 6326
rect 21560 6322 21588 7414
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 20916 5030 20944 5578
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 21008 4010 21036 5578
rect 21468 5370 21496 6258
rect 21836 6118 21864 7772
rect 21916 7754 21968 7760
rect 22020 6202 22048 7840
rect 22020 6174 22140 6202
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21652 5914 21680 6054
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 21640 5908 21692 5914
rect 22112 5896 22140 6174
rect 22296 5914 22324 7840
rect 22468 6316 22520 6322
rect 22468 6258 22520 6264
rect 21640 5850 21692 5856
rect 22020 5868 22140 5896
rect 22284 5908 22336 5914
rect 21916 5636 21968 5642
rect 21916 5578 21968 5584
rect 21928 5370 21956 5578
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21468 3534 21496 5170
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21560 4282 21588 4558
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21652 4214 21680 5170
rect 22020 5114 22048 5868
rect 22284 5850 22336 5856
rect 22480 5817 22508 6258
rect 22466 5808 22522 5817
rect 22466 5743 22522 5752
rect 22466 5672 22522 5681
rect 22466 5607 22468 5616
rect 22520 5607 22522 5616
rect 22468 5578 22520 5584
rect 22020 5086 22232 5114
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 22204 4758 22232 5086
rect 22468 5024 22520 5030
rect 22468 4966 22520 4972
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22192 4752 22244 4758
rect 22192 4694 22244 4700
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 21836 4026 21864 4558
rect 22192 4480 22244 4486
rect 22192 4422 22244 4428
rect 22284 4480 22336 4486
rect 22284 4422 22336 4428
rect 22204 4146 22232 4422
rect 22296 4282 22324 4422
rect 22388 4282 22416 4762
rect 22284 4276 22336 4282
rect 22284 4218 22336 4224
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22480 4214 22508 4966
rect 22572 4826 22600 7840
rect 22848 5914 22876 7840
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 23032 6225 23060 6258
rect 23018 6216 23074 6225
rect 23018 6151 23074 6160
rect 22836 5908 22888 5914
rect 23124 5896 23152 7840
rect 23400 6066 23428 7840
rect 23480 7812 23532 7818
rect 23480 7754 23532 7760
rect 23492 6458 23520 7754
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23400 6038 23612 6066
rect 23480 5908 23532 5914
rect 23124 5868 23480 5896
rect 22836 5850 22888 5856
rect 23480 5850 23532 5856
rect 23018 5672 23074 5681
rect 23018 5607 23020 5616
rect 23072 5607 23074 5616
rect 23020 5578 23072 5584
rect 23584 5370 23612 6038
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 22560 4820 22612 4826
rect 22560 4762 22612 4768
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 21652 3998 21864 4026
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21652 1358 21680 3998
rect 22560 3936 22612 3942
rect 22560 3878 22612 3884
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 22572 3738 22600 3878
rect 22848 3738 22876 3878
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22940 2990 22968 5170
rect 23676 4826 23704 7840
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23664 4820 23716 4826
rect 23664 4762 23716 4768
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 23020 4548 23072 4554
rect 23020 4490 23072 4496
rect 23032 4185 23060 4490
rect 23018 4176 23074 4185
rect 23018 4111 23074 4120
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 19156 1352 19208 1358
rect 19156 1294 19208 1300
rect 19248 1352 19300 1358
rect 20168 1352 20220 1358
rect 19248 1294 19300 1300
rect 20088 1312 20168 1340
rect 18512 1284 18564 1290
rect 18512 1226 18564 1232
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 18144 1012 18196 1018
rect 18144 954 18196 960
rect 18892 190 19012 218
rect 18892 160 18920 190
rect 15290 54 15424 82
rect 14094 0 14150 54
rect 15290 0 15346 54
rect 16486 0 16542 160
rect 17682 0 17738 160
rect 18878 0 18934 160
rect 18984 82 19012 190
rect 19260 82 19288 1294
rect 20088 160 20116 1312
rect 20168 1294 20220 1300
rect 20720 1352 20772 1358
rect 20720 1294 20772 1300
rect 21364 1352 21416 1358
rect 21364 1294 21416 1300
rect 21640 1352 21692 1358
rect 21640 1294 21692 1300
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 18984 54 19288 82
rect 20074 0 20130 160
rect 21270 82 21326 160
rect 21376 82 21404 1294
rect 21270 54 21404 82
rect 22466 82 22522 160
rect 22572 82 22600 1294
rect 23492 1290 23520 4558
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23676 4282 23704 4422
rect 23664 4276 23716 4282
rect 23664 4218 23716 4224
rect 23768 3670 23796 5170
rect 23860 5098 23888 7942
rect 23938 7840 23994 7942
rect 24214 7840 24270 8000
rect 24490 7970 24546 8000
rect 24766 7970 24822 8000
rect 24320 7942 24546 7970
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 24044 5658 24072 6258
rect 23940 5636 23992 5642
rect 24044 5630 24164 5658
rect 23940 5578 23992 5584
rect 23848 5092 23900 5098
rect 23848 5034 23900 5040
rect 23848 4548 23900 4554
rect 23848 4490 23900 4496
rect 23860 3738 23888 4490
rect 23848 3732 23900 3738
rect 23848 3674 23900 3680
rect 23756 3664 23808 3670
rect 23756 3606 23808 3612
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23676 3194 23704 3470
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23860 2650 23888 3402
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 23952 2582 23980 5578
rect 24032 5568 24084 5574
rect 24032 5510 24084 5516
rect 24044 5302 24072 5510
rect 24032 5296 24084 5302
rect 24032 5238 24084 5244
rect 24136 4570 24164 5630
rect 24044 4542 24164 4570
rect 23940 2576 23992 2582
rect 23940 2518 23992 2524
rect 24044 2378 24072 4542
rect 24228 4146 24256 7840
rect 24320 5030 24348 7942
rect 24490 7840 24546 7942
rect 24596 7942 24822 7970
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 24596 4146 24624 7942
rect 24766 7840 24822 7942
rect 25042 7840 25098 8000
rect 25318 7840 25374 8000
rect 25594 7840 25650 8000
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 25056 5166 25084 7840
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 24136 3194 24164 3878
rect 25332 3738 25360 7840
rect 25608 5914 25636 7840
rect 25596 5908 25648 5914
rect 25596 5850 25648 5856
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 24032 2372 24084 2378
rect 24032 2314 24084 2320
rect 24228 2106 24256 2382
rect 24216 2100 24268 2106
rect 24216 2042 24268 2048
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24136 1562 24164 1906
rect 24124 1556 24176 1562
rect 24124 1498 24176 1504
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 23480 1284 23532 1290
rect 23480 1226 23532 1232
rect 23676 190 23796 218
rect 23676 160 23704 190
rect 22466 54 22600 82
rect 21270 0 21326 54
rect 22466 0 22522 54
rect 23662 0 23718 160
rect 23768 82 23796 190
rect 23952 82 23980 1294
rect 24320 1290 24348 2994
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24492 1352 24544 1358
rect 24492 1294 24544 1300
rect 24308 1284 24360 1290
rect 24308 1226 24360 1232
rect 23768 54 23980 82
rect 24504 82 24532 1294
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 24858 82 24914 160
rect 24504 54 24914 82
rect 24858 0 24914 54
<< via2 >>
rect 2502 5228 2558 5264
rect 2502 5208 2504 5228
rect 2504 5208 2556 5228
rect 2556 5208 2558 5228
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 1766 4548 1822 4584
rect 1766 4528 1768 4548
rect 1768 4528 1820 4548
rect 1820 4528 1822 4548
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 6274 5072 6330 5128
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 9678 5752 9734 5808
rect 10138 5616 10194 5672
rect 9770 5344 9826 5400
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 11058 6180 11114 6216
rect 11058 6160 11060 6180
rect 11060 6160 11112 6180
rect 11112 6160 11114 6180
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 11978 5344 12034 5400
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 12622 6316 12678 6352
rect 12622 6296 12624 6316
rect 12624 6296 12676 6316
rect 12676 6296 12678 6316
rect 12714 5616 12770 5672
rect 14002 6296 14058 6352
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 14370 5208 14426 5264
rect 16118 6180 16174 6216
rect 16118 6160 16120 6180
rect 16120 6160 16172 6180
rect 16172 6160 16174 6180
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 17314 5788 17316 5808
rect 17316 5788 17368 5808
rect 17368 5788 17370 5808
rect 17314 5752 17370 5788
rect 18234 6296 18290 6352
rect 18418 5480 18474 5536
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 18786 6296 18842 6352
rect 18694 5616 18750 5672
rect 18970 5616 19026 5672
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 19246 5364 19302 5400
rect 19246 5344 19248 5364
rect 19248 5344 19300 5364
rect 19300 5344 19302 5364
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 15198 4528 15254 4584
rect 8574 2524 8576 2544
rect 8576 2524 8628 2544
rect 8628 2524 8630 2544
rect 8574 2488 8630 2524
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 7286 1944 7342 2000
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 12346 2352 12402 2408
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 10966 1808 11022 1864
rect 14554 1400 14610 1456
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 20074 5092 20130 5128
rect 20074 5072 20076 5092
rect 20076 5072 20128 5092
rect 20128 5072 20130 5092
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 22466 5752 22522 5808
rect 22466 5636 22522 5672
rect 22466 5616 22468 5636
rect 22468 5616 22520 5636
rect 22520 5616 22522 5636
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 23018 6160 23074 6216
rect 23018 5636 23074 5672
rect 23018 5616 23020 5636
rect 23020 5616 23072 5636
rect 23072 5616 23074 5636
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 23018 4120 23074 4176
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
<< metal3 >>
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 12617 6354 12683 6357
rect 13997 6354 14063 6357
rect 12617 6352 14063 6354
rect 12617 6296 12622 6352
rect 12678 6296 14002 6352
rect 14058 6296 14063 6352
rect 12617 6294 14063 6296
rect 12617 6291 12683 6294
rect 13997 6291 14063 6294
rect 18229 6354 18295 6357
rect 18781 6354 18847 6357
rect 18229 6352 18847 6354
rect 18229 6296 18234 6352
rect 18290 6296 18786 6352
rect 18842 6296 18847 6352
rect 18229 6294 18847 6296
rect 18229 6291 18295 6294
rect 18781 6291 18847 6294
rect 11053 6218 11119 6221
rect 16113 6218 16179 6221
rect 11053 6216 16179 6218
rect 11053 6160 11058 6216
rect 11114 6160 16118 6216
rect 16174 6160 16179 6216
rect 11053 6158 16179 6160
rect 11053 6155 11119 6158
rect 16113 6155 16179 6158
rect 19742 6156 19748 6220
rect 19812 6218 19818 6220
rect 23013 6218 23079 6221
rect 19812 6216 23079 6218
rect 19812 6160 23018 6216
rect 23074 6160 23079 6216
rect 19812 6158 23079 6160
rect 19812 6156 19818 6158
rect 23013 6155 23079 6158
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 9673 5810 9739 5813
rect 17309 5810 17375 5813
rect 9673 5808 17375 5810
rect 9673 5752 9678 5808
rect 9734 5752 17314 5808
rect 17370 5752 17375 5808
rect 9673 5750 17375 5752
rect 9673 5747 9739 5750
rect 17309 5747 17375 5750
rect 19558 5748 19564 5812
rect 19628 5810 19634 5812
rect 22461 5810 22527 5813
rect 19628 5808 22527 5810
rect 19628 5752 22466 5808
rect 22522 5752 22527 5808
rect 19628 5750 22527 5752
rect 19628 5748 19634 5750
rect 22461 5747 22527 5750
rect 10133 5674 10199 5677
rect 12709 5674 12775 5677
rect 18689 5674 18755 5677
rect 10133 5672 12775 5674
rect 10133 5616 10138 5672
rect 10194 5616 12714 5672
rect 12770 5616 12775 5672
rect 10133 5614 12775 5616
rect 10133 5611 10199 5614
rect 12709 5611 12775 5614
rect 18462 5672 18755 5674
rect 18462 5616 18694 5672
rect 18750 5616 18755 5672
rect 18462 5614 18755 5616
rect 18462 5541 18522 5614
rect 18689 5611 18755 5614
rect 18965 5674 19031 5677
rect 18965 5672 19258 5674
rect 18965 5616 18970 5672
rect 19026 5616 19258 5672
rect 18965 5614 19258 5616
rect 18965 5611 19031 5614
rect 18413 5536 18522 5541
rect 18413 5480 18418 5536
rect 18474 5480 18522 5536
rect 18413 5478 18522 5480
rect 18413 5475 18479 5478
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 19198 5405 19258 5614
rect 22134 5612 22140 5676
rect 22204 5674 22210 5676
rect 22461 5674 22527 5677
rect 22204 5672 22527 5674
rect 22204 5616 22466 5672
rect 22522 5616 22527 5672
rect 22204 5614 22527 5616
rect 22204 5612 22210 5614
rect 22461 5611 22527 5614
rect 22686 5612 22692 5676
rect 22756 5674 22762 5676
rect 23013 5674 23079 5677
rect 22756 5672 23079 5674
rect 22756 5616 23018 5672
rect 23074 5616 23079 5672
rect 22756 5614 23079 5616
rect 22756 5612 22762 5614
rect 23013 5611 23079 5614
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 9765 5402 9831 5405
rect 11973 5402 12039 5405
rect 9765 5400 12039 5402
rect 9765 5344 9770 5400
rect 9826 5344 11978 5400
rect 12034 5344 12039 5400
rect 9765 5342 12039 5344
rect 19198 5400 19307 5405
rect 19198 5344 19246 5400
rect 19302 5344 19307 5400
rect 19198 5342 19307 5344
rect 9765 5339 9831 5342
rect 11973 5339 12039 5342
rect 19241 5339 19307 5342
rect 2497 5266 2563 5269
rect 14365 5266 14431 5269
rect 2497 5264 14431 5266
rect 2497 5208 2502 5264
rect 2558 5208 14370 5264
rect 14426 5208 14431 5264
rect 2497 5206 14431 5208
rect 2497 5203 2563 5206
rect 14365 5203 14431 5206
rect 6269 5130 6335 5133
rect 20069 5130 20135 5133
rect 6269 5128 20135 5130
rect 6269 5072 6274 5128
rect 6330 5072 20074 5128
rect 20130 5072 20135 5128
rect 6269 5070 20135 5072
rect 6269 5067 6335 5070
rect 20069 5067 20135 5070
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 1761 4586 1827 4589
rect 15193 4586 15259 4589
rect 1761 4584 15259 4586
rect 1761 4528 1766 4584
rect 1822 4528 15198 4584
rect 15254 4528 15259 4584
rect 1761 4526 15259 4528
rect 1761 4523 1827 4526
rect 15193 4523 15259 4526
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 17902 4116 17908 4180
rect 17972 4178 17978 4180
rect 23013 4178 23079 4181
rect 17972 4176 23079 4178
rect 17972 4120 23018 4176
rect 23074 4120 23079 4176
rect 17972 4118 23079 4120
rect 17972 4116 17978 4118
rect 23013 4115 23079 4118
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 8569 2546 8635 2549
rect 19742 2546 19748 2548
rect 8569 2544 19748 2546
rect 8569 2488 8574 2544
rect 8630 2488 19748 2544
rect 8569 2486 19748 2488
rect 8569 2483 8635 2486
rect 19742 2484 19748 2486
rect 19812 2484 19818 2548
rect 12341 2410 12407 2413
rect 22134 2410 22140 2412
rect 12341 2408 22140 2410
rect 12341 2352 12346 2408
rect 12402 2352 22140 2408
rect 12341 2350 22140 2352
rect 12341 2347 12407 2350
rect 22134 2348 22140 2350
rect 22204 2348 22210 2412
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 7281 2002 7347 2005
rect 19558 2002 19564 2004
rect 7281 2000 19564 2002
rect 7281 1944 7286 2000
rect 7342 1944 19564 2000
rect 7281 1942 19564 1944
rect 7281 1939 7347 1942
rect 19558 1940 19564 1942
rect 19628 1940 19634 2004
rect 10961 1866 11027 1869
rect 17902 1866 17908 1868
rect 10961 1864 17908 1866
rect 10961 1808 10966 1864
rect 11022 1808 17908 1864
rect 10961 1806 17908 1808
rect 10961 1803 11027 1806
rect 17902 1804 17908 1806
rect 17972 1804 17978 1868
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 14549 1458 14615 1461
rect 22686 1458 22692 1460
rect 14549 1456 22692 1458
rect 14549 1400 14554 1456
rect 14610 1400 22692 1456
rect 14549 1398 22692 1400
rect 14549 1395 14615 1398
rect 22686 1396 22692 1398
rect 22756 1396 22762 1460
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
<< via3 >>
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 19748 6156 19812 6220
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 19564 5748 19628 5812
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 22140 5612 22204 5676
rect 22692 5612 22756 5676
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 17908 4116 17972 4180
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 19748 2484 19812 2548
rect 22140 2348 22204 2412
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 19564 1940 19628 2004
rect 17908 1804 17972 1868
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 22692 1396 22756 1460
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
<< metal4 >>
rect 3911 6016 4231 6576
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 3911 1040 4231 1600
rect 6878 6560 7198 6576
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 6878 2208 7198 3232
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 6016 10165 6576
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 12812 6560 13132 6576
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12812 2208 13132 3232
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 6016 16099 6576
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 18746 6560 19066 6576
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 19747 6220 19813 6221
rect 19747 6156 19748 6220
rect 19812 6156 19813 6220
rect 19747 6155 19813 6156
rect 19563 5812 19629 5813
rect 19563 5748 19564 5812
rect 19628 5748 19629 5812
rect 19563 5747 19629 5748
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 17907 4180 17973 4181
rect 17907 4116 17908 4180
rect 17972 4116 17973 4180
rect 17907 4115 17973 4116
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 15779 1664 16099 2688
rect 17910 1869 17970 4115
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18746 2208 19066 3232
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 17907 1868 17973 1869
rect 17907 1804 17908 1868
rect 17972 1804 17973 1868
rect 17907 1803 17973 1804
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 18746 1120 19066 2144
rect 19566 2005 19626 5747
rect 19750 2549 19810 6155
rect 21713 6016 22033 6576
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 24680 6560 25000 6576
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 22139 5676 22205 5677
rect 22139 5612 22140 5676
rect 22204 5612 22205 5676
rect 22139 5611 22205 5612
rect 22691 5676 22757 5677
rect 22691 5612 22692 5676
rect 22756 5612 22757 5676
rect 22691 5611 22757 5612
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 19747 2548 19813 2549
rect 19747 2484 19748 2548
rect 19812 2484 19813 2548
rect 19747 2483 19813 2484
rect 19563 2004 19629 2005
rect 19563 1940 19564 2004
rect 19628 1940 19629 2004
rect 19563 1939 19629 1940
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 1664 22033 2688
rect 22142 2413 22202 5611
rect 22139 2412 22205 2413
rect 22139 2348 22140 2412
rect 22204 2348 22205 2412
rect 22139 2347 22205 2348
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 21713 1040 22033 1600
rect 22694 1461 22754 5611
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 22691 1460 22757 1461
rect 22691 1396 22692 1460
rect 22756 1396 22757 1460
rect 22691 1395 22757 1396
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 8096 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _08_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _09_
timestamp 1688980957
transform -1 0 20332 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _10_
timestamp 1688980957
transform -1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _11_
timestamp 1688980957
transform -1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 6900 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform -1 0 5888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform -1 0 9936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform -1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 2576 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform -1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _28_
timestamp 1688980957
transform -1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _29_
timestamp 1688980957
transform -1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _30_
timestamp 1688980957
transform -1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _31_
timestamp 1688980957
transform -1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _32_
timestamp 1688980957
transform -1 0 12880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 12144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _35_
timestamp 1688980957
transform -1 0 11316 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform -1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform -1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _38_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _39_
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _40_
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _41_
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _42_
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _43_
timestamp 1688980957
transform 1 0 12144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _44_
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _45_
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _46_
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform -1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform -1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform -1 0 19504 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform -1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform -1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform -1 0 21712 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_23 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_49
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54
timestamp 1688980957
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_70
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_76
timestamp 1688980957
transform 1 0 8096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_96
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_100
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_122
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_128
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_148
timestamp 1688980957
transform 1 0 14720 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_154
timestamp 1688980957
transform 1 0 15272 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_158
timestamp 1688980957
transform 1 0 15640 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1688980957
transform 1 0 16376 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_180
timestamp 1688980957
transform 1 0 17664 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_190
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 1688980957
transform 1 0 18952 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_206
timestamp 1688980957
transform 1 0 20056 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_210
timestamp 1688980957
transform 1 0 20424 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_236
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_240
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_244
timestamp 1688980957
transform 1 0 23552 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_62
timestamp 1688980957
transform 1 0 6808 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_70
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_76
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_89
timestamp 1688980957
transform 1 0 9292 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_97
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_102
timestamp 1688980957
transform 1 0 10488 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1688980957
transform 1 0 11224 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_119
timestamp 1688980957
transform 1 0 12052 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_128
timestamp 1688980957
transform 1 0 12880 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_136
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_141
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_200
timestamp 1688980957
transform 1 0 19504 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_212
timestamp 1688980957
transform 1 0 20608 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_253
timestamp 1688980957
transform 1 0 24380 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_68
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_76
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_91
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_95
timestamp 1688980957
transform 1 0 9844 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_103
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_108
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_119
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_123
timestamp 1688980957
transform 1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_131
timestamp 1688980957
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_147
timestamp 1688980957
transform 1 0 14628 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_155
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_159
timestamp 1688980957
transform 1 0 15732 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_171
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_183
timestamp 1688980957
transform 1 0 17940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_206
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_218
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_230
timestamp 1688980957
transform 1 0 22264 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_242
timestamp 1688980957
transform 1 0 23368 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_248
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_187
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_196
timestamp 1688980957
transform 1 0 19136 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_208
timestamp 1688980957
transform 1 0 20240 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_220
timestamp 1688980957
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_245
timestamp 1688980957
transform 1 0 23644 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_10
timestamp 1688980957
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_22
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_202
timestamp 1688980957
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_214
timestamp 1688980957
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_226
timestamp 1688980957
transform 1 0 21896 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_234
timestamp 1688980957
transform 1 0 22632 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_238
timestamp 1688980957
transform 1 0 23000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_242
timestamp 1688980957
transform 1 0 23368 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_17
timestamp 1688980957
transform 1 0 2668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_29
timestamp 1688980957
transform 1 0 3772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_41
timestamp 1688980957
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_200
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_209
timestamp 1688980957
transform 1 0 20332 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_253
timestamp 1688980957
transform 1 0 24380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_25
timestamp 1688980957
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_174
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_186
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_200
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_212
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_220
timestamp 1688980957
transform 1 0 21344 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_23
timestamp 1688980957
transform 1 0 3220 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_40
timestamp 1688980957
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_66
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_85
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_102
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_116
timestamp 1688980957
transform 1 0 11776 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_128
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_140
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_152
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_201
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_209
timestamp 1688980957
transform 1 0 20332 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_216
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_251
timestamp 1688980957
transform 1 0 24196 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_70
timestamp 1688980957
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_128
timestamp 1688980957
transform 1 0 12880 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_154
timestamp 1688980957
transform 1 0 15272 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_194
timestamp 1688980957
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_224
timestamp 1688980957
transform 1 0 21712 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1688980957
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_206
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 14444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 15364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 19504 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 20424 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 21620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 22816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 24288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 6072 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 8464 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 9660 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 10672 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 12052 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 13248 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 10212 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform -1 0 10488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform -1 0 18768 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform -1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform -1 0 19320 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform -1 0 19596 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform -1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  inst_clk_buf
timestamp 1688980957
transform -1 0 18952 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._00_
timestamp 1688980957
transform -1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._01_
timestamp 1688980957
transform 1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._02_
timestamp 1688980957
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._03_
timestamp 1688980957
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._04_
timestamp 1688980957
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._05_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._06_
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._07_
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._08_
timestamp 1688980957
transform -1 0 12604 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._09_
timestamp 1688980957
transform -1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._10_
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._11_
timestamp 1688980957
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._12_
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._13_
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._14_
timestamp 1688980957
transform 1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._15_
timestamp 1688980957
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._16_
timestamp 1688980957
transform -1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._17_
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._18_
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._19_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._20_
timestamp 1688980957
transform -1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._21_
timestamp 1688980957
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._22_
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._23_
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._24_
timestamp 1688980957
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._25_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._26_
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._27_
timestamp 1688980957
transform -1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._28_
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix._29_
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._30_
timestamp 1688980957
transform -1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._31_
timestamp 1688980957
transform -1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform -1 0 18400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform -1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform -1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 23460 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 23644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 21988 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 23000 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform -1 0 23644 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1688980957
transform 1 0 23552 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform -1 0 23092 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 20884 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 22908 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 22356 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 22356 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 22908 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform -1 0 3220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform -1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform -1 0 2668 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform -1 0 2116 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform -1 0 2024 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform -1 0 2576 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform -1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform -1 0 2576 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform -1 0 3680 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform -1 0 3128 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output91 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform -1 0 4508 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform -1 0 3680 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform -1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform -1 0 5336 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform -1 0 4600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform -1 0 5152 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform -1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform -1 0 8280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform -1 0 8832 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform -1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform -1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform -1 0 6440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform -1 0 6716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform -1 0 6992 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform -1 0 6256 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform -1 0 7544 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform -1 0 7360 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 7728 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform -1 0 8832 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 20148 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform -1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform -1 0 10948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform -1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform -1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform -1 0 8740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform -1 0 9936 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform -1 0 11224 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform -1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform -1 0 13524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10._0_
timestamp 1688980957
transform -1 0 14720 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11._0_
timestamp 1688980957
transform -1 0 22356 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform -1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform -1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform -1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform -1 0 20976 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform -1 0 22080 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform -1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform -1 0 23552 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform -1 0 19504 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform -1 0 19688 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform -1 0 12052 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform -1 0 6808 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform -1 0 8096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform -1 0 9292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform -1 0 10488 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform -1 0 11776 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform -1 0 12880 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform -1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform -1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform -1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform -1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform -1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform -1 0 21712 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 24104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform -1 0 24380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 130 592
<< labels >>
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 14094 0 14150 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 15290 0 15346 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 17682 0 17738 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 18878 0 18934 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 21270 0 21326 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 22466 0 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 24858 0 24914 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 3330 0 3386 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 4526 0 4582 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 6918 0 6974 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 8114 0 8170 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 10506 0 10562 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 11702 0 11758 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 20350 7840 20406 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 23110 7840 23166 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 23386 7840 23442 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 23662 7840 23718 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 23938 7840 23994 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 24214 7840 24270 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 24490 7840 24546 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 24766 7840 24822 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 25042 7840 25098 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 25318 7840 25374 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 25594 7840 25650 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 20626 7840 20682 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 20902 7840 20958 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 21178 7840 21234 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 21454 7840 21510 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 21730 7840 21786 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 22006 7840 22062 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 22282 7840 22338 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 22558 7840 22614 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 22834 7840 22890 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 202 7840 258 8000 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 478 7840 534 8000 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 754 7840 810 8000 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 1030 7840 1086 8000 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 1306 7840 1362 8000 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 1582 7840 1638 8000 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 1858 7840 1914 8000 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 2134 7840 2190 8000 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 2410 7840 2466 8000 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 2686 7840 2742 8000 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 2962 7840 3018 8000 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 3238 7840 3294 8000 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 3514 7840 3570 8000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 3790 7840 3846 8000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 4066 7840 4122 8000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 4342 7840 4398 8000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 4618 7840 4674 8000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 4894 7840 4950 8000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 5170 7840 5226 8000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 5446 7840 5502 8000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 5722 7840 5778 8000 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 8482 7840 8538 8000 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 8758 7840 8814 8000 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 9034 7840 9090 8000 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 9310 7840 9366 8000 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 9586 7840 9642 8000 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 9862 7840 9918 8000 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 5998 7840 6054 8000 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 6274 7840 6330 8000 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 6550 7840 6606 8000 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 6826 7840 6882 8000 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 7102 7840 7158 8000 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 7378 7840 7434 8000 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 7654 7840 7710 8000 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 7930 7840 7986 8000 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 8206 7840 8262 8000 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 10138 7840 10194 8000 0 FreeSans 224 90 0 0 S1END[0]
port 76 nsew signal input
flabel metal2 s 10414 7840 10470 8000 0 FreeSans 224 90 0 0 S1END[1]
port 77 nsew signal input
flabel metal2 s 10690 7840 10746 8000 0 FreeSans 224 90 0 0 S1END[2]
port 78 nsew signal input
flabel metal2 s 10966 7840 11022 8000 0 FreeSans 224 90 0 0 S1END[3]
port 79 nsew signal input
flabel metal2 s 11242 7840 11298 8000 0 FreeSans 224 90 0 0 S2END[0]
port 80 nsew signal input
flabel metal2 s 11518 7840 11574 8000 0 FreeSans 224 90 0 0 S2END[1]
port 81 nsew signal input
flabel metal2 s 11794 7840 11850 8000 0 FreeSans 224 90 0 0 S2END[2]
port 82 nsew signal input
flabel metal2 s 12070 7840 12126 8000 0 FreeSans 224 90 0 0 S2END[3]
port 83 nsew signal input
flabel metal2 s 12346 7840 12402 8000 0 FreeSans 224 90 0 0 S2END[4]
port 84 nsew signal input
flabel metal2 s 12622 7840 12678 8000 0 FreeSans 224 90 0 0 S2END[5]
port 85 nsew signal input
flabel metal2 s 12898 7840 12954 8000 0 FreeSans 224 90 0 0 S2END[6]
port 86 nsew signal input
flabel metal2 s 13174 7840 13230 8000 0 FreeSans 224 90 0 0 S2END[7]
port 87 nsew signal input
flabel metal2 s 13450 7840 13506 8000 0 FreeSans 224 90 0 0 S2MID[0]
port 88 nsew signal input
flabel metal2 s 13726 7840 13782 8000 0 FreeSans 224 90 0 0 S2MID[1]
port 89 nsew signal input
flabel metal2 s 14002 7840 14058 8000 0 FreeSans 224 90 0 0 S2MID[2]
port 90 nsew signal input
flabel metal2 s 14278 7840 14334 8000 0 FreeSans 224 90 0 0 S2MID[3]
port 91 nsew signal input
flabel metal2 s 14554 7840 14610 8000 0 FreeSans 224 90 0 0 S2MID[4]
port 92 nsew signal input
flabel metal2 s 14830 7840 14886 8000 0 FreeSans 224 90 0 0 S2MID[5]
port 93 nsew signal input
flabel metal2 s 15106 7840 15162 8000 0 FreeSans 224 90 0 0 S2MID[6]
port 94 nsew signal input
flabel metal2 s 15382 7840 15438 8000 0 FreeSans 224 90 0 0 S2MID[7]
port 95 nsew signal input
flabel metal2 s 15658 7840 15714 8000 0 FreeSans 224 90 0 0 S4END[0]
port 96 nsew signal input
flabel metal2 s 18418 7840 18474 8000 0 FreeSans 224 90 0 0 S4END[10]
port 97 nsew signal input
flabel metal2 s 18694 7840 18750 8000 0 FreeSans 224 90 0 0 S4END[11]
port 98 nsew signal input
flabel metal2 s 18970 7840 19026 8000 0 FreeSans 224 90 0 0 S4END[12]
port 99 nsew signal input
flabel metal2 s 19246 7840 19302 8000 0 FreeSans 224 90 0 0 S4END[13]
port 100 nsew signal input
flabel metal2 s 19522 7840 19578 8000 0 FreeSans 224 90 0 0 S4END[14]
port 101 nsew signal input
flabel metal2 s 19798 7840 19854 8000 0 FreeSans 224 90 0 0 S4END[15]
port 102 nsew signal input
flabel metal2 s 15934 7840 15990 8000 0 FreeSans 224 90 0 0 S4END[1]
port 103 nsew signal input
flabel metal2 s 16210 7840 16266 8000 0 FreeSans 224 90 0 0 S4END[2]
port 104 nsew signal input
flabel metal2 s 16486 7840 16542 8000 0 FreeSans 224 90 0 0 S4END[3]
port 105 nsew signal input
flabel metal2 s 16762 7840 16818 8000 0 FreeSans 224 90 0 0 S4END[4]
port 106 nsew signal input
flabel metal2 s 17038 7840 17094 8000 0 FreeSans 224 90 0 0 S4END[5]
port 107 nsew signal input
flabel metal2 s 17314 7840 17370 8000 0 FreeSans 224 90 0 0 S4END[6]
port 108 nsew signal input
flabel metal2 s 17590 7840 17646 8000 0 FreeSans 224 90 0 0 S4END[7]
port 109 nsew signal input
flabel metal2 s 17866 7840 17922 8000 0 FreeSans 224 90 0 0 S4END[8]
port 110 nsew signal input
flabel metal2 s 18142 7840 18198 8000 0 FreeSans 224 90 0 0 S4END[9]
port 111 nsew signal input
flabel metal2 s 938 0 994 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 20074 7840 20130 8000 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6878 1040 7198 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9845 1040 10165 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15779 1040 16099 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21713 1040 22033 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 13052 6528 13052 6528 0 VGND
rlabel metal1 12972 5984 12972 5984 0 VPWR
rlabel metal2 2215 68 2215 68 0 FrameStrobe[0]
rlabel metal2 14175 68 14175 68 0 FrameStrobe[10]
rlabel metal2 15371 68 15371 68 0 FrameStrobe[11]
rlabel metal2 16514 704 16514 704 0 FrameStrobe[12]
rlabel metal2 17710 704 17710 704 0 FrameStrobe[13]
rlabel metal2 18906 143 18906 143 0 FrameStrobe[14]
rlabel metal2 20102 704 20102 704 0 FrameStrobe[15]
rlabel metal2 21351 68 21351 68 0 FrameStrobe[16]
rlabel metal2 22547 68 22547 68 0 FrameStrobe[17]
rlabel metal2 23690 143 23690 143 0 FrameStrobe[18]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[19]
rlabel metal2 3358 704 3358 704 0 FrameStrobe[1]
rlabel metal2 4607 68 4607 68 0 FrameStrobe[2]
rlabel metal2 5750 704 5750 704 0 FrameStrobe[3]
rlabel metal2 7137 68 7137 68 0 FrameStrobe[4]
rlabel metal2 8142 704 8142 704 0 FrameStrobe[5]
rlabel metal2 9338 704 9338 704 0 FrameStrobe[6]
rlabel metal2 10481 68 10481 68 0 FrameStrobe[7]
rlabel metal2 11730 704 11730 704 0 FrameStrobe[8]
rlabel metal2 12827 68 12827 68 0 FrameStrobe[9]
rlabel metal2 20378 7473 20378 7473 0 FrameStrobe_O[0]
rlabel metal2 23138 6912 23138 6912 0 FrameStrobe_O[10]
rlabel metal2 23414 6997 23414 6997 0 FrameStrobe_O[11]
rlabel metal2 23690 6368 23690 6368 0 FrameStrobe_O[12]
rlabel metal1 22494 5134 22494 5134 0 FrameStrobe_O[13]
rlabel metal1 23598 4046 23598 4046 0 FrameStrobe_O[14]
rlabel metal1 23874 4998 23874 4998 0 FrameStrobe_O[15]
rlabel metal1 24288 4046 24288 4046 0 FrameStrobe_O[16]
rlabel metal1 23874 5134 23874 5134 0 FrameStrobe_O[17]
rlabel metal1 24748 3706 24748 3706 0 FrameStrobe_O[18]
rlabel metal1 23920 5814 23920 5814 0 FrameStrobe_O[19]
rlabel metal2 20654 6878 20654 6878 0 FrameStrobe_O[1]
rlabel metal2 21029 7956 21029 7956 0 FrameStrobe_O[2]
rlabel metal2 21305 7956 21305 7956 0 FrameStrobe_O[3]
rlabel metal2 21482 7864 21482 7864 0 FrameStrobe_O[4]
rlabel metal2 21857 7956 21857 7956 0 FrameStrobe_O[5]
rlabel metal2 22034 7065 22034 7065 0 FrameStrobe_O[6]
rlabel metal2 22310 6912 22310 6912 0 FrameStrobe_O[7]
rlabel metal2 22586 6368 22586 6368 0 FrameStrobe_O[8]
rlabel metal2 22862 6912 22862 6912 0 FrameStrobe_O[9]
rlabel metal1 3404 4794 3404 4794 0 Inst_S_term_RAM_IO_switch_matrix.N1BEG0
rlabel metal1 2806 4624 2806 4624 0 Inst_S_term_RAM_IO_switch_matrix.N1BEG1
rlabel metal1 1978 3502 1978 3502 0 Inst_S_term_RAM_IO_switch_matrix.N1BEG2
rlabel metal1 1702 3536 1702 3536 0 Inst_S_term_RAM_IO_switch_matrix.N1BEG3
rlabel metal1 15410 6222 15410 6222 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG0
rlabel metal1 14582 6324 14582 6324 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG1
rlabel metal1 14030 6290 14030 6290 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG2
rlabel via1 12838 6294 12838 6294 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG3
rlabel metal1 12696 5678 12696 5678 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG4
rlabel metal1 12374 5712 12374 5712 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG5
rlabel metal1 11132 6290 11132 6290 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG6
rlabel metal1 11178 5202 11178 5202 0 Inst_S_term_RAM_IO_switch_matrix.N2BEG7
rlabel metal1 9614 5712 9614 5712 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb0
rlabel metal1 8372 5202 8372 5202 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb1
rlabel metal1 6394 4998 6394 4998 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb2
rlabel metal1 4554 4794 4554 4794 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb3
rlabel metal1 4830 5202 4830 5202 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb4
rlabel metal1 5474 5202 5474 5202 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb5
rlabel metal1 4738 7446 4738 7446 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb6
rlabel metal1 6210 5202 6210 5202 0 Inst_S_term_RAM_IO_switch_matrix.N2BEGb7
rlabel metal1 20700 5678 20700 5678 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 20194 5202 20194 5202 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG1
rlabel metal1 17756 6290 17756 6290 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG10
rlabel metal1 17204 6290 17204 6290 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG11
rlabel metal1 15594 5712 15594 5712 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG12
rlabel metal1 9338 5168 9338 5168 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG13
rlabel metal2 9614 5678 9614 5678 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG14
rlabel metal1 9936 5202 9936 5202 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG15
rlabel metal1 19780 5678 19780 5678 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 19550 5678 19550 5678 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG3
rlabel metal2 8050 7072 8050 7072 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG4
rlabel metal1 7682 7650 7682 7650 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG5
rlabel metal2 7774 6494 7774 6494 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG6
rlabel metal1 5658 5712 5658 5712 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG7
rlabel metal2 8786 6715 8786 6715 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG8
rlabel metal1 8878 5134 8878 5134 0 Inst_S_term_RAM_IO_switch_matrix.N4BEG9
rlabel metal2 230 7201 230 7201 0 N1BEG[0]
rlabel metal2 506 7150 506 7150 0 N1BEG[1]
rlabel metal2 782 6334 782 6334 0 N1BEG[2]
rlabel metal2 1058 5926 1058 5926 0 N1BEG[3]
rlabel metal2 1334 6368 1334 6368 0 N2BEG[0]
rlabel metal2 1610 6606 1610 6606 0 N2BEG[1]
rlabel metal2 1886 6640 1886 6640 0 N2BEG[2]
rlabel metal2 2162 6912 2162 6912 0 N2BEG[3]
rlabel metal2 2385 7956 2385 7956 0 N2BEG[4]
rlabel metal2 2714 6912 2714 6912 0 N2BEG[5]
rlabel metal1 2668 6426 2668 6426 0 N2BEG[6]
rlabel metal2 3266 6912 3266 6912 0 N2BEG[7]
rlabel metal1 3036 6222 3036 6222 0 N2BEGb[0]
rlabel metal1 3542 5338 3542 5338 0 N2BEGb[1]
rlabel metal2 3995 7956 3995 7956 0 N2BEGb[2]
rlabel metal1 3772 6426 3772 6426 0 N2BEGb[3]
rlabel metal2 4600 5338 4600 5338 0 N2BEGb[4]
rlabel metal2 4922 6912 4922 6912 0 N2BEGb[5]
rlabel metal1 4370 6392 4370 6392 0 N2BEGb[6]
rlabel metal1 5106 6426 5106 6426 0 N2BEGb[7]
rlabel metal1 5612 6426 5612 6426 0 N4BEG[0]
rlabel metal1 8280 6426 8280 6426 0 N4BEG[10]
rlabel metal2 8602 7191 8602 7191 0 N4BEG[11]
rlabel metal1 9108 5882 9108 5882 0 N4BEG[12]
rlabel metal2 9338 7184 9338 7184 0 N4BEG[13]
rlabel metal2 9614 7150 9614 7150 0 N4BEG[14]
rlabel metal2 9890 7184 9890 7184 0 N4BEG[15]
rlabel metal2 6026 6912 6026 6912 0 N4BEG[1]
rlabel metal1 6394 6426 6394 6426 0 N4BEG[2]
rlabel metal2 6578 6912 6578 6912 0 N4BEG[3]
rlabel metal1 6394 6086 6394 6086 0 N4BEG[4]
rlabel metal2 7130 7337 7130 7337 0 N4BEG[5]
rlabel metal1 7268 6426 7268 6426 0 N4BEG[6]
rlabel metal2 7590 7191 7590 7191 0 N4BEG[7]
rlabel metal2 7958 6912 7958 6912 0 N4BEG[8]
rlabel metal2 8234 6912 8234 6912 0 N4BEG[9]
rlabel metal2 10166 7677 10166 7677 0 S1END[0]
rlabel metal2 10442 6810 10442 6810 0 S1END[1]
rlabel metal2 10718 7269 10718 7269 0 S1END[2]
rlabel metal2 10994 6810 10994 6810 0 S1END[3]
rlabel metal2 11270 7269 11270 7269 0 S2END[0]
rlabel metal2 11546 6810 11546 6810 0 S2END[1]
rlabel metal2 11822 6810 11822 6810 0 S2END[2]
rlabel metal2 12098 6810 12098 6810 0 S2END[3]
rlabel metal2 12374 7626 12374 7626 0 S2END[4]
rlabel metal1 12282 6324 12282 6324 0 S2END[5]
rlabel metal2 13025 7956 13025 7956 0 S2END[6]
rlabel metal2 13202 7864 13202 7864 0 S2END[7]
rlabel metal2 13478 7116 13478 7116 0 S2MID[0]
rlabel metal2 13701 7956 13701 7956 0 S2MID[1]
rlabel metal2 14129 7956 14129 7956 0 S2MID[2]
rlabel metal2 14306 6810 14306 6810 0 S2MID[3]
rlabel metal2 14582 6810 14582 6810 0 S2MID[4]
rlabel metal2 14858 7388 14858 7388 0 S2MID[5]
rlabel metal2 15134 7184 15134 7184 0 S2MID[6]
rlabel metal2 15410 6776 15410 6776 0 S2MID[7]
rlabel metal2 15686 7405 15686 7405 0 S4END[0]
rlabel metal2 18499 7956 18499 7956 0 S4END[10]
rlabel metal2 18722 7286 18722 7286 0 S4END[11]
rlabel metal2 19097 7956 19097 7956 0 S4END[12]
rlabel metal2 19274 6725 19274 6725 0 S4END[13]
rlabel metal2 19550 7150 19550 7150 0 S4END[14]
rlabel metal2 19826 7269 19826 7269 0 S4END[15]
rlabel metal2 15962 7388 15962 7388 0 S4END[1]
rlabel metal2 16238 6776 16238 6776 0 S4END[2]
rlabel metal2 16514 7473 16514 7473 0 S4END[3]
rlabel metal2 16790 7388 16790 7388 0 S4END[4]
rlabel metal2 17066 7286 17066 7286 0 S4END[5]
rlabel metal2 17342 7184 17342 7184 0 S4END[6]
rlabel metal2 17618 7609 17618 7609 0 S4END[7]
rlabel metal2 17841 7956 17841 7956 0 S4END[8]
rlabel metal2 18170 7320 18170 7320 0 S4END[9]
rlabel metal2 966 704 966 704 0 UserCLK
rlabel metal2 20102 7184 20102 7184 0 UserCLKo
rlabel metal2 2438 1700 2438 1700 0 net1
rlabel metal1 23552 1326 23552 1326 0 net10
rlabel metal1 9108 6358 9108 6358 0 net100
rlabel metal1 9338 5712 9338 5712 0 net101
rlabel metal1 9246 5338 9246 5338 0 net102
rlabel metal1 10212 5066 10212 5066 0 net103
rlabel metal2 10166 5423 10166 5423 0 net104
rlabel metal2 6302 5355 6302 5355 0 net105
rlabel metal1 6791 6290 6791 6290 0 net106
rlabel metal1 6854 5576 6854 5576 0 net107
rlabel metal1 6118 6324 6118 6324 0 net108
rlabel metal1 7360 5338 7360 5338 0 net109
rlabel metal1 24288 1190 24288 1190 0 net11
rlabel metal1 7544 5338 7544 5338 0 net110
rlabel metal1 6371 5814 6371 5814 0 net111
rlabel metal2 7866 5474 7866 5474 0 net112
rlabel metal2 8694 5474 8694 5474 0 net113
rlabel metal1 18722 1190 18722 1190 0 net114
rlabel metal2 3634 2108 3634 2108 0 net12
rlabel metal2 4830 1088 4830 1088 0 net13
rlabel metal1 6210 1326 6210 1326 0 net14
rlabel metal1 7268 1326 7268 1326 0 net15
rlabel metal1 8464 1326 8464 1326 0 net16
rlabel metal1 9660 1326 9660 1326 0 net17
rlabel metal1 10994 1292 10994 1292 0 net18
rlabel metal1 12052 1326 12052 1326 0 net19
rlabel metal1 14444 1326 14444 1326 0 net2
rlabel metal1 13248 1326 13248 1326 0 net20
rlabel metal2 10258 4658 10258 4658 0 net21
rlabel metal2 5014 5712 5014 5712 0 net22
rlabel metal1 3358 4556 3358 4556 0 net23
rlabel metal1 3266 4624 3266 4624 0 net24
rlabel metal1 6578 5134 6578 5134 0 net25
rlabel metal1 11040 5678 11040 5678 0 net26
rlabel metal1 6670 5202 6670 5202 0 net27
rlabel metal1 6854 6120 6854 6120 0 net28
rlabel metal2 5934 6018 5934 6018 0 net29
rlabel metal1 15594 1258 15594 1258 0 net3
rlabel metal1 6854 5236 6854 5236 0 net30
rlabel metal1 8602 5236 8602 5236 0 net31
rlabel metal1 10166 5644 10166 5644 0 net32
rlabel metal1 11316 5678 11316 5678 0 net33
rlabel metal1 11362 6256 11362 6256 0 net34
rlabel metal1 11822 6358 11822 6358 0 net35
rlabel metal1 14214 5542 14214 5542 0 net36
rlabel metal1 13892 5882 13892 5882 0 net37
rlabel metal1 14306 6222 14306 6222 0 net38
rlabel metal1 15134 6324 15134 6324 0 net39
rlabel metal1 16882 1258 16882 1258 0 net4
rlabel metal2 15686 6086 15686 6086 0 net40
rlabel metal1 9844 5678 9844 5678 0 net41
rlabel metal1 18676 5338 18676 5338 0 net42
rlabel metal1 19458 6324 19458 6324 0 net43
rlabel metal1 19596 5066 19596 5066 0 net44
rlabel metal1 19780 5338 19780 5338 0 net45
rlabel metal1 20286 5712 20286 5712 0 net46
rlabel metal1 21068 4998 21068 4998 0 net47
rlabel metal2 16514 6086 16514 6086 0 net48
rlabel metal1 16928 5882 16928 5882 0 net49
rlabel metal1 18032 1190 18032 1190 0 net5
rlabel metal1 16146 5712 16146 5712 0 net50
rlabel metal1 17434 6324 17434 6324 0 net51
rlabel metal1 17986 6256 17986 6256 0 net52
rlabel metal1 17526 5746 17526 5746 0 net53
rlabel metal1 17802 5644 17802 5644 0 net54
rlabel metal1 18078 5712 18078 5712 0 net55
rlabel metal1 18400 5678 18400 5678 0 net56
rlabel metal1 1610 1224 1610 1224 0 net57
rlabel metal1 20424 2618 20424 2618 0 net58
rlabel metal1 19826 2550 19826 2550 0 net59
rlabel metal1 19320 1190 19320 1190 0 net6
rlabel metal1 23368 3638 23368 3638 0 net60
rlabel metal1 23598 3706 23598 3706 0 net61
rlabel metal1 19458 4216 19458 4216 0 net62
rlabel metal1 21390 5032 21390 5032 0 net63
rlabel metal1 23782 5270 23782 5270 0 net64
rlabel metal1 23644 4114 23644 4114 0 net65
rlabel metal1 23414 2822 23414 2822 0 net66
rlabel metal1 23966 2618 23966 2618 0 net67
rlabel metal1 21804 5338 21804 5338 0 net68
rlabel metal1 20654 3978 20654 3978 0 net69
rlabel metal1 20562 1190 20562 1190 0 net7
rlabel metal1 11960 2618 11960 2618 0 net70
rlabel metal2 7314 2125 7314 2125 0 net71
rlabel via2 8602 2533 8602 2533 0 net72
rlabel metal1 9798 2312 9798 2312 0 net73
rlabel metal2 10994 2057 10994 2057 0 net74
rlabel metal2 12374 2329 12374 2329 0 net75
rlabel metal2 13478 3570 13478 3570 0 net76
rlabel metal2 14582 1853 14582 1853 0 net77
rlabel metal1 3404 5270 3404 5270 0 net78
rlabel metal1 2438 4794 2438 4794 0 net79
rlabel metal1 21620 1190 21620 1190 0 net8
rlabel metal1 2024 3706 2024 3706 0 net80
rlabel metal2 1518 3910 1518 3910 0 net81
rlabel via2 1794 4539 1794 4539 0 net82
rlabel via2 2530 5219 2530 5219 0 net83
rlabel metal1 1978 4556 1978 4556 0 net84
rlabel metal1 1886 5746 1886 5746 0 net85
rlabel metal1 2944 5610 2944 5610 0 net86
rlabel metal1 2990 5712 2990 5712 0 net87
rlabel metal1 2668 6358 2668 6358 0 net88
rlabel metal1 4048 5678 4048 5678 0 net89
rlabel metal1 23138 1190 23138 1190 0 net9
rlabel metal1 2990 6324 2990 6324 0 net90
rlabel metal2 6762 4896 6762 4896 0 net91
rlabel metal1 4370 5576 4370 5576 0 net92
rlabel metal1 3772 4998 3772 4998 0 net93
rlabel metal1 4784 5270 4784 5270 0 net94
rlabel metal2 5198 5474 5198 5474 0 net95
rlabel metal1 4508 5882 4508 5882 0 net96
rlabel metal2 5842 5814 5842 5814 0 net97
rlabel metal1 5796 6358 5796 6358 0 net98
rlabel metal1 8234 6358 8234 6358 0 net99
rlabel metal1 19044 1938 19044 1938 0 strobe_inbuf_0.X
rlabel metal1 19274 3162 19274 3162 0 strobe_inbuf_1.X
rlabel metal1 14812 1530 14812 1530 0 strobe_inbuf_10.X
rlabel metal1 22402 4148 22402 4148 0 strobe_inbuf_11.X
rlabel metal2 18630 4250 18630 4250 0 strobe_inbuf_12.X
rlabel metal1 18446 3162 18446 3162 0 strobe_inbuf_13.X
rlabel metal1 19642 4794 19642 4794 0 strobe_inbuf_14.X
rlabel metal1 21206 5338 21206 5338 0 strobe_inbuf_15.X
rlabel metal2 22218 4284 22218 4284 0 strobe_inbuf_16.X
rlabel metal1 24334 4148 24334 4148 0 strobe_inbuf_17.X
rlabel metal1 23828 1530 23828 1530 0 strobe_inbuf_18.X
rlabel metal1 23920 2890 23920 2890 0 strobe_inbuf_19.X
rlabel metal1 11270 1190 11270 1190 0 strobe_inbuf_2.X
rlabel metal2 6578 1734 6578 1734 0 strobe_inbuf_3.X
rlabel metal1 7682 1530 7682 1530 0 strobe_inbuf_4.X
rlabel metal1 8878 1530 8878 1530 0 strobe_inbuf_5.X
rlabel metal1 10074 1530 10074 1530 0 strobe_inbuf_6.X
rlabel metal1 11362 1530 11362 1530 0 strobe_inbuf_7.X
rlabel metal1 12466 1530 12466 1530 0 strobe_inbuf_8.X
rlabel metal1 13662 1190 13662 1190 0 strobe_inbuf_9.X
rlabel metal1 19642 2074 19642 2074 0 strobe_outbuf_0.X
rlabel metal1 19872 3706 19872 3706 0 strobe_outbuf_1.X
rlabel metal1 15318 2074 15318 2074 0 strobe_outbuf_10.X
rlabel metal1 22678 3502 22678 3502 0 strobe_outbuf_11.X
rlabel metal1 23000 3502 23000 3502 0 strobe_outbuf_12.X
rlabel metal1 19044 3706 19044 3706 0 strobe_outbuf_13.X
rlabel metal1 20470 5168 20470 5168 0 strobe_outbuf_14.X
rlabel metal2 21666 5984 21666 5984 0 strobe_outbuf_15.X
rlabel metal2 21574 4420 21574 4420 0 strobe_outbuf_16.X
rlabel metal1 24104 3026 24104 3026 0 strobe_outbuf_17.X
rlabel metal1 24288 2074 24288 2074 0 strobe_outbuf_18.X
rlabel metal1 22494 3366 22494 3366 0 strobe_outbuf_19.X
rlabel metal1 11914 2074 11914 2074 0 strobe_outbuf_2.X
rlabel metal2 6762 2244 6762 2244 0 strobe_outbuf_3.X
rlabel metal1 8234 2074 8234 2074 0 strobe_outbuf_4.X
rlabel metal1 9430 2074 9430 2074 0 strobe_outbuf_5.X
rlabel metal1 10626 2074 10626 2074 0 strobe_outbuf_6.X
rlabel metal1 11730 2040 11730 2040 0 strobe_outbuf_7.X
rlabel metal1 13064 2074 13064 2074 0 strobe_outbuf_8.X
rlabel metal1 14214 2074 14214 2074 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 8000
<< end >>
