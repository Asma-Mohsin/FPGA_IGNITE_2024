VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BlockRAM_1KB
  CLASS BLOCK ;
  FOREIGN BlockRAM_1KB ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 446.230 ;
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END C0
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END C3
  PIN C4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END C4
  PIN C5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END C5
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 457.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 566.080 -7.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 454.000 566.080 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 562.980 -11.020 566.080 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.340 -11.020 25.940 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 420.480 179.540 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 421.100 333.140 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 420.480 486.740 457.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 30.030 566.080 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 183.210 566.080 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 336.390 566.080 337.990 ;
    END
    PORT
      LAYER met4 ;
        RECT 537.860 10.640 539.460 435.440 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 452.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 561.280 -3.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 449.200 561.280 452.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.180 -6.220 561.280 452.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -11.020 22.640 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 420.480 176.240 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 420.480 329.840 457.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 420.480 483.440 457.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 26.730 566.080 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 179.910 566.080 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 333.090 566.080 334.690 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.180 10.640 535.780 435.440 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END clk
  PIN rd_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 442.230 438.290 446.230 ;
    END
  END rd_addr[0]
  PIN rd_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 105.440 550.000 106.040 ;
    END
  END rd_addr[1]
  PIN rd_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 98.640 550.000 99.240 ;
    END
  END rd_addr[2]
  PIN rd_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 91.840 550.000 92.440 ;
    END
  END rd_addr[3]
  PIN rd_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END rd_addr[4]
  PIN rd_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END rd_addr[5]
  PIN rd_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END rd_addr[6]
  PIN rd_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END rd_addr[7]
  PIN rd_data[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END rd_data[0]
  PIN rd_data[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END rd_data[10]
  PIN rd_data[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END rd_data[11]
  PIN rd_data[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END rd_data[12]
  PIN rd_data[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END rd_data[13]
  PIN rd_data[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END rd_data[14]
  PIN rd_data[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END rd_data[15]
  PIN rd_data[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END rd_data[16]
  PIN rd_data[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END rd_data[17]
  PIN rd_data[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END rd_data[18]
  PIN rd_data[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END rd_data[19]
  PIN rd_data[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END rd_data[1]
  PIN rd_data[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 280.230 442.230 280.510 446.230 ;
    END
  END rd_data[20]
  PIN rd_data[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 486.310 442.230 486.590 446.230 ;
    END
  END rd_data[21]
  PIN rd_data[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 354.290 442.230 354.570 446.230 ;
    END
  END rd_data[22]
  PIN rd_data[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 231.930 442.230 232.210 446.230 ;
    END
  END rd_data[23]
  PIN rd_data[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 257.690 442.230 257.970 446.230 ;
    END
  END rd_data[24]
  PIN rd_data[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 305.990 442.230 306.270 446.230 ;
    END
  END rd_data[25]
  PIN rd_data[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 502.410 442.230 502.690 446.230 ;
    END
  END rd_data[26]
  PIN rd_data[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 476.650 442.230 476.930 446.230 ;
    END
  END rd_data[27]
  PIN rd_data[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 415.470 442.230 415.750 446.230 ;
    END
  END rd_data[28]
  PIN rd_data[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 546.000 428.440 550.000 429.040 ;
    END
  END rd_data[29]
  PIN rd_data[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END rd_data[2]
  PIN rd_data[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END rd_data[30]
  PIN rd_data[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END rd_data[31]
  PIN rd_data[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END rd_data[7]
  PIN rd_data[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END rd_data[8]
  PIN rd_data[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END rd_data[9]
  PIN wr_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wr_addr[0]
  PIN wr_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END wr_addr[1]
  PIN wr_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END wr_addr[2]
  PIN wr_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END wr_addr[3]
  PIN wr_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END wr_addr[4]
  PIN wr_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END wr_addr[5]
  PIN wr_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wr_addr[6]
  PIN wr_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wr_addr[7]
  PIN wr_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END wr_data[0]
  PIN wr_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END wr_data[10]
  PIN wr_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END wr_data[11]
  PIN wr_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wr_data[15]
  PIN wr_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wr_data[19]
  PIN wr_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END wr_data[1]
  PIN wr_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wr_data[29]
  PIN wr_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END wr_data[2]
  PIN wr_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END wr_data[31]
  PIN wr_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END wr_data[7]
  PIN wr_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END wr_data[8]
  PIN wr_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END wr_data[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 544.370 435.285 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 435.285 ;
      LAYER met1 ;
        RECT 0.070 9.560 544.180 440.260 ;
      LAYER met2 ;
        RECT 0.100 441.950 231.650 442.410 ;
        RECT 232.490 441.950 257.410 442.410 ;
        RECT 258.250 441.950 279.950 442.410 ;
        RECT 280.790 441.950 305.710 442.410 ;
        RECT 306.550 441.950 354.010 442.410 ;
        RECT 354.850 441.950 415.190 442.410 ;
        RECT 416.030 441.950 437.730 442.410 ;
        RECT 438.570 441.950 476.370 442.410 ;
        RECT 477.210 441.950 486.030 442.410 ;
        RECT 486.870 441.950 502.130 442.410 ;
        RECT 502.970 441.950 542.250 442.410 ;
        RECT 0.100 4.280 542.250 441.950 ;
        RECT 0.100 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 25.570 4.280 ;
        RECT 26.410 4.000 115.730 4.280 ;
        RECT 116.570 4.000 450.610 4.280 ;
        RECT 451.450 4.000 453.830 4.280 ;
        RECT 454.670 4.000 457.050 4.280 ;
        RECT 457.890 4.000 460.270 4.280 ;
        RECT 461.110 4.000 542.250 4.280 ;
      LAYER met3 ;
        RECT 1.445 432.840 546.000 441.145 ;
        RECT 4.400 431.440 546.000 432.840 ;
        RECT 1.445 429.440 546.000 431.440 ;
        RECT 4.400 428.040 545.600 429.440 ;
        RECT 1.445 426.040 546.000 428.040 ;
        RECT 4.400 424.640 546.000 426.040 ;
        RECT 1.445 422.640 546.000 424.640 ;
        RECT 4.400 421.240 546.000 422.640 ;
        RECT 1.445 415.840 546.000 421.240 ;
        RECT 4.400 414.440 546.000 415.840 ;
        RECT 1.445 412.440 546.000 414.440 ;
        RECT 4.400 411.040 546.000 412.440 ;
        RECT 1.445 409.040 546.000 411.040 ;
        RECT 4.400 407.640 546.000 409.040 ;
        RECT 1.445 402.240 546.000 407.640 ;
        RECT 4.400 400.840 546.000 402.240 ;
        RECT 1.445 388.640 546.000 400.840 ;
        RECT 4.400 387.240 546.000 388.640 ;
        RECT 1.445 385.240 546.000 387.240 ;
        RECT 4.400 383.840 546.000 385.240 ;
        RECT 1.445 381.840 546.000 383.840 ;
        RECT 4.400 380.440 546.000 381.840 ;
        RECT 1.445 375.040 546.000 380.440 ;
        RECT 4.400 373.640 546.000 375.040 ;
        RECT 1.445 371.640 546.000 373.640 ;
        RECT 4.400 370.240 546.000 371.640 ;
        RECT 1.445 361.440 546.000 370.240 ;
        RECT 4.400 360.040 546.000 361.440 ;
        RECT 1.445 347.840 546.000 360.040 ;
        RECT 4.400 346.440 546.000 347.840 ;
        RECT 1.445 344.440 546.000 346.440 ;
        RECT 4.400 343.040 546.000 344.440 ;
        RECT 1.445 341.040 546.000 343.040 ;
        RECT 4.400 339.640 546.000 341.040 ;
        RECT 1.445 330.840 546.000 339.640 ;
        RECT 4.400 329.440 546.000 330.840 ;
        RECT 1.445 327.440 546.000 329.440 ;
        RECT 4.400 326.040 546.000 327.440 ;
        RECT 1.445 324.040 546.000 326.040 ;
        RECT 4.400 322.640 546.000 324.040 ;
        RECT 1.445 293.440 546.000 322.640 ;
        RECT 4.400 292.040 546.000 293.440 ;
        RECT 1.445 290.040 546.000 292.040 ;
        RECT 4.400 288.640 546.000 290.040 ;
        RECT 1.445 283.240 546.000 288.640 ;
        RECT 4.400 281.840 546.000 283.240 ;
        RECT 1.445 276.440 546.000 281.840 ;
        RECT 4.400 275.040 546.000 276.440 ;
        RECT 1.445 269.640 546.000 275.040 ;
        RECT 4.400 268.240 546.000 269.640 ;
        RECT 1.445 259.440 546.000 268.240 ;
        RECT 4.400 258.040 546.000 259.440 ;
        RECT 1.445 232.240 546.000 258.040 ;
        RECT 4.400 230.840 546.000 232.240 ;
        RECT 1.445 228.840 546.000 230.840 ;
        RECT 4.400 227.440 546.000 228.840 ;
        RECT 1.445 208.440 546.000 227.440 ;
        RECT 4.400 207.040 546.000 208.440 ;
        RECT 1.445 205.040 546.000 207.040 ;
        RECT 4.400 203.640 546.000 205.040 ;
        RECT 1.445 201.640 546.000 203.640 ;
        RECT 4.400 200.240 546.000 201.640 ;
        RECT 1.445 194.840 546.000 200.240 ;
        RECT 4.400 193.440 546.000 194.840 ;
        RECT 1.445 188.040 546.000 193.440 ;
        RECT 4.400 186.640 546.000 188.040 ;
        RECT 1.445 184.640 546.000 186.640 ;
        RECT 4.400 183.240 546.000 184.640 ;
        RECT 1.445 181.240 546.000 183.240 ;
        RECT 4.400 179.840 546.000 181.240 ;
        RECT 1.445 177.840 546.000 179.840 ;
        RECT 4.400 176.440 546.000 177.840 ;
        RECT 1.445 174.440 546.000 176.440 ;
        RECT 4.400 173.040 546.000 174.440 ;
        RECT 1.445 171.040 546.000 173.040 ;
        RECT 4.400 169.640 546.000 171.040 ;
        RECT 1.445 167.640 546.000 169.640 ;
        RECT 4.400 166.240 546.000 167.640 ;
        RECT 1.445 164.240 546.000 166.240 ;
        RECT 4.400 162.840 546.000 164.240 ;
        RECT 1.445 160.840 546.000 162.840 ;
        RECT 4.400 159.440 546.000 160.840 ;
        RECT 1.445 157.440 546.000 159.440 ;
        RECT 4.400 156.040 546.000 157.440 ;
        RECT 1.445 154.040 546.000 156.040 ;
        RECT 4.400 152.640 546.000 154.040 ;
        RECT 1.445 150.640 546.000 152.640 ;
        RECT 4.400 149.240 546.000 150.640 ;
        RECT 1.445 147.240 546.000 149.240 ;
        RECT 4.400 145.840 546.000 147.240 ;
        RECT 1.445 143.840 546.000 145.840 ;
        RECT 4.400 142.440 546.000 143.840 ;
        RECT 1.445 140.440 546.000 142.440 ;
        RECT 4.400 139.040 546.000 140.440 ;
        RECT 1.445 133.640 546.000 139.040 ;
        RECT 4.400 132.240 546.000 133.640 ;
        RECT 1.445 120.040 546.000 132.240 ;
        RECT 4.400 118.640 546.000 120.040 ;
        RECT 1.445 113.240 546.000 118.640 ;
        RECT 4.400 111.840 546.000 113.240 ;
        RECT 1.445 109.840 546.000 111.840 ;
        RECT 4.400 108.440 546.000 109.840 ;
        RECT 1.445 106.440 546.000 108.440 ;
        RECT 4.400 105.040 545.600 106.440 ;
        RECT 1.445 103.040 546.000 105.040 ;
        RECT 4.400 101.640 546.000 103.040 ;
        RECT 1.445 99.640 546.000 101.640 ;
        RECT 4.400 98.240 545.600 99.640 ;
        RECT 1.445 96.240 546.000 98.240 ;
        RECT 4.400 94.840 546.000 96.240 ;
        RECT 1.445 92.840 546.000 94.840 ;
        RECT 4.400 91.440 545.600 92.840 ;
        RECT 1.445 89.440 546.000 91.440 ;
        RECT 4.400 88.040 546.000 89.440 ;
        RECT 1.445 55.440 546.000 88.040 ;
        RECT 4.400 54.040 546.000 55.440 ;
        RECT 1.445 52.040 546.000 54.040 ;
        RECT 4.400 50.640 546.000 52.040 ;
        RECT 1.445 48.640 546.000 50.640 ;
        RECT 4.400 47.240 546.000 48.640 ;
        RECT 1.445 38.440 546.000 47.240 ;
        RECT 4.400 37.040 546.000 38.440 ;
        RECT 1.445 35.040 546.000 37.040 ;
        RECT 4.400 33.640 546.000 35.040 ;
        RECT 1.445 31.640 546.000 33.640 ;
        RECT 4.400 30.240 546.000 31.640 ;
        RECT 1.445 18.040 546.000 30.240 ;
        RECT 4.400 16.640 546.000 18.040 ;
        RECT 1.445 14.640 546.000 16.640 ;
        RECT 4.400 13.240 546.000 14.640 ;
        RECT 1.445 5.620 546.000 13.240 ;
      LAYER met4 ;
        RECT 2.135 5.615 20.640 440.465 ;
        RECT 23.040 5.615 23.940 440.465 ;
        RECT 26.340 420.080 174.240 440.465 ;
        RECT 176.640 420.080 177.540 440.465 ;
        RECT 179.940 420.080 327.840 440.465 ;
        RECT 330.240 420.700 331.140 440.465 ;
        RECT 333.540 420.700 481.440 440.465 ;
        RECT 330.240 420.080 481.440 420.700 ;
        RECT 483.840 420.080 484.740 440.465 ;
        RECT 487.140 420.080 519.160 440.465 ;
        RECT 26.340 5.615 519.160 420.080 ;
      LAYER met5 ;
        RECT 33.700 339.590 276.340 434.300 ;
        RECT 33.700 186.410 276.340 331.490 ;
        RECT 33.700 33.230 276.340 178.310 ;
        RECT 33.700 11.100 276.340 25.130 ;
  END
END BlockRAM_1KB
END LIBRARY

