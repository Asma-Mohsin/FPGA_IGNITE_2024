// This is the unpowered netlist.
module S_term_single (Co,
    UIO_BOT_UIN0,
    UIO_BOT_UIN1,
    UIO_BOT_UIN10,
    UIO_BOT_UIN11,
    UIO_BOT_UIN12,
    UIO_BOT_UIN13,
    UIO_BOT_UIN14,
    UIO_BOT_UIN15,
    UIO_BOT_UIN16,
    UIO_BOT_UIN17,
    UIO_BOT_UIN18,
    UIO_BOT_UIN19,
    UIO_BOT_UIN2,
    UIO_BOT_UIN3,
    UIO_BOT_UIN4,
    UIO_BOT_UIN5,
    UIO_BOT_UIN6,
    UIO_BOT_UIN7,
    UIO_BOT_UIN8,
    UIO_BOT_UIN9,
    UIO_BOT_UOUT0,
    UIO_BOT_UOUT1,
    UIO_BOT_UOUT10,
    UIO_BOT_UOUT11,
    UIO_BOT_UOUT12,
    UIO_BOT_UOUT13,
    UIO_BOT_UOUT14,
    UIO_BOT_UOUT15,
    UIO_BOT_UOUT16,
    UIO_BOT_UOUT17,
    UIO_BOT_UOUT18,
    UIO_BOT_UOUT19,
    UIO_BOT_UOUT2,
    UIO_BOT_UOUT3,
    UIO_BOT_UOUT4,
    UIO_BOT_UOUT5,
    UIO_BOT_UOUT6,
    UIO_BOT_UOUT7,
    UIO_BOT_UOUT8,
    UIO_BOT_UOUT9,
    UserCLK,
    UserCLKo,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N2BEG,
    N2BEGb,
    N4BEG,
    NN4BEG,
    S1END,
    S2END,
    S2MID,
    S4END,
    SS4END);
 output Co;
 input UIO_BOT_UIN0;
 input UIO_BOT_UIN1;
 input UIO_BOT_UIN10;
 input UIO_BOT_UIN11;
 input UIO_BOT_UIN12;
 input UIO_BOT_UIN13;
 input UIO_BOT_UIN14;
 input UIO_BOT_UIN15;
 input UIO_BOT_UIN16;
 input UIO_BOT_UIN17;
 input UIO_BOT_UIN18;
 input UIO_BOT_UIN19;
 input UIO_BOT_UIN2;
 input UIO_BOT_UIN3;
 input UIO_BOT_UIN4;
 input UIO_BOT_UIN5;
 input UIO_BOT_UIN6;
 input UIO_BOT_UIN7;
 input UIO_BOT_UIN8;
 input UIO_BOT_UIN9;
 output UIO_BOT_UOUT0;
 output UIO_BOT_UOUT1;
 output UIO_BOT_UOUT10;
 output UIO_BOT_UOUT11;
 output UIO_BOT_UOUT12;
 output UIO_BOT_UOUT13;
 output UIO_BOT_UOUT14;
 output UIO_BOT_UOUT15;
 output UIO_BOT_UOUT16;
 output UIO_BOT_UOUT17;
 output UIO_BOT_UOUT18;
 output UIO_BOT_UOUT19;
 output UIO_BOT_UOUT2;
 output UIO_BOT_UOUT3;
 output UIO_BOT_UOUT4;
 output UIO_BOT_UOUT5;
 output UIO_BOT_UOUT6;
 output UIO_BOT_UOUT7;
 output UIO_BOT_UOUT8;
 output UIO_BOT_UOUT9;
 input UserCLK;
 output UserCLKo;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 output [15:0] N4BEG;
 output [15:0] NN4BEG;
 input [3:0] S1END;
 input [7:0] S2END;
 input [7:0] S2MID;
 input [15:0] S4END;
 input [15:0] SS4END;

 wire net183;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_ef_sc_hd__decap_12 FILLER_0_0_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_85 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__conb_1 S_term_single_183 (.LO(net183));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__clkbuf_1 _01_ (.A(net16),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(net17),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(net18),
    .X(net107));
 sky130_fd_sc_hd__buf_1 _04_ (.A(net19),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 _05_ (.A(net20),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(net2),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_2 _07_ (.A(net3),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_2 _08_ (.A(net4),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_2 _09_ (.A(net5),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 _10_ (.A(net6),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_2 _11_ (.A(net7),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 _12_ (.A(net8),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 _13_ (.A(net9),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 _14_ (.A(net10),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_2 _15_ (.A(net11),
    .X(net100));
 sky130_fd_sc_hd__buf_1 _16_ (.A(net24),
    .X(net110));
 sky130_fd_sc_hd__buf_1 _17_ (.A(net23),
    .X(net111));
 sky130_fd_sc_hd__buf_1 _18_ (.A(net22),
    .X(net112));
 sky130_fd_sc_hd__buf_1 _19_ (.A(net21),
    .X(net113));
 sky130_fd_sc_hd__buf_1 _20_ (.A(net40),
    .X(net114));
 sky130_fd_sc_hd__buf_1 _21_ (.A(net39),
    .X(net115));
 sky130_fd_sc_hd__buf_1 _22_ (.A(net38),
    .X(net116));
 sky130_fd_sc_hd__buf_1 _23_ (.A(net37),
    .X(net117));
 sky130_fd_sc_hd__buf_1 _24_ (.A(net36),
    .X(net118));
 sky130_fd_sc_hd__buf_1 _25_ (.A(net35),
    .X(net119));
 sky130_fd_sc_hd__buf_1 _26_ (.A(net34),
    .X(net120));
 sky130_fd_sc_hd__buf_1 _27_ (.A(net33),
    .X(net121));
 sky130_fd_sc_hd__buf_1 _28_ (.A(net32),
    .X(net122));
 sky130_fd_sc_hd__buf_1 _29_ (.A(net31),
    .X(net123));
 sky130_fd_sc_hd__buf_1 _30_ (.A(net30),
    .X(net124));
 sky130_fd_sc_hd__buf_1 _31_ (.A(net29),
    .X(net125));
 sky130_fd_sc_hd__buf_1 _32_ (.A(net28),
    .X(net126));
 sky130_fd_sc_hd__buf_1 _33_ (.A(net27),
    .X(net127));
 sky130_fd_sc_hd__buf_1 _34_ (.A(net26),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _35_ (.A(net25),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _36_ (.A(net76),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _37_ (.A(net75),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _38_ (.A(net74),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _39_ (.A(net73),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _40_ (.A(net72),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _41_ (.A(net71),
    .X(net141));
 sky130_fd_sc_hd__buf_1 _42_ (.A(net88),
    .X(net142));
 sky130_fd_sc_hd__buf_1 _43_ (.A(net87),
    .X(net143));
 sky130_fd_sc_hd__buf_1 _44_ (.A(net86),
    .X(net144));
 sky130_fd_sc_hd__buf_1 _45_ (.A(net85),
    .X(net145));
 sky130_fd_sc_hd__buf_1 _46_ (.A(net84),
    .X(net131));
 sky130_fd_sc_hd__buf_1 _47_ (.A(net83),
    .X(net132));
 sky130_fd_sc_hd__buf_1 _48_ (.A(net82),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _49_ (.A(net81),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _50_ (.A(net70),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _51_ (.A(net69),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _52_ (.A(net80),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _53_ (.A(net79),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _54_ (.A(net78),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _55_ (.A(net77),
    .X(net155));
 sky130_fd_sc_hd__buf_1 _56_ (.A(net43),
    .X(net156));
 sky130_fd_sc_hd__buf_1 _57_ (.A(net42),
    .X(net157));
 sky130_fd_sc_hd__buf_1 _58_ (.A(net52),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _59_ (.A(net51),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _60_ (.A(net50),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _61_ (.A(net49),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _62_ (.A(net48),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _63_ (.A(net47),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _64_ (.A(net46),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _65_ (.A(net45),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _66_ (.A(net44),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _67_ (.A(net41),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _68_ (.A(net59),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _69_ (.A(net58),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _70_ (.A(net64),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _71_ (.A(net63),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _72_ (.A(net62),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 _73_ (.A(net61),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _74_ (.A(net60),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _75_ (.A(net53),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _76_ (.A(net46),
    .X(net170));
 sky130_fd_sc_hd__buf_1 _77_ (.A(net45),
    .X(net171));
 sky130_fd_sc_hd__buf_1 _78_ (.A(net44),
    .X(net172));
 sky130_fd_sc_hd__buf_1 _79_ (.A(net41),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _80_ (.A(net57),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _81_ (.A(net56),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _82_ (.A(net55),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _83_ (.A(net54),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 _84_ (.A(net68),
    .X(net178));
 sky130_fd_sc_hd__buf_1 _85_ (.A(net67),
    .X(net179));
 sky130_fd_sc_hd__buf_1 _86_ (.A(net66),
    .X(net180));
 sky130_fd_sc_hd__buf_1 _87_ (.A(net65),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _88_ (.A(net89),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _89_ (.A(net1),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 _90_ (.A(net12),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _91_ (.A(net13),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _92_ (.A(net14),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 _93_ (.A(net15),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(FrameStrobe[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(FrameStrobe[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(FrameStrobe[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(FrameStrobe[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(FrameStrobe[2]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(FrameStrobe[3]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(FrameStrobe[4]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(FrameStrobe[5]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(FrameStrobe[6]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(FrameStrobe[7]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(FrameStrobe[8]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(FrameStrobe[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(FrameStrobe[9]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(S1END[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(S1END[1]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(S1END[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(S1END[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(S2END[0]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(S2END[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(S2END[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(S2END[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(S2END[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(FrameStrobe[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(S2END[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(S2END[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(S2END[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(S2MID[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(S2MID[1]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(S2MID[2]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(S2MID[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(S2MID[4]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(S2MID[5]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(S2MID[6]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(FrameStrobe[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(S2MID[7]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(S4END[0]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(S4END[10]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(S4END[11]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(S4END[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(S4END[2]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(S4END[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(S4END[4]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(S4END[5]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(S4END[6]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(FrameStrobe[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(S4END[7]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(S4END[8]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(S4END[9]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(SS4END[0]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(SS4END[10]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(SS4END[11]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(SS4END[12]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(SS4END[13]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(SS4END[14]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(SS4END[15]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(FrameStrobe[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(SS4END[1]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(SS4END[2]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(SS4END[3]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(SS4END[4]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(SS4END[5]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(SS4END[6]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(SS4END[7]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(SS4END[8]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(SS4END[9]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(UIO_BOT_UIN0),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(FrameStrobe[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(UIO_BOT_UIN1),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(UIO_BOT_UIN10),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(UIO_BOT_UIN11),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(UIO_BOT_UIN12),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(UIO_BOT_UIN13),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(UIO_BOT_UIN14),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(UIO_BOT_UIN15),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(UIO_BOT_UIN16),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(UIO_BOT_UIN17),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(UIO_BOT_UIN18),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(FrameStrobe[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(UIO_BOT_UIN19),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(UIO_BOT_UIN2),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(UIO_BOT_UIN3),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(UIO_BOT_UIN4),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(UIO_BOT_UIN5),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(UIO_BOT_UIN6),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(UIO_BOT_UIN7),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(UIO_BOT_UIN8),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(UIO_BOT_UIN9),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(UserCLK),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(FrameStrobe[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output100 (.A(net100),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output101 (.A(net101),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__clkbuf_4 output102 (.A(net102),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output103 (.A(net103),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output104 (.A(net104),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output105 (.A(net105),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output106 (.A(net106),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output107 (.A(net107),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output108 (.A(net108),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output109 (.A(net109),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output110 (.A(net110),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output111 (.A(net111),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output112 (.A(net112),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output113 (.A(net113),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output114 (.A(net114),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output115 (.A(net115),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output116 (.A(net116),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output117 (.A(net117),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output118 (.A(net118),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output119 (.A(net119),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output120 (.A(net120),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output121 (.A(net121),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output122 (.A(net122),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output123 (.A(net123),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output124 (.A(net124),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output125 (.A(net125),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output126 (.A(net126),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output127 (.A(net127),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output128 (.A(net128),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output129 (.A(net129),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output130 (.A(net130),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output131 (.A(net131),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output132 (.A(net132),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output133 (.A(net133),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output134 (.A(net134),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output135 (.A(net135),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output136 (.A(net136),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output137 (.A(net137),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output138 (.A(net138),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output139 (.A(net139),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output140 (.A(net140),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output141 (.A(net141),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output142 (.A(net142),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output143 (.A(net143),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output144 (.A(net144),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output145 (.A(net145),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output146 (.A(net146),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output147 (.A(net147),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output148 (.A(net148),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output149 (.A(net149),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output150 (.A(net150),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output151 (.A(net151),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output152 (.A(net152),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output153 (.A(net153),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output154 (.A(net154),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output155 (.A(net155),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output156 (.A(net156),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output157 (.A(net157),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output158 (.A(net158),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output159 (.A(net159),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output160 (.A(net160),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output161 (.A(net161),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output162 (.A(net162),
    .X(UIO_BOT_UOUT0));
 sky130_fd_sc_hd__clkbuf_4 output163 (.A(net163),
    .X(UIO_BOT_UOUT1));
 sky130_fd_sc_hd__clkbuf_4 output164 (.A(net164),
    .X(UIO_BOT_UOUT10));
 sky130_fd_sc_hd__clkbuf_4 output165 (.A(net165),
    .X(UIO_BOT_UOUT11));
 sky130_fd_sc_hd__clkbuf_4 output166 (.A(net166),
    .X(UIO_BOT_UOUT12));
 sky130_fd_sc_hd__clkbuf_4 output167 (.A(net167),
    .X(UIO_BOT_UOUT13));
 sky130_fd_sc_hd__clkbuf_4 output168 (.A(net168),
    .X(UIO_BOT_UOUT14));
 sky130_fd_sc_hd__clkbuf_4 output169 (.A(net169),
    .X(UIO_BOT_UOUT15));
 sky130_fd_sc_hd__clkbuf_4 output170 (.A(net170),
    .X(UIO_BOT_UOUT16));
 sky130_fd_sc_hd__clkbuf_4 output171 (.A(net171),
    .X(UIO_BOT_UOUT17));
 sky130_fd_sc_hd__clkbuf_4 output172 (.A(net172),
    .X(UIO_BOT_UOUT18));
 sky130_fd_sc_hd__clkbuf_4 output173 (.A(net173),
    .X(UIO_BOT_UOUT19));
 sky130_fd_sc_hd__clkbuf_4 output174 (.A(net174),
    .X(UIO_BOT_UOUT2));
 sky130_fd_sc_hd__clkbuf_4 output175 (.A(net175),
    .X(UIO_BOT_UOUT3));
 sky130_fd_sc_hd__clkbuf_4 output176 (.A(net176),
    .X(UIO_BOT_UOUT4));
 sky130_fd_sc_hd__clkbuf_4 output177 (.A(net177),
    .X(UIO_BOT_UOUT5));
 sky130_fd_sc_hd__clkbuf_4 output178 (.A(net178),
    .X(UIO_BOT_UOUT6));
 sky130_fd_sc_hd__clkbuf_4 output179 (.A(net179),
    .X(UIO_BOT_UOUT7));
 sky130_fd_sc_hd__clkbuf_4 output180 (.A(net180),
    .X(UIO_BOT_UOUT8));
 sky130_fd_sc_hd__clkbuf_4 output181 (.A(net181),
    .X(UIO_BOT_UOUT9));
 sky130_fd_sc_hd__clkbuf_4 output182 (.A(net182),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output90 (.A(net90),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output91 (.A(net91),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output92 (.A(net92),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output93 (.A(net93),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output94 (.A(net94),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output95 (.A(net95),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output96 (.A(net96),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output97 (.A(net97),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output98 (.A(net98),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output99 (.A(net99),
    .X(FrameStrobe_O[18]));
 assign Co = net183;
endmodule

