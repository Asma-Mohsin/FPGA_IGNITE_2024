magic
tech sky130A
magscale 1 2
timestamp 1732489753
<< obsli1 >>
rect 1104 1071 24840 6545
<< obsm1 >>
rect 290 892 25654 7948
<< metal2 >>
rect 202 7840 258 8000
rect 478 7840 534 8000
rect 754 7840 810 8000
rect 1030 7840 1086 8000
rect 1306 7840 1362 8000
rect 1582 7840 1638 8000
rect 1858 7840 1914 8000
rect 2134 7840 2190 8000
rect 2410 7840 2466 8000
rect 2686 7840 2742 8000
rect 2962 7840 3018 8000
rect 3238 7840 3294 8000
rect 3514 7840 3570 8000
rect 3790 7840 3846 8000
rect 4066 7840 4122 8000
rect 4342 7840 4398 8000
rect 4618 7840 4674 8000
rect 4894 7840 4950 8000
rect 5170 7840 5226 8000
rect 5446 7840 5502 8000
rect 5722 7840 5778 8000
rect 5998 7840 6054 8000
rect 6274 7840 6330 8000
rect 6550 7840 6606 8000
rect 6826 7840 6882 8000
rect 7102 7840 7158 8000
rect 7378 7840 7434 8000
rect 7654 7840 7710 8000
rect 7930 7840 7986 8000
rect 8206 7840 8262 8000
rect 8482 7840 8538 8000
rect 8758 7840 8814 8000
rect 9034 7840 9090 8000
rect 9310 7840 9366 8000
rect 9586 7840 9642 8000
rect 9862 7840 9918 8000
rect 10138 7840 10194 8000
rect 10414 7840 10470 8000
rect 10690 7840 10746 8000
rect 10966 7840 11022 8000
rect 11242 7840 11298 8000
rect 11518 7840 11574 8000
rect 11794 7840 11850 8000
rect 12070 7840 12126 8000
rect 12346 7840 12402 8000
rect 12622 7840 12678 8000
rect 12898 7840 12954 8000
rect 13174 7840 13230 8000
rect 13450 7840 13506 8000
rect 13726 7840 13782 8000
rect 14002 7840 14058 8000
rect 14278 7840 14334 8000
rect 14554 7840 14610 8000
rect 14830 7840 14886 8000
rect 15106 7840 15162 8000
rect 15382 7840 15438 8000
rect 15658 7840 15714 8000
rect 15934 7840 15990 8000
rect 16210 7840 16266 8000
rect 16486 7840 16542 8000
rect 16762 7840 16818 8000
rect 17038 7840 17094 8000
rect 17314 7840 17370 8000
rect 17590 7840 17646 8000
rect 17866 7840 17922 8000
rect 18142 7840 18198 8000
rect 18418 7840 18474 8000
rect 18694 7840 18750 8000
rect 18970 7840 19026 8000
rect 19246 7840 19302 8000
rect 19522 7840 19578 8000
rect 19798 7840 19854 8000
rect 20074 7840 20130 8000
rect 20350 7840 20406 8000
rect 20626 7840 20682 8000
rect 20902 7840 20958 8000
rect 21178 7840 21234 8000
rect 21454 7840 21510 8000
rect 21730 7840 21786 8000
rect 22006 7840 22062 8000
rect 22282 7840 22338 8000
rect 22558 7840 22614 8000
rect 22834 7840 22890 8000
rect 23110 7840 23166 8000
rect 23386 7840 23442 8000
rect 23662 7840 23718 8000
rect 23938 7840 23994 8000
rect 24214 7840 24270 8000
rect 24490 7840 24546 8000
rect 24766 7840 24822 8000
rect 25042 7840 25098 8000
rect 25318 7840 25374 8000
rect 25594 7840 25650 8000
rect 938 0 994 160
rect 2134 0 2190 160
rect 3330 0 3386 160
rect 4526 0 4582 160
rect 5722 0 5778 160
rect 6918 0 6974 160
rect 8114 0 8170 160
rect 9310 0 9366 160
rect 10506 0 10562 160
rect 11702 0 11758 160
rect 12898 0 12954 160
rect 14094 0 14150 160
rect 15290 0 15346 160
rect 16486 0 16542 160
rect 17682 0 17738 160
rect 18878 0 18934 160
rect 20074 0 20130 160
rect 21270 0 21326 160
rect 22466 0 22522 160
rect 23662 0 23718 160
rect 24858 0 24914 160
<< obsm2 >>
rect 314 7784 422 7970
rect 590 7784 698 7970
rect 866 7784 974 7970
rect 1142 7784 1250 7970
rect 1418 7784 1526 7970
rect 1694 7784 1802 7970
rect 1970 7784 2078 7970
rect 2246 7784 2354 7970
rect 2522 7784 2630 7970
rect 2798 7784 2906 7970
rect 3074 7784 3182 7970
rect 3350 7784 3458 7970
rect 3626 7784 3734 7970
rect 3902 7784 4010 7970
rect 4178 7784 4286 7970
rect 4454 7784 4562 7970
rect 4730 7784 4838 7970
rect 5006 7784 5114 7970
rect 5282 7784 5390 7970
rect 5558 7784 5666 7970
rect 5834 7784 5942 7970
rect 6110 7784 6218 7970
rect 6386 7784 6494 7970
rect 6662 7784 6770 7970
rect 6938 7784 7046 7970
rect 7214 7784 7322 7970
rect 7490 7784 7598 7970
rect 7766 7784 7874 7970
rect 8042 7784 8150 7970
rect 8318 7784 8426 7970
rect 8594 7784 8702 7970
rect 8870 7784 8978 7970
rect 9146 7784 9254 7970
rect 9422 7784 9530 7970
rect 9698 7784 9806 7970
rect 9974 7784 10082 7970
rect 10250 7784 10358 7970
rect 10526 7784 10634 7970
rect 10802 7784 10910 7970
rect 11078 7784 11186 7970
rect 11354 7784 11462 7970
rect 11630 7784 11738 7970
rect 11906 7784 12014 7970
rect 12182 7784 12290 7970
rect 12458 7784 12566 7970
rect 12734 7784 12842 7970
rect 13010 7784 13118 7970
rect 13286 7784 13394 7970
rect 13562 7784 13670 7970
rect 13838 7784 13946 7970
rect 14114 7784 14222 7970
rect 14390 7784 14498 7970
rect 14666 7784 14774 7970
rect 14942 7784 15050 7970
rect 15218 7784 15326 7970
rect 15494 7784 15602 7970
rect 15770 7784 15878 7970
rect 16046 7784 16154 7970
rect 16322 7784 16430 7970
rect 16598 7784 16706 7970
rect 16874 7784 16982 7970
rect 17150 7784 17258 7970
rect 17426 7784 17534 7970
rect 17702 7784 17810 7970
rect 17978 7784 18086 7970
rect 18254 7784 18362 7970
rect 18530 7784 18638 7970
rect 18806 7784 18914 7970
rect 19082 7784 19190 7970
rect 19358 7784 19466 7970
rect 19634 7784 19742 7970
rect 19910 7784 20018 7970
rect 20186 7784 20294 7970
rect 20462 7784 20570 7970
rect 20738 7784 20846 7970
rect 21014 7784 21122 7970
rect 21290 7784 21398 7970
rect 21566 7784 21674 7970
rect 21842 7784 21950 7970
rect 22118 7784 22226 7970
rect 22394 7784 22502 7970
rect 22670 7784 22778 7970
rect 22946 7784 23054 7970
rect 23222 7784 23330 7970
rect 23498 7784 23606 7970
rect 23774 7784 23882 7970
rect 24050 7784 24158 7970
rect 24326 7784 24434 7970
rect 24602 7784 24710 7970
rect 24878 7784 24986 7970
rect 25154 7784 25262 7970
rect 25430 7784 25538 7970
rect 216 216 25648 7784
rect 216 54 882 216
rect 1050 54 2078 216
rect 2246 54 3274 216
rect 3442 54 4470 216
rect 4638 54 5666 216
rect 5834 54 6862 216
rect 7030 54 8058 216
rect 8226 54 9254 216
rect 9422 54 10450 216
rect 10618 54 11646 216
rect 11814 54 12842 216
rect 13010 54 14038 216
rect 14206 54 15234 216
rect 15402 54 16430 216
rect 16598 54 17626 216
rect 17794 54 18822 216
rect 18990 54 20018 216
rect 20186 54 21214 216
rect 21382 54 22410 216
rect 22578 54 23606 216
rect 23774 54 24802 216
rect 24970 54 25648 216
<< obsm3 >>
rect 1761 1055 24998 6561
<< metal4 >>
rect 3911 1040 4231 6576
rect 6878 1040 7198 6576
rect 9845 1040 10165 6576
rect 12812 1040 13132 6576
rect 15779 1040 16099 6576
rect 18746 1040 19066 6576
rect 21713 1040 22033 6576
rect 24680 1040 25000 6576
<< obsm4 >>
rect 17907 1395 18666 6221
rect 19146 1395 21633 6221
rect 22113 1395 22757 6221
<< labels >>
rlabel metal2 s 2134 0 2190 160 6 FrameStrobe[0]
port 1 nsew signal input
rlabel metal2 s 14094 0 14150 160 6 FrameStrobe[10]
port 2 nsew signal input
rlabel metal2 s 15290 0 15346 160 6 FrameStrobe[11]
port 3 nsew signal input
rlabel metal2 s 16486 0 16542 160 6 FrameStrobe[12]
port 4 nsew signal input
rlabel metal2 s 17682 0 17738 160 6 FrameStrobe[13]
port 5 nsew signal input
rlabel metal2 s 18878 0 18934 160 6 FrameStrobe[14]
port 6 nsew signal input
rlabel metal2 s 20074 0 20130 160 6 FrameStrobe[15]
port 7 nsew signal input
rlabel metal2 s 21270 0 21326 160 6 FrameStrobe[16]
port 8 nsew signal input
rlabel metal2 s 22466 0 22522 160 6 FrameStrobe[17]
port 9 nsew signal input
rlabel metal2 s 23662 0 23718 160 6 FrameStrobe[18]
port 10 nsew signal input
rlabel metal2 s 24858 0 24914 160 6 FrameStrobe[19]
port 11 nsew signal input
rlabel metal2 s 3330 0 3386 160 6 FrameStrobe[1]
port 12 nsew signal input
rlabel metal2 s 4526 0 4582 160 6 FrameStrobe[2]
port 13 nsew signal input
rlabel metal2 s 5722 0 5778 160 6 FrameStrobe[3]
port 14 nsew signal input
rlabel metal2 s 6918 0 6974 160 6 FrameStrobe[4]
port 15 nsew signal input
rlabel metal2 s 8114 0 8170 160 6 FrameStrobe[5]
port 16 nsew signal input
rlabel metal2 s 9310 0 9366 160 6 FrameStrobe[6]
port 17 nsew signal input
rlabel metal2 s 10506 0 10562 160 6 FrameStrobe[7]
port 18 nsew signal input
rlabel metal2 s 11702 0 11758 160 6 FrameStrobe[8]
port 19 nsew signal input
rlabel metal2 s 12898 0 12954 160 6 FrameStrobe[9]
port 20 nsew signal input
rlabel metal2 s 20350 7840 20406 8000 6 FrameStrobe_O[0]
port 21 nsew signal output
rlabel metal2 s 23110 7840 23166 8000 6 FrameStrobe_O[10]
port 22 nsew signal output
rlabel metal2 s 23386 7840 23442 8000 6 FrameStrobe_O[11]
port 23 nsew signal output
rlabel metal2 s 23662 7840 23718 8000 6 FrameStrobe_O[12]
port 24 nsew signal output
rlabel metal2 s 23938 7840 23994 8000 6 FrameStrobe_O[13]
port 25 nsew signal output
rlabel metal2 s 24214 7840 24270 8000 6 FrameStrobe_O[14]
port 26 nsew signal output
rlabel metal2 s 24490 7840 24546 8000 6 FrameStrobe_O[15]
port 27 nsew signal output
rlabel metal2 s 24766 7840 24822 8000 6 FrameStrobe_O[16]
port 28 nsew signal output
rlabel metal2 s 25042 7840 25098 8000 6 FrameStrobe_O[17]
port 29 nsew signal output
rlabel metal2 s 25318 7840 25374 8000 6 FrameStrobe_O[18]
port 30 nsew signal output
rlabel metal2 s 25594 7840 25650 8000 6 FrameStrobe_O[19]
port 31 nsew signal output
rlabel metal2 s 20626 7840 20682 8000 6 FrameStrobe_O[1]
port 32 nsew signal output
rlabel metal2 s 20902 7840 20958 8000 6 FrameStrobe_O[2]
port 33 nsew signal output
rlabel metal2 s 21178 7840 21234 8000 6 FrameStrobe_O[3]
port 34 nsew signal output
rlabel metal2 s 21454 7840 21510 8000 6 FrameStrobe_O[4]
port 35 nsew signal output
rlabel metal2 s 21730 7840 21786 8000 6 FrameStrobe_O[5]
port 36 nsew signal output
rlabel metal2 s 22006 7840 22062 8000 6 FrameStrobe_O[6]
port 37 nsew signal output
rlabel metal2 s 22282 7840 22338 8000 6 FrameStrobe_O[7]
port 38 nsew signal output
rlabel metal2 s 22558 7840 22614 8000 6 FrameStrobe_O[8]
port 39 nsew signal output
rlabel metal2 s 22834 7840 22890 8000 6 FrameStrobe_O[9]
port 40 nsew signal output
rlabel metal2 s 202 7840 258 8000 6 N1BEG[0]
port 41 nsew signal output
rlabel metal2 s 478 7840 534 8000 6 N1BEG[1]
port 42 nsew signal output
rlabel metal2 s 754 7840 810 8000 6 N1BEG[2]
port 43 nsew signal output
rlabel metal2 s 1030 7840 1086 8000 6 N1BEG[3]
port 44 nsew signal output
rlabel metal2 s 1306 7840 1362 8000 6 N2BEG[0]
port 45 nsew signal output
rlabel metal2 s 1582 7840 1638 8000 6 N2BEG[1]
port 46 nsew signal output
rlabel metal2 s 1858 7840 1914 8000 6 N2BEG[2]
port 47 nsew signal output
rlabel metal2 s 2134 7840 2190 8000 6 N2BEG[3]
port 48 nsew signal output
rlabel metal2 s 2410 7840 2466 8000 6 N2BEG[4]
port 49 nsew signal output
rlabel metal2 s 2686 7840 2742 8000 6 N2BEG[5]
port 50 nsew signal output
rlabel metal2 s 2962 7840 3018 8000 6 N2BEG[6]
port 51 nsew signal output
rlabel metal2 s 3238 7840 3294 8000 6 N2BEG[7]
port 52 nsew signal output
rlabel metal2 s 3514 7840 3570 8000 6 N2BEGb[0]
port 53 nsew signal output
rlabel metal2 s 3790 7840 3846 8000 6 N2BEGb[1]
port 54 nsew signal output
rlabel metal2 s 4066 7840 4122 8000 6 N2BEGb[2]
port 55 nsew signal output
rlabel metal2 s 4342 7840 4398 8000 6 N2BEGb[3]
port 56 nsew signal output
rlabel metal2 s 4618 7840 4674 8000 6 N2BEGb[4]
port 57 nsew signal output
rlabel metal2 s 4894 7840 4950 8000 6 N2BEGb[5]
port 58 nsew signal output
rlabel metal2 s 5170 7840 5226 8000 6 N2BEGb[6]
port 59 nsew signal output
rlabel metal2 s 5446 7840 5502 8000 6 N2BEGb[7]
port 60 nsew signal output
rlabel metal2 s 5722 7840 5778 8000 6 N4BEG[0]
port 61 nsew signal output
rlabel metal2 s 8482 7840 8538 8000 6 N4BEG[10]
port 62 nsew signal output
rlabel metal2 s 8758 7840 8814 8000 6 N4BEG[11]
port 63 nsew signal output
rlabel metal2 s 9034 7840 9090 8000 6 N4BEG[12]
port 64 nsew signal output
rlabel metal2 s 9310 7840 9366 8000 6 N4BEG[13]
port 65 nsew signal output
rlabel metal2 s 9586 7840 9642 8000 6 N4BEG[14]
port 66 nsew signal output
rlabel metal2 s 9862 7840 9918 8000 6 N4BEG[15]
port 67 nsew signal output
rlabel metal2 s 5998 7840 6054 8000 6 N4BEG[1]
port 68 nsew signal output
rlabel metal2 s 6274 7840 6330 8000 6 N4BEG[2]
port 69 nsew signal output
rlabel metal2 s 6550 7840 6606 8000 6 N4BEG[3]
port 70 nsew signal output
rlabel metal2 s 6826 7840 6882 8000 6 N4BEG[4]
port 71 nsew signal output
rlabel metal2 s 7102 7840 7158 8000 6 N4BEG[5]
port 72 nsew signal output
rlabel metal2 s 7378 7840 7434 8000 6 N4BEG[6]
port 73 nsew signal output
rlabel metal2 s 7654 7840 7710 8000 6 N4BEG[7]
port 74 nsew signal output
rlabel metal2 s 7930 7840 7986 8000 6 N4BEG[8]
port 75 nsew signal output
rlabel metal2 s 8206 7840 8262 8000 6 N4BEG[9]
port 76 nsew signal output
rlabel metal2 s 10138 7840 10194 8000 6 S1END[0]
port 77 nsew signal input
rlabel metal2 s 10414 7840 10470 8000 6 S1END[1]
port 78 nsew signal input
rlabel metal2 s 10690 7840 10746 8000 6 S1END[2]
port 79 nsew signal input
rlabel metal2 s 10966 7840 11022 8000 6 S1END[3]
port 80 nsew signal input
rlabel metal2 s 11242 7840 11298 8000 6 S2END[0]
port 81 nsew signal input
rlabel metal2 s 11518 7840 11574 8000 6 S2END[1]
port 82 nsew signal input
rlabel metal2 s 11794 7840 11850 8000 6 S2END[2]
port 83 nsew signal input
rlabel metal2 s 12070 7840 12126 8000 6 S2END[3]
port 84 nsew signal input
rlabel metal2 s 12346 7840 12402 8000 6 S2END[4]
port 85 nsew signal input
rlabel metal2 s 12622 7840 12678 8000 6 S2END[5]
port 86 nsew signal input
rlabel metal2 s 12898 7840 12954 8000 6 S2END[6]
port 87 nsew signal input
rlabel metal2 s 13174 7840 13230 8000 6 S2END[7]
port 88 nsew signal input
rlabel metal2 s 13450 7840 13506 8000 6 S2MID[0]
port 89 nsew signal input
rlabel metal2 s 13726 7840 13782 8000 6 S2MID[1]
port 90 nsew signal input
rlabel metal2 s 14002 7840 14058 8000 6 S2MID[2]
port 91 nsew signal input
rlabel metal2 s 14278 7840 14334 8000 6 S2MID[3]
port 92 nsew signal input
rlabel metal2 s 14554 7840 14610 8000 6 S2MID[4]
port 93 nsew signal input
rlabel metal2 s 14830 7840 14886 8000 6 S2MID[5]
port 94 nsew signal input
rlabel metal2 s 15106 7840 15162 8000 6 S2MID[6]
port 95 nsew signal input
rlabel metal2 s 15382 7840 15438 8000 6 S2MID[7]
port 96 nsew signal input
rlabel metal2 s 15658 7840 15714 8000 6 S4END[0]
port 97 nsew signal input
rlabel metal2 s 18418 7840 18474 8000 6 S4END[10]
port 98 nsew signal input
rlabel metal2 s 18694 7840 18750 8000 6 S4END[11]
port 99 nsew signal input
rlabel metal2 s 18970 7840 19026 8000 6 S4END[12]
port 100 nsew signal input
rlabel metal2 s 19246 7840 19302 8000 6 S4END[13]
port 101 nsew signal input
rlabel metal2 s 19522 7840 19578 8000 6 S4END[14]
port 102 nsew signal input
rlabel metal2 s 19798 7840 19854 8000 6 S4END[15]
port 103 nsew signal input
rlabel metal2 s 15934 7840 15990 8000 6 S4END[1]
port 104 nsew signal input
rlabel metal2 s 16210 7840 16266 8000 6 S4END[2]
port 105 nsew signal input
rlabel metal2 s 16486 7840 16542 8000 6 S4END[3]
port 106 nsew signal input
rlabel metal2 s 16762 7840 16818 8000 6 S4END[4]
port 107 nsew signal input
rlabel metal2 s 17038 7840 17094 8000 6 S4END[5]
port 108 nsew signal input
rlabel metal2 s 17314 7840 17370 8000 6 S4END[6]
port 109 nsew signal input
rlabel metal2 s 17590 7840 17646 8000 6 S4END[7]
port 110 nsew signal input
rlabel metal2 s 17866 7840 17922 8000 6 S4END[8]
port 111 nsew signal input
rlabel metal2 s 18142 7840 18198 8000 6 S4END[9]
port 112 nsew signal input
rlabel metal2 s 938 0 994 160 6 UserCLK
port 113 nsew signal input
rlabel metal2 s 20074 7840 20130 8000 6 UserCLKo
port 114 nsew signal output
rlabel metal4 s 6878 1040 7198 6576 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 12812 1040 13132 6576 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 18746 1040 19066 6576 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 24680 1040 25000 6576 6 VGND
port 115 nsew ground bidirectional
rlabel metal4 s 3911 1040 4231 6576 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 9845 1040 10165 6576 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 15779 1040 16099 6576 6 VPWR
port 116 nsew power bidirectional
rlabel metal4 s 21713 1040 22033 6576 6 VPWR
port 116 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 26000 8000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 464816
string GDS_FILE /home/asma/Desktop/FPGA_IGNITE_2024/openlane/S_term_RAMIO_redo/runs/24_11_24_23_07/results/signoff/S_term_RAM_IO.magic.gds
string GDS_START 37874
<< end >>

