VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_single
  CLASS BLOCK ;
  FOREIGN S_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 182.000 ;
  PIN Co
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.000 181.300 104.380 182.000 ;
    END
  END Co
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 46.040 0.000 46.420 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 50.180 0.000 50.560 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 53.860 0.000 54.240 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 0.000 58.380 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 62.140 0.000 62.520 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 66.280 0.000 66.660 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 69.960 0.000 70.340 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.100 0.000 74.480 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 78.240 0.000 78.620 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.380 0.000 82.760 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 9.700 0.000 10.080 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 13.840 0.000 14.220 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 17.520 0.000 17.900 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 21.660 0.000 22.040 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 25.800 0.000 26.180 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.940 0.000 30.320 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 33.620 0.000 34.000 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.760 0.000 38.140 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.900 0.000 42.280 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 206.120 181.300 206.500 182.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 225.440 181.300 225.820 182.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 227.280 181.300 227.660 182.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 229.120 181.300 229.500 182.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 230.960 181.300 231.340 182.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 233.260 181.300 233.640 182.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 235.100 181.300 235.480 182.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 236.940 181.300 237.320 182.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 238.780 181.300 239.160 182.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 240.620 181.300 241.000 182.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 242.920 181.300 243.300 182.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 207.960 181.300 208.340 182.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 209.800 181.300 210.180 182.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 211.640 181.300 212.020 182.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 213.940 181.300 214.320 182.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 215.780 181.300 216.160 182.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 217.620 181.300 218.000 182.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.460 181.300 219.840 182.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 221.300 181.300 221.680 182.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 223.600 181.300 223.980 182.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 3.720 181.300 4.100 182.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 5.560 181.300 5.940 182.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 7.400 181.300 7.780 182.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 9.240 181.300 9.620 182.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 11.080 181.300 11.460 182.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 13.380 181.300 13.760 182.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 15.220 181.300 15.600 182.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.060 181.300 17.440 182.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 18.900 181.300 19.280 182.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 20.740 181.300 21.120 182.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 22.580 181.300 22.960 182.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.880 181.300 25.260 182.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 26.720 181.300 27.100 182.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 28.560 181.300 28.940 182.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 30.400 181.300 30.780 182.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.240 181.300 32.620 182.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 34.540 181.300 34.920 182.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.380 181.300 36.760 182.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.220 181.300 38.600 182.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 40.060 181.300 40.440 182.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 41.900 181.300 42.280 182.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 61.220 181.300 61.600 182.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.520 181.300 63.900 182.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.360 181.300 65.740 182.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.200 181.300 67.580 182.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.040 181.300 69.420 182.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.880 181.300 71.260 182.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.200 181.300 44.580 182.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.040 181.300 46.420 182.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.880 181.300 48.260 182.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 49.720 181.300 50.100 182.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.560 181.300 51.940 182.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 53.860 181.300 54.240 182.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 55.700 181.300 56.080 182.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 57.540 181.300 57.920 182.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.380 181.300 59.760 182.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 73.180 181.300 73.560 182.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 92.040 181.300 92.420 182.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.340 181.300 94.720 182.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.180 181.300 96.560 182.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.020 181.300 98.400 182.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.860 181.300 100.240 182.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 101.700 181.300 102.080 182.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.020 181.300 75.400 182.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 76.860 181.300 77.240 182.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.700 181.300 79.080 182.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.540 181.300 80.920 182.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.380 181.300 82.760 182.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.680 181.300 85.060 182.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 181.300 86.900 182.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.360 181.300 88.740 182.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.200 181.300 90.580 182.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 105.840 181.300 106.220 182.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 107.680 181.300 108.060 182.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 109.520 181.300 109.900 182.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 111.360 181.300 111.740 182.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 128.840 181.300 129.220 182.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 130.680 181.300 131.060 182.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 132.980 181.300 133.360 182.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 134.820 181.300 135.200 182.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.660 181.300 137.040 182.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 138.500 181.300 138.880 182.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 140.340 181.300 140.720 182.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 142.180 181.300 142.560 182.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 113.660 181.300 114.040 182.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 115.500 181.300 115.880 182.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 117.340 181.300 117.720 182.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 119.180 181.300 119.560 182.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 121.020 181.300 121.400 182.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 123.320 181.300 123.700 182.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 125.160 181.300 125.540 182.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 127.000 181.300 127.380 182.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.480 181.300 144.860 182.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.800 181.300 164.180 182.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.640 181.300 166.020 182.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.480 181.300 167.860 182.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.320 181.300 169.700 182.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.160 181.300 171.540 182.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.460 181.300 173.840 182.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 181.300 146.700 182.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 148.160 181.300 148.540 182.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 150.000 181.300 150.380 182.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 151.840 181.300 152.220 182.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 154.140 181.300 154.520 182.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 155.980 181.300 156.360 182.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 157.820 181.300 158.200 182.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 159.660 181.300 160.040 182.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 161.500 181.300 161.880 182.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 175.300 181.300 175.680 182.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 194.620 181.300 195.000 182.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 196.460 181.300 196.840 182.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 198.300 181.300 198.680 182.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 200.140 181.300 200.520 182.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 201.980 181.300 202.360 182.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 204.280 181.300 204.660 182.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 177.140 181.300 177.520 182.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 178.980 181.300 179.360 182.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.820 181.300 181.200 182.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 183.120 181.300 183.500 182.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 184.960 181.300 185.340 182.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 186.800 181.300 187.180 182.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 188.640 181.300 189.020 182.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.480 181.300 190.860 182.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 192.780 181.300 193.160 182.000 ;
    END
  END SS4END[9]
  PIN UIO_BOT_UIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.020 0.000 167.400 0.700 ;
    END
  END UIO_BOT_UIN0
  PIN UIO_BOT_UIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 171.160 0.000 171.540 0.700 ;
    END
  END UIO_BOT_UIN1
  PIN UIO_BOT_UIN10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 174.840 0.000 175.220 0.700 ;
    END
  END UIO_BOT_UIN10
  PIN UIO_BOT_UIN11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 178.980 0.000 179.360 0.700 ;
    END
  END UIO_BOT_UIN11
  PIN UIO_BOT_UIN12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.120 0.000 183.500 0.700 ;
    END
  END UIO_BOT_UIN12
  PIN UIO_BOT_UIN13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 187.260 0.000 187.640 0.700 ;
    END
  END UIO_BOT_UIN13
  PIN UIO_BOT_UIN14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 190.940 0.000 191.320 0.700 ;
    END
  END UIO_BOT_UIN14
  PIN UIO_BOT_UIN15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 195.080 0.000 195.460 0.700 ;
    END
  END UIO_BOT_UIN15
  PIN UIO_BOT_UIN16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 199.220 0.000 199.600 0.700 ;
    END
  END UIO_BOT_UIN16
  PIN UIO_BOT_UIN17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 203.360 0.000 203.740 0.700 ;
    END
  END UIO_BOT_UIN17
  PIN UIO_BOT_UIN18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 207.040 0.000 207.420 0.700 ;
    END
  END UIO_BOT_UIN18
  PIN UIO_BOT_UIN19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 211.180 0.000 211.560 0.700 ;
    END
  END UIO_BOT_UIN19
  PIN UIO_BOT_UIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 215.320 0.000 215.700 0.700 ;
    END
  END UIO_BOT_UIN2
  PIN UIO_BOT_UIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 219.460 0.000 219.840 0.700 ;
    END
  END UIO_BOT_UIN3
  PIN UIO_BOT_UIN4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 223.600 0.000 223.980 0.700 ;
    END
  END UIO_BOT_UIN4
  PIN UIO_BOT_UIN5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 227.280 0.000 227.660 0.700 ;
    END
  END UIO_BOT_UIN5
  PIN UIO_BOT_UIN6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 231.420 0.000 231.800 0.700 ;
    END
  END UIO_BOT_UIN6
  PIN UIO_BOT_UIN7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 235.560 0.000 235.940 0.700 ;
    END
  END UIO_BOT_UIN7
  PIN UIO_BOT_UIN8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 239.700 0.000 240.080 0.700 ;
    END
  END UIO_BOT_UIN8
  PIN UIO_BOT_UIN9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 243.380 0.000 243.760 0.700 ;
    END
  END UIO_BOT_UIN9
  PIN UIO_BOT_UOUT0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.060 0.000 86.440 0.700 ;
    END
  END UIO_BOT_UOUT0
  PIN UIO_BOT_UOUT1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 90.200 0.000 90.580 0.700 ;
    END
  END UIO_BOT_UOUT1
  PIN UIO_BOT_UOUT10
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.340 0.000 94.720 0.700 ;
    END
  END UIO_BOT_UOUT10
  PIN UIO_BOT_UOUT11
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 0.000 98.860 0.700 ;
    END
  END UIO_BOT_UOUT11
  PIN UIO_BOT_UOUT12
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 102.620 0.000 103.000 0.700 ;
    END
  END UIO_BOT_UOUT12
  PIN UIO_BOT_UOUT13
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.300 0.000 106.680 0.700 ;
    END
  END UIO_BOT_UOUT13
  PIN UIO_BOT_UOUT14
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 110.440 0.000 110.820 0.700 ;
    END
  END UIO_BOT_UOUT14
  PIN UIO_BOT_UOUT15
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.580 0.000 114.960 0.700 ;
    END
  END UIO_BOT_UOUT15
  PIN UIO_BOT_UOUT16
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 118.720 0.000 119.100 0.700 ;
    END
  END UIO_BOT_UOUT16
  PIN UIO_BOT_UOUT17
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 122.400 0.000 122.780 0.700 ;
    END
  END UIO_BOT_UOUT17
  PIN UIO_BOT_UOUT18
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 126.540 0.000 126.920 0.700 ;
    END
  END UIO_BOT_UOUT18
  PIN UIO_BOT_UOUT19
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.680 0.000 131.060 0.700 ;
    END
  END UIO_BOT_UOUT19
  PIN UIO_BOT_UOUT2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 134.820 0.000 135.200 0.700 ;
    END
  END UIO_BOT_UOUT2
  PIN UIO_BOT_UOUT3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.500 0.000 138.880 0.700 ;
    END
  END UIO_BOT_UOUT3
  PIN UIO_BOT_UOUT4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 142.640 0.000 143.020 0.700 ;
    END
  END UIO_BOT_UOUT4
  PIN UIO_BOT_UOUT5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 0.000 147.160 0.700 ;
    END
  END UIO_BOT_UOUT5
  PIN UIO_BOT_UOUT6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.920 0.000 151.300 0.700 ;
    END
  END UIO_BOT_UOUT6
  PIN UIO_BOT_UOUT7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 155.060 0.000 155.440 0.700 ;
    END
  END UIO_BOT_UOUT7
  PIN UIO_BOT_UOUT8
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 158.740 0.000 159.120 0.700 ;
    END
  END UIO_BOT_UOUT8
  PIN UIO_BOT_UOUT9
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.880 0.000 163.260 0.700 ;
    END
  END UIO_BOT_UOUT9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 0.700 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.580 5.200 22.180 177.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 5.200 175.780 177.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 21.290 244.960 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 174.470 244.960 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.880 5.200 25.480 177.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.480 5.200 179.080 177.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.820 24.590 244.960 26.190 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.060 5.355 244.720 176.885 ;
      LAYER met1 ;
        RECT 5.060 2.420 244.720 179.140 ;
      LAYER met2 ;
        RECT 4.380 181.020 5.280 181.300 ;
        RECT 6.220 181.020 7.120 181.300 ;
        RECT 8.060 181.020 8.960 181.300 ;
        RECT 9.900 181.020 10.800 181.300 ;
        RECT 11.740 181.020 13.100 181.300 ;
        RECT 14.040 181.020 14.940 181.300 ;
        RECT 15.880 181.020 16.780 181.300 ;
        RECT 17.720 181.020 18.620 181.300 ;
        RECT 19.560 181.020 20.460 181.300 ;
        RECT 21.400 181.020 22.300 181.300 ;
        RECT 23.240 181.020 24.600 181.300 ;
        RECT 25.540 181.020 26.440 181.300 ;
        RECT 27.380 181.020 28.280 181.300 ;
        RECT 29.220 181.020 30.120 181.300 ;
        RECT 31.060 181.020 31.960 181.300 ;
        RECT 32.900 181.020 34.260 181.300 ;
        RECT 35.200 181.020 36.100 181.300 ;
        RECT 37.040 181.020 37.940 181.300 ;
        RECT 38.880 181.020 39.780 181.300 ;
        RECT 40.720 181.020 41.620 181.300 ;
        RECT 42.560 181.020 43.920 181.300 ;
        RECT 44.860 181.020 45.760 181.300 ;
        RECT 46.700 181.020 47.600 181.300 ;
        RECT 48.540 181.020 49.440 181.300 ;
        RECT 50.380 181.020 51.280 181.300 ;
        RECT 52.220 181.020 53.580 181.300 ;
        RECT 54.520 181.020 55.420 181.300 ;
        RECT 56.360 181.020 57.260 181.300 ;
        RECT 58.200 181.020 59.100 181.300 ;
        RECT 60.040 181.020 60.940 181.300 ;
        RECT 61.880 181.020 63.240 181.300 ;
        RECT 64.180 181.020 65.080 181.300 ;
        RECT 66.020 181.020 66.920 181.300 ;
        RECT 67.860 181.020 68.760 181.300 ;
        RECT 69.700 181.020 70.600 181.300 ;
        RECT 71.540 181.020 72.900 181.300 ;
        RECT 73.840 181.020 74.740 181.300 ;
        RECT 75.680 181.020 76.580 181.300 ;
        RECT 77.520 181.020 78.420 181.300 ;
        RECT 79.360 181.020 80.260 181.300 ;
        RECT 81.200 181.020 82.100 181.300 ;
        RECT 83.040 181.020 84.400 181.300 ;
        RECT 85.340 181.020 86.240 181.300 ;
        RECT 87.180 181.020 88.080 181.300 ;
        RECT 89.020 181.020 89.920 181.300 ;
        RECT 90.860 181.020 91.760 181.300 ;
        RECT 92.700 181.020 94.060 181.300 ;
        RECT 95.000 181.020 95.900 181.300 ;
        RECT 96.840 181.020 97.740 181.300 ;
        RECT 98.680 181.020 99.580 181.300 ;
        RECT 100.520 181.020 101.420 181.300 ;
        RECT 102.360 181.020 103.720 181.300 ;
        RECT 104.660 181.020 105.560 181.300 ;
        RECT 106.500 181.020 107.400 181.300 ;
        RECT 108.340 181.020 109.240 181.300 ;
        RECT 110.180 181.020 111.080 181.300 ;
        RECT 112.020 181.020 113.380 181.300 ;
        RECT 114.320 181.020 115.220 181.300 ;
        RECT 116.160 181.020 117.060 181.300 ;
        RECT 118.000 181.020 118.900 181.300 ;
        RECT 119.840 181.020 120.740 181.300 ;
        RECT 121.680 181.020 123.040 181.300 ;
        RECT 123.980 181.020 124.880 181.300 ;
        RECT 125.820 181.020 126.720 181.300 ;
        RECT 127.660 181.020 128.560 181.300 ;
        RECT 129.500 181.020 130.400 181.300 ;
        RECT 131.340 181.020 132.700 181.300 ;
        RECT 133.640 181.020 134.540 181.300 ;
        RECT 135.480 181.020 136.380 181.300 ;
        RECT 137.320 181.020 138.220 181.300 ;
        RECT 139.160 181.020 140.060 181.300 ;
        RECT 141.000 181.020 141.900 181.300 ;
        RECT 142.840 181.020 144.200 181.300 ;
        RECT 145.140 181.020 146.040 181.300 ;
        RECT 146.980 181.020 147.880 181.300 ;
        RECT 148.820 181.020 149.720 181.300 ;
        RECT 150.660 181.020 151.560 181.300 ;
        RECT 152.500 181.020 153.860 181.300 ;
        RECT 154.800 181.020 155.700 181.300 ;
        RECT 156.640 181.020 157.540 181.300 ;
        RECT 158.480 181.020 159.380 181.300 ;
        RECT 160.320 181.020 161.220 181.300 ;
        RECT 162.160 181.020 163.520 181.300 ;
        RECT 164.460 181.020 165.360 181.300 ;
        RECT 166.300 181.020 167.200 181.300 ;
        RECT 168.140 181.020 169.040 181.300 ;
        RECT 169.980 181.020 170.880 181.300 ;
        RECT 171.820 181.020 173.180 181.300 ;
        RECT 174.120 181.020 175.020 181.300 ;
        RECT 175.960 181.020 176.860 181.300 ;
        RECT 177.800 181.020 178.700 181.300 ;
        RECT 179.640 181.020 180.540 181.300 ;
        RECT 181.480 181.020 182.840 181.300 ;
        RECT 183.780 181.020 184.680 181.300 ;
        RECT 185.620 181.020 186.520 181.300 ;
        RECT 187.460 181.020 188.360 181.300 ;
        RECT 189.300 181.020 190.200 181.300 ;
        RECT 191.140 181.020 192.500 181.300 ;
        RECT 193.440 181.020 194.340 181.300 ;
        RECT 195.280 181.020 196.180 181.300 ;
        RECT 197.120 181.020 198.020 181.300 ;
        RECT 198.960 181.020 199.860 181.300 ;
        RECT 200.800 181.020 201.700 181.300 ;
        RECT 202.640 181.020 204.000 181.300 ;
        RECT 204.940 181.020 205.840 181.300 ;
        RECT 206.780 181.020 207.680 181.300 ;
        RECT 208.620 181.020 209.520 181.300 ;
        RECT 210.460 181.020 211.360 181.300 ;
        RECT 212.300 181.020 213.660 181.300 ;
        RECT 214.600 181.020 215.500 181.300 ;
        RECT 216.440 181.020 217.340 181.300 ;
        RECT 218.280 181.020 219.180 181.300 ;
        RECT 220.120 181.020 221.020 181.300 ;
        RECT 221.960 181.020 223.320 181.300 ;
        RECT 224.260 181.020 225.160 181.300 ;
        RECT 226.100 181.020 227.000 181.300 ;
        RECT 227.940 181.020 228.840 181.300 ;
        RECT 229.780 181.020 230.680 181.300 ;
        RECT 231.620 181.020 232.980 181.300 ;
        RECT 233.920 181.020 234.820 181.300 ;
        RECT 235.760 181.020 236.660 181.300 ;
        RECT 237.600 181.020 238.500 181.300 ;
        RECT 239.440 181.020 240.340 181.300 ;
        RECT 241.280 181.020 242.640 181.300 ;
        RECT 243.580 181.020 243.700 181.300 ;
        RECT 3.840 0.980 243.700 181.020 ;
        RECT 3.840 0.270 5.280 0.980 ;
        RECT 6.220 0.270 9.420 0.980 ;
        RECT 10.360 0.270 13.560 0.980 ;
        RECT 14.500 0.270 17.240 0.980 ;
        RECT 18.180 0.270 21.380 0.980 ;
        RECT 22.320 0.270 25.520 0.980 ;
        RECT 26.460 0.270 29.660 0.980 ;
        RECT 30.600 0.270 33.340 0.980 ;
        RECT 34.280 0.270 37.480 0.980 ;
        RECT 38.420 0.270 41.620 0.980 ;
        RECT 42.560 0.270 45.760 0.980 ;
        RECT 46.700 0.270 49.900 0.980 ;
        RECT 50.840 0.270 53.580 0.980 ;
        RECT 54.520 0.270 57.720 0.980 ;
        RECT 58.660 0.270 61.860 0.980 ;
        RECT 62.800 0.270 66.000 0.980 ;
        RECT 66.940 0.270 69.680 0.980 ;
        RECT 70.620 0.270 73.820 0.980 ;
        RECT 74.760 0.270 77.960 0.980 ;
        RECT 78.900 0.270 82.100 0.980 ;
        RECT 83.040 0.270 85.780 0.980 ;
        RECT 86.720 0.270 89.920 0.980 ;
        RECT 90.860 0.270 94.060 0.980 ;
        RECT 95.000 0.270 98.200 0.980 ;
        RECT 99.140 0.270 102.340 0.980 ;
        RECT 103.280 0.270 106.020 0.980 ;
        RECT 106.960 0.270 109.290 0.980 ;
        RECT 110.130 0.270 110.160 0.980 ;
        RECT 111.100 0.270 112.510 0.980 ;
        RECT 113.350 0.270 114.300 0.980 ;
        RECT 115.240 0.270 118.440 0.980 ;
        RECT 119.380 0.270 122.120 0.980 ;
        RECT 123.060 0.270 126.260 0.980 ;
        RECT 127.200 0.270 130.400 0.980 ;
        RECT 131.340 0.270 134.540 0.980 ;
        RECT 135.480 0.270 138.220 0.980 ;
        RECT 139.160 0.270 142.360 0.980 ;
        RECT 143.300 0.270 146.500 0.980 ;
        RECT 147.440 0.270 150.640 0.980 ;
        RECT 151.580 0.270 154.780 0.980 ;
        RECT 155.720 0.270 158.460 0.980 ;
        RECT 159.400 0.270 162.600 0.980 ;
        RECT 163.540 0.270 166.740 0.980 ;
        RECT 167.680 0.270 170.880 0.980 ;
        RECT 171.820 0.270 174.560 0.980 ;
        RECT 175.500 0.270 178.700 0.980 ;
        RECT 179.640 0.270 182.840 0.980 ;
        RECT 183.780 0.270 186.980 0.980 ;
        RECT 187.920 0.270 190.660 0.980 ;
        RECT 191.600 0.270 194.800 0.980 ;
        RECT 195.740 0.270 198.940 0.980 ;
        RECT 199.880 0.270 203.080 0.980 ;
        RECT 204.020 0.270 206.760 0.980 ;
        RECT 207.700 0.270 210.900 0.980 ;
        RECT 211.840 0.270 215.040 0.980 ;
        RECT 215.980 0.270 219.180 0.980 ;
        RECT 220.120 0.270 223.320 0.980 ;
        RECT 224.260 0.270 227.000 0.980 ;
        RECT 227.940 0.270 231.140 0.980 ;
        RECT 232.080 0.270 235.280 0.980 ;
        RECT 236.220 0.270 239.420 0.980 ;
        RECT 240.360 0.270 243.100 0.980 ;
      LAYER met3 ;
        RECT 20.590 5.275 209.235 176.965 ;
      LAYER met4 ;
        RECT 113.455 38.935 128.505 110.665 ;
  END
END S_term_single
END LIBRARY

