module LUT4AB (Ci,
    Co,
    UserCLK,
    UserCLKo,
    vccd1,
    vssd1,
    E1BEG,
    E1END,
    E2BEG,
    E2BEGb,
    E2END,
    E2MID,
    E6BEG,
    E6END,
    EE4BEG,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    NN4BEG,
    NN4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    SS4BEG,
    SS4END,
    W1BEG,
    W1END,
    W2BEG,
    W2BEGb,
    W2END,
    W2MID,
    W6BEG,
    W6END,
    WW4BEG,
    WW4END);
 input Ci;
 output Co;
 input UserCLK;
 output UserCLKo;
 input vccd1;
 input vssd1;
 output [3:0] E1BEG;
 input [3:0] E1END;
 output [7:0] E2BEG;
 output [7:0] E2BEGb;
 input [7:0] E2END;
 input [7:0] E2MID;
 output [11:0] E6BEG;
 input [11:0] E6END;
 output [15:0] EE4BEG;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [15:0] NN4BEG;
 input [15:0] NN4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [15:0] SS4BEG;
 input [15:0] SS4END;
 output [3:0] W1BEG;
 input [3:0] W1END;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 input [7:0] W2END;
 input [7:0] W2MID;
 output [11:0] W6BEG;
 input [11:0] W6END;
 output [15:0] WW4BEG;
 input [15:0] WW4END;

 wire A;
 wire B;
 wire C;
 wire \ConfigBits[0] ;
 wire \ConfigBits[100] ;
 wire \ConfigBits[101] ;
 wire \ConfigBits[102] ;
 wire \ConfigBits[103] ;
 wire \ConfigBits[104] ;
 wire \ConfigBits[105] ;
 wire \ConfigBits[106] ;
 wire \ConfigBits[107] ;
 wire \ConfigBits[108] ;
 wire \ConfigBits[109] ;
 wire \ConfigBits[10] ;
 wire \ConfigBits[110] ;
 wire \ConfigBits[111] ;
 wire \ConfigBits[112] ;
 wire \ConfigBits[113] ;
 wire \ConfigBits[114] ;
 wire \ConfigBits[115] ;
 wire \ConfigBits[116] ;
 wire \ConfigBits[117] ;
 wire \ConfigBits[118] ;
 wire \ConfigBits[119] ;
 wire \ConfigBits[11] ;
 wire \ConfigBits[120] ;
 wire \ConfigBits[121] ;
 wire \ConfigBits[122] ;
 wire \ConfigBits[123] ;
 wire \ConfigBits[124] ;
 wire \ConfigBits[125] ;
 wire \ConfigBits[126] ;
 wire \ConfigBits[127] ;
 wire \ConfigBits[128] ;
 wire \ConfigBits[129] ;
 wire \ConfigBits[12] ;
 wire \ConfigBits[130] ;
 wire \ConfigBits[131] ;
 wire \ConfigBits[132] ;
 wire \ConfigBits[133] ;
 wire \ConfigBits[134] ;
 wire \ConfigBits[135] ;
 wire \ConfigBits[136] ;
 wire \ConfigBits[137] ;
 wire \ConfigBits[138] ;
 wire \ConfigBits[139] ;
 wire \ConfigBits[13] ;
 wire \ConfigBits[140] ;
 wire \ConfigBits[141] ;
 wire \ConfigBits[142] ;
 wire \ConfigBits[143] ;
 wire \ConfigBits[144] ;
 wire \ConfigBits[145] ;
 wire \ConfigBits[146] ;
 wire \ConfigBits[147] ;
 wire \ConfigBits[148] ;
 wire \ConfigBits[149] ;
 wire \ConfigBits[14] ;
 wire \ConfigBits[150] ;
 wire \ConfigBits[151] ;
 wire \ConfigBits[152] ;
 wire \ConfigBits[153] ;
 wire \ConfigBits[154] ;
 wire \ConfigBits[155] ;
 wire \ConfigBits[156] ;
 wire \ConfigBits[157] ;
 wire \ConfigBits[158] ;
 wire \ConfigBits[159] ;
 wire \ConfigBits[15] ;
 wire \ConfigBits[160] ;
 wire \ConfigBits[161] ;
 wire \ConfigBits[162] ;
 wire \ConfigBits[163] ;
 wire \ConfigBits[164] ;
 wire \ConfigBits[165] ;
 wire \ConfigBits[166] ;
 wire \ConfigBits[167] ;
 wire \ConfigBits[168] ;
 wire \ConfigBits[169] ;
 wire \ConfigBits[16] ;
 wire \ConfigBits[170] ;
 wire \ConfigBits[171] ;
 wire \ConfigBits[172] ;
 wire \ConfigBits[173] ;
 wire \ConfigBits[174] ;
 wire \ConfigBits[175] ;
 wire \ConfigBits[176] ;
 wire \ConfigBits[177] ;
 wire \ConfigBits[178] ;
 wire \ConfigBits[179] ;
 wire \ConfigBits[17] ;
 wire \ConfigBits[180] ;
 wire \ConfigBits[181] ;
 wire \ConfigBits[182] ;
 wire \ConfigBits[183] ;
 wire \ConfigBits[184] ;
 wire \ConfigBits[185] ;
 wire \ConfigBits[186] ;
 wire \ConfigBits[187] ;
 wire \ConfigBits[188] ;
 wire \ConfigBits[189] ;
 wire \ConfigBits[18] ;
 wire \ConfigBits[190] ;
 wire \ConfigBits[191] ;
 wire \ConfigBits[192] ;
 wire \ConfigBits[193] ;
 wire \ConfigBits[194] ;
 wire \ConfigBits[195] ;
 wire \ConfigBits[196] ;
 wire \ConfigBits[197] ;
 wire \ConfigBits[198] ;
 wire \ConfigBits[199] ;
 wire \ConfigBits[19] ;
 wire \ConfigBits[1] ;
 wire \ConfigBits[200] ;
 wire \ConfigBits[201] ;
 wire \ConfigBits[202] ;
 wire \ConfigBits[203] ;
 wire \ConfigBits[204] ;
 wire \ConfigBits[205] ;
 wire \ConfigBits[206] ;
 wire \ConfigBits[207] ;
 wire \ConfigBits[208] ;
 wire \ConfigBits[209] ;
 wire \ConfigBits[20] ;
 wire \ConfigBits[210] ;
 wire \ConfigBits[211] ;
 wire \ConfigBits[212] ;
 wire \ConfigBits[213] ;
 wire \ConfigBits[214] ;
 wire \ConfigBits[215] ;
 wire \ConfigBits[216] ;
 wire \ConfigBits[217] ;
 wire \ConfigBits[218] ;
 wire \ConfigBits[219] ;
 wire \ConfigBits[21] ;
 wire \ConfigBits[220] ;
 wire \ConfigBits[221] ;
 wire \ConfigBits[222] ;
 wire \ConfigBits[223] ;
 wire \ConfigBits[224] ;
 wire \ConfigBits[225] ;
 wire \ConfigBits[226] ;
 wire \ConfigBits[227] ;
 wire \ConfigBits[228] ;
 wire \ConfigBits[229] ;
 wire \ConfigBits[22] ;
 wire \ConfigBits[230] ;
 wire \ConfigBits[231] ;
 wire \ConfigBits[232] ;
 wire \ConfigBits[233] ;
 wire \ConfigBits[234] ;
 wire \ConfigBits[235] ;
 wire \ConfigBits[236] ;
 wire \ConfigBits[237] ;
 wire \ConfigBits[238] ;
 wire \ConfigBits[239] ;
 wire \ConfigBits[23] ;
 wire \ConfigBits[240] ;
 wire \ConfigBits[241] ;
 wire \ConfigBits[242] ;
 wire \ConfigBits[243] ;
 wire \ConfigBits[244] ;
 wire \ConfigBits[245] ;
 wire \ConfigBits[246] ;
 wire \ConfigBits[247] ;
 wire \ConfigBits[248] ;
 wire \ConfigBits[249] ;
 wire \ConfigBits[24] ;
 wire \ConfigBits[250] ;
 wire \ConfigBits[251] ;
 wire \ConfigBits[252] ;
 wire \ConfigBits[253] ;
 wire \ConfigBits[254] ;
 wire \ConfigBits[255] ;
 wire \ConfigBits[256] ;
 wire \ConfigBits[257] ;
 wire \ConfigBits[258] ;
 wire \ConfigBits[259] ;
 wire \ConfigBits[25] ;
 wire \ConfigBits[260] ;
 wire \ConfigBits[261] ;
 wire \ConfigBits[262] ;
 wire \ConfigBits[263] ;
 wire \ConfigBits[264] ;
 wire \ConfigBits[265] ;
 wire \ConfigBits[266] ;
 wire \ConfigBits[267] ;
 wire \ConfigBits[268] ;
 wire \ConfigBits[269] ;
 wire \ConfigBits[26] ;
 wire \ConfigBits[270] ;
 wire \ConfigBits[271] ;
 wire \ConfigBits[272] ;
 wire \ConfigBits[273] ;
 wire \ConfigBits[274] ;
 wire \ConfigBits[275] ;
 wire \ConfigBits[276] ;
 wire \ConfigBits[277] ;
 wire \ConfigBits[278] ;
 wire \ConfigBits[279] ;
 wire \ConfigBits[27] ;
 wire \ConfigBits[280] ;
 wire \ConfigBits[281] ;
 wire \ConfigBits[282] ;
 wire \ConfigBits[283] ;
 wire \ConfigBits[284] ;
 wire \ConfigBits[285] ;
 wire \ConfigBits[286] ;
 wire \ConfigBits[287] ;
 wire \ConfigBits[288] ;
 wire \ConfigBits[289] ;
 wire \ConfigBits[28] ;
 wire \ConfigBits[290] ;
 wire \ConfigBits[291] ;
 wire \ConfigBits[292] ;
 wire \ConfigBits[293] ;
 wire \ConfigBits[294] ;
 wire \ConfigBits[295] ;
 wire \ConfigBits[296] ;
 wire \ConfigBits[297] ;
 wire \ConfigBits[298] ;
 wire \ConfigBits[299] ;
 wire \ConfigBits[29] ;
 wire \ConfigBits[2] ;
 wire \ConfigBits[300] ;
 wire \ConfigBits[301] ;
 wire \ConfigBits[302] ;
 wire \ConfigBits[303] ;
 wire \ConfigBits[304] ;
 wire \ConfigBits[305] ;
 wire \ConfigBits[306] ;
 wire \ConfigBits[307] ;
 wire \ConfigBits[308] ;
 wire \ConfigBits[309] ;
 wire \ConfigBits[30] ;
 wire \ConfigBits[310] ;
 wire \ConfigBits[311] ;
 wire \ConfigBits[312] ;
 wire \ConfigBits[313] ;
 wire \ConfigBits[314] ;
 wire \ConfigBits[315] ;
 wire \ConfigBits[316] ;
 wire \ConfigBits[317] ;
 wire \ConfigBits[318] ;
 wire \ConfigBits[319] ;
 wire \ConfigBits[31] ;
 wire \ConfigBits[320] ;
 wire \ConfigBits[321] ;
 wire \ConfigBits[322] ;
 wire \ConfigBits[323] ;
 wire \ConfigBits[324] ;
 wire \ConfigBits[325] ;
 wire \ConfigBits[326] ;
 wire \ConfigBits[327] ;
 wire \ConfigBits[328] ;
 wire \ConfigBits[329] ;
 wire \ConfigBits[32] ;
 wire \ConfigBits[330] ;
 wire \ConfigBits[331] ;
 wire \ConfigBits[332] ;
 wire \ConfigBits[333] ;
 wire \ConfigBits[334] ;
 wire \ConfigBits[335] ;
 wire \ConfigBits[336] ;
 wire \ConfigBits[337] ;
 wire \ConfigBits[338] ;
 wire \ConfigBits[339] ;
 wire \ConfigBits[33] ;
 wire \ConfigBits[340] ;
 wire \ConfigBits[341] ;
 wire \ConfigBits[342] ;
 wire \ConfigBits[343] ;
 wire \ConfigBits[344] ;
 wire \ConfigBits[345] ;
 wire \ConfigBits[346] ;
 wire \ConfigBits[347] ;
 wire \ConfigBits[348] ;
 wire \ConfigBits[349] ;
 wire \ConfigBits[34] ;
 wire \ConfigBits[350] ;
 wire \ConfigBits[351] ;
 wire \ConfigBits[352] ;
 wire \ConfigBits[353] ;
 wire \ConfigBits[354] ;
 wire \ConfigBits[355] ;
 wire \ConfigBits[356] ;
 wire \ConfigBits[357] ;
 wire \ConfigBits[358] ;
 wire \ConfigBits[359] ;
 wire \ConfigBits[35] ;
 wire \ConfigBits[360] ;
 wire \ConfigBits[361] ;
 wire \ConfigBits[362] ;
 wire \ConfigBits[363] ;
 wire \ConfigBits[364] ;
 wire \ConfigBits[365] ;
 wire \ConfigBits[366] ;
 wire \ConfigBits[367] ;
 wire \ConfigBits[368] ;
 wire \ConfigBits[369] ;
 wire \ConfigBits[36] ;
 wire \ConfigBits[370] ;
 wire \ConfigBits[371] ;
 wire \ConfigBits[372] ;
 wire \ConfigBits[373] ;
 wire \ConfigBits[374] ;
 wire \ConfigBits[375] ;
 wire \ConfigBits[376] ;
 wire \ConfigBits[377] ;
 wire \ConfigBits[378] ;
 wire \ConfigBits[379] ;
 wire \ConfigBits[37] ;
 wire \ConfigBits[380] ;
 wire \ConfigBits[381] ;
 wire \ConfigBits[382] ;
 wire \ConfigBits[383] ;
 wire \ConfigBits[384] ;
 wire \ConfigBits[385] ;
 wire \ConfigBits[386] ;
 wire \ConfigBits[387] ;
 wire \ConfigBits[388] ;
 wire \ConfigBits[389] ;
 wire \ConfigBits[38] ;
 wire \ConfigBits[390] ;
 wire \ConfigBits[391] ;
 wire \ConfigBits[392] ;
 wire \ConfigBits[393] ;
 wire \ConfigBits[394] ;
 wire \ConfigBits[395] ;
 wire \ConfigBits[396] ;
 wire \ConfigBits[397] ;
 wire \ConfigBits[398] ;
 wire \ConfigBits[399] ;
 wire \ConfigBits[39] ;
 wire \ConfigBits[3] ;
 wire \ConfigBits[400] ;
 wire \ConfigBits[401] ;
 wire \ConfigBits[402] ;
 wire \ConfigBits[403] ;
 wire \ConfigBits[404] ;
 wire \ConfigBits[405] ;
 wire \ConfigBits[406] ;
 wire \ConfigBits[407] ;
 wire \ConfigBits[408] ;
 wire \ConfigBits[409] ;
 wire \ConfigBits[40] ;
 wire \ConfigBits[410] ;
 wire \ConfigBits[411] ;
 wire \ConfigBits[412] ;
 wire \ConfigBits[413] ;
 wire \ConfigBits[414] ;
 wire \ConfigBits[415] ;
 wire \ConfigBits[416] ;
 wire \ConfigBits[417] ;
 wire \ConfigBits[418] ;
 wire \ConfigBits[419] ;
 wire \ConfigBits[41] ;
 wire \ConfigBits[420] ;
 wire \ConfigBits[421] ;
 wire \ConfigBits[422] ;
 wire \ConfigBits[423] ;
 wire \ConfigBits[424] ;
 wire \ConfigBits[425] ;
 wire \ConfigBits[426] ;
 wire \ConfigBits[427] ;
 wire \ConfigBits[428] ;
 wire \ConfigBits[429] ;
 wire \ConfigBits[42] ;
 wire \ConfigBits[430] ;
 wire \ConfigBits[431] ;
 wire \ConfigBits[432] ;
 wire \ConfigBits[433] ;
 wire \ConfigBits[434] ;
 wire \ConfigBits[435] ;
 wire \ConfigBits[436] ;
 wire \ConfigBits[437] ;
 wire \ConfigBits[438] ;
 wire \ConfigBits[439] ;
 wire \ConfigBits[43] ;
 wire \ConfigBits[440] ;
 wire \ConfigBits[441] ;
 wire \ConfigBits[442] ;
 wire \ConfigBits[443] ;
 wire \ConfigBits[444] ;
 wire \ConfigBits[445] ;
 wire \ConfigBits[446] ;
 wire \ConfigBits[447] ;
 wire \ConfigBits[448] ;
 wire \ConfigBits[449] ;
 wire \ConfigBits[44] ;
 wire \ConfigBits[450] ;
 wire \ConfigBits[451] ;
 wire \ConfigBits[452] ;
 wire \ConfigBits[453] ;
 wire \ConfigBits[454] ;
 wire \ConfigBits[455] ;
 wire \ConfigBits[456] ;
 wire \ConfigBits[457] ;
 wire \ConfigBits[458] ;
 wire \ConfigBits[459] ;
 wire \ConfigBits[45] ;
 wire \ConfigBits[460] ;
 wire \ConfigBits[461] ;
 wire \ConfigBits[462] ;
 wire \ConfigBits[463] ;
 wire \ConfigBits[464] ;
 wire \ConfigBits[465] ;
 wire \ConfigBits[466] ;
 wire \ConfigBits[467] ;
 wire \ConfigBits[468] ;
 wire \ConfigBits[469] ;
 wire \ConfigBits[46] ;
 wire \ConfigBits[470] ;
 wire \ConfigBits[471] ;
 wire \ConfigBits[472] ;
 wire \ConfigBits[473] ;
 wire \ConfigBits[474] ;
 wire \ConfigBits[475] ;
 wire \ConfigBits[476] ;
 wire \ConfigBits[477] ;
 wire \ConfigBits[478] ;
 wire \ConfigBits[479] ;
 wire \ConfigBits[47] ;
 wire \ConfigBits[480] ;
 wire \ConfigBits[481] ;
 wire \ConfigBits[482] ;
 wire \ConfigBits[483] ;
 wire \ConfigBits[484] ;
 wire \ConfigBits[485] ;
 wire \ConfigBits[486] ;
 wire \ConfigBits[487] ;
 wire \ConfigBits[488] ;
 wire \ConfigBits[489] ;
 wire \ConfigBits[48] ;
 wire \ConfigBits[490] ;
 wire \ConfigBits[491] ;
 wire \ConfigBits[492] ;
 wire \ConfigBits[493] ;
 wire \ConfigBits[494] ;
 wire \ConfigBits[495] ;
 wire \ConfigBits[496] ;
 wire \ConfigBits[497] ;
 wire \ConfigBits[498] ;
 wire \ConfigBits[499] ;
 wire \ConfigBits[49] ;
 wire \ConfigBits[4] ;
 wire \ConfigBits[500] ;
 wire \ConfigBits[501] ;
 wire \ConfigBits[502] ;
 wire \ConfigBits[503] ;
 wire \ConfigBits[504] ;
 wire \ConfigBits[505] ;
 wire \ConfigBits[506] ;
 wire \ConfigBits[507] ;
 wire \ConfigBits[508] ;
 wire \ConfigBits[509] ;
 wire \ConfigBits[50] ;
 wire \ConfigBits[510] ;
 wire \ConfigBits[511] ;
 wire \ConfigBits[512] ;
 wire \ConfigBits[513] ;
 wire \ConfigBits[514] ;
 wire \ConfigBits[515] ;
 wire \ConfigBits[516] ;
 wire \ConfigBits[517] ;
 wire \ConfigBits[518] ;
 wire \ConfigBits[519] ;
 wire \ConfigBits[51] ;
 wire \ConfigBits[520] ;
 wire \ConfigBits[521] ;
 wire \ConfigBits[522] ;
 wire \ConfigBits[523] ;
 wire \ConfigBits[524] ;
 wire \ConfigBits[525] ;
 wire \ConfigBits[526] ;
 wire \ConfigBits[527] ;
 wire \ConfigBits[528] ;
 wire \ConfigBits[529] ;
 wire \ConfigBits[52] ;
 wire \ConfigBits[530] ;
 wire \ConfigBits[531] ;
 wire \ConfigBits[532] ;
 wire \ConfigBits[533] ;
 wire \ConfigBits[534] ;
 wire \ConfigBits[535] ;
 wire \ConfigBits[536] ;
 wire \ConfigBits[537] ;
 wire \ConfigBits[538] ;
 wire \ConfigBits[539] ;
 wire \ConfigBits[53] ;
 wire \ConfigBits[540] ;
 wire \ConfigBits[541] ;
 wire \ConfigBits[542] ;
 wire \ConfigBits[543] ;
 wire \ConfigBits[544] ;
 wire \ConfigBits[545] ;
 wire \ConfigBits[546] ;
 wire \ConfigBits[547] ;
 wire \ConfigBits[548] ;
 wire \ConfigBits[549] ;
 wire \ConfigBits[54] ;
 wire \ConfigBits[550] ;
 wire \ConfigBits[551] ;
 wire \ConfigBits[552] ;
 wire \ConfigBits[553] ;
 wire \ConfigBits[554] ;
 wire \ConfigBits[555] ;
 wire \ConfigBits[556] ;
 wire \ConfigBits[557] ;
 wire \ConfigBits[558] ;
 wire \ConfigBits[559] ;
 wire \ConfigBits[55] ;
 wire \ConfigBits[560] ;
 wire \ConfigBits[561] ;
 wire \ConfigBits[562] ;
 wire \ConfigBits[563] ;
 wire \ConfigBits[564] ;
 wire \ConfigBits[565] ;
 wire \ConfigBits[566] ;
 wire \ConfigBits[567] ;
 wire \ConfigBits[568] ;
 wire \ConfigBits[569] ;
 wire \ConfigBits[56] ;
 wire \ConfigBits[570] ;
 wire \ConfigBits[571] ;
 wire \ConfigBits[572] ;
 wire \ConfigBits[573] ;
 wire \ConfigBits[574] ;
 wire \ConfigBits[575] ;
 wire \ConfigBits[576] ;
 wire \ConfigBits[577] ;
 wire \ConfigBits[578] ;
 wire \ConfigBits[579] ;
 wire \ConfigBits[57] ;
 wire \ConfigBits[580] ;
 wire \ConfigBits[581] ;
 wire \ConfigBits[582] ;
 wire \ConfigBits[583] ;
 wire \ConfigBits[584] ;
 wire \ConfigBits[585] ;
 wire \ConfigBits[586] ;
 wire \ConfigBits[587] ;
 wire \ConfigBits[588] ;
 wire \ConfigBits[589] ;
 wire \ConfigBits[58] ;
 wire \ConfigBits[590] ;
 wire \ConfigBits[591] ;
 wire \ConfigBits[592] ;
 wire \ConfigBits[593] ;
 wire \ConfigBits[594] ;
 wire \ConfigBits[595] ;
 wire \ConfigBits[596] ;
 wire \ConfigBits[597] ;
 wire \ConfigBits[598] ;
 wire \ConfigBits[599] ;
 wire \ConfigBits[59] ;
 wire \ConfigBits[5] ;
 wire \ConfigBits[600] ;
 wire \ConfigBits[601] ;
 wire \ConfigBits[602] ;
 wire \ConfigBits[603] ;
 wire \ConfigBits[604] ;
 wire \ConfigBits[605] ;
 wire \ConfigBits[606] ;
 wire \ConfigBits[607] ;
 wire \ConfigBits[608] ;
 wire \ConfigBits[609] ;
 wire \ConfigBits[60] ;
 wire \ConfigBits[610] ;
 wire \ConfigBits[611] ;
 wire \ConfigBits[612] ;
 wire \ConfigBits[613] ;
 wire \ConfigBits[614] ;
 wire \ConfigBits[615] ;
 wire \ConfigBits[61] ;
 wire \ConfigBits[62] ;
 wire \ConfigBits[63] ;
 wire \ConfigBits[64] ;
 wire \ConfigBits[65] ;
 wire \ConfigBits[66] ;
 wire \ConfigBits[67] ;
 wire \ConfigBits[68] ;
 wire \ConfigBits[69] ;
 wire \ConfigBits[6] ;
 wire \ConfigBits[70] ;
 wire \ConfigBits[71] ;
 wire \ConfigBits[72] ;
 wire \ConfigBits[73] ;
 wire \ConfigBits[74] ;
 wire \ConfigBits[75] ;
 wire \ConfigBits[76] ;
 wire \ConfigBits[77] ;
 wire \ConfigBits[78] ;
 wire \ConfigBits[79] ;
 wire \ConfigBits[7] ;
 wire \ConfigBits[80] ;
 wire \ConfigBits[81] ;
 wire \ConfigBits[82] ;
 wire \ConfigBits[83] ;
 wire \ConfigBits[84] ;
 wire \ConfigBits[85] ;
 wire \ConfigBits[86] ;
 wire \ConfigBits[87] ;
 wire \ConfigBits[88] ;
 wire \ConfigBits[89] ;
 wire \ConfigBits[8] ;
 wire \ConfigBits[90] ;
 wire \ConfigBits[91] ;
 wire \ConfigBits[92] ;
 wire \ConfigBits[93] ;
 wire \ConfigBits[94] ;
 wire \ConfigBits[95] ;
 wire \ConfigBits[96] ;
 wire \ConfigBits[97] ;
 wire \ConfigBits[98] ;
 wire \ConfigBits[99] ;
 wire \ConfigBits[9] ;
 wire \ConfigBits_N[0] ;
 wire \ConfigBits_N[100] ;
 wire \ConfigBits_N[101] ;
 wire \ConfigBits_N[102] ;
 wire \ConfigBits_N[103] ;
 wire \ConfigBits_N[104] ;
 wire \ConfigBits_N[105] ;
 wire \ConfigBits_N[106] ;
 wire \ConfigBits_N[107] ;
 wire \ConfigBits_N[108] ;
 wire \ConfigBits_N[109] ;
 wire \ConfigBits_N[10] ;
 wire \ConfigBits_N[110] ;
 wire \ConfigBits_N[111] ;
 wire \ConfigBits_N[112] ;
 wire \ConfigBits_N[113] ;
 wire \ConfigBits_N[114] ;
 wire \ConfigBits_N[115] ;
 wire \ConfigBits_N[116] ;
 wire \ConfigBits_N[117] ;
 wire \ConfigBits_N[118] ;
 wire \ConfigBits_N[119] ;
 wire \ConfigBits_N[11] ;
 wire \ConfigBits_N[120] ;
 wire \ConfigBits_N[121] ;
 wire \ConfigBits_N[122] ;
 wire \ConfigBits_N[123] ;
 wire \ConfigBits_N[124] ;
 wire \ConfigBits_N[125] ;
 wire \ConfigBits_N[126] ;
 wire \ConfigBits_N[127] ;
 wire \ConfigBits_N[128] ;
 wire \ConfigBits_N[129] ;
 wire \ConfigBits_N[12] ;
 wire \ConfigBits_N[130] ;
 wire \ConfigBits_N[131] ;
 wire \ConfigBits_N[132] ;
 wire \ConfigBits_N[133] ;
 wire \ConfigBits_N[134] ;
 wire \ConfigBits_N[135] ;
 wire \ConfigBits_N[136] ;
 wire \ConfigBits_N[137] ;
 wire \ConfigBits_N[138] ;
 wire \ConfigBits_N[139] ;
 wire \ConfigBits_N[13] ;
 wire \ConfigBits_N[140] ;
 wire \ConfigBits_N[141] ;
 wire \ConfigBits_N[142] ;
 wire \ConfigBits_N[143] ;
 wire \ConfigBits_N[144] ;
 wire \ConfigBits_N[145] ;
 wire \ConfigBits_N[146] ;
 wire \ConfigBits_N[147] ;
 wire \ConfigBits_N[148] ;
 wire \ConfigBits_N[149] ;
 wire \ConfigBits_N[14] ;
 wire \ConfigBits_N[150] ;
 wire \ConfigBits_N[151] ;
 wire \ConfigBits_N[152] ;
 wire \ConfigBits_N[153] ;
 wire \ConfigBits_N[154] ;
 wire \ConfigBits_N[155] ;
 wire \ConfigBits_N[156] ;
 wire \ConfigBits_N[157] ;
 wire \ConfigBits_N[158] ;
 wire \ConfigBits_N[159] ;
 wire \ConfigBits_N[15] ;
 wire \ConfigBits_N[160] ;
 wire \ConfigBits_N[161] ;
 wire \ConfigBits_N[162] ;
 wire \ConfigBits_N[163] ;
 wire \ConfigBits_N[164] ;
 wire \ConfigBits_N[165] ;
 wire \ConfigBits_N[166] ;
 wire \ConfigBits_N[167] ;
 wire \ConfigBits_N[168] ;
 wire \ConfigBits_N[169] ;
 wire \ConfigBits_N[16] ;
 wire \ConfigBits_N[170] ;
 wire \ConfigBits_N[171] ;
 wire \ConfigBits_N[172] ;
 wire \ConfigBits_N[173] ;
 wire \ConfigBits_N[174] ;
 wire \ConfigBits_N[175] ;
 wire \ConfigBits_N[176] ;
 wire \ConfigBits_N[177] ;
 wire \ConfigBits_N[178] ;
 wire \ConfigBits_N[179] ;
 wire \ConfigBits_N[17] ;
 wire \ConfigBits_N[180] ;
 wire \ConfigBits_N[181] ;
 wire \ConfigBits_N[182] ;
 wire \ConfigBits_N[183] ;
 wire \ConfigBits_N[184] ;
 wire \ConfigBits_N[185] ;
 wire \ConfigBits_N[186] ;
 wire \ConfigBits_N[187] ;
 wire \ConfigBits_N[188] ;
 wire \ConfigBits_N[189] ;
 wire \ConfigBits_N[18] ;
 wire \ConfigBits_N[190] ;
 wire \ConfigBits_N[191] ;
 wire \ConfigBits_N[192] ;
 wire \ConfigBits_N[193] ;
 wire \ConfigBits_N[194] ;
 wire \ConfigBits_N[195] ;
 wire \ConfigBits_N[196] ;
 wire \ConfigBits_N[197] ;
 wire \ConfigBits_N[198] ;
 wire \ConfigBits_N[199] ;
 wire \ConfigBits_N[19] ;
 wire \ConfigBits_N[1] ;
 wire \ConfigBits_N[200] ;
 wire \ConfigBits_N[201] ;
 wire \ConfigBits_N[202] ;
 wire \ConfigBits_N[203] ;
 wire \ConfigBits_N[204] ;
 wire \ConfigBits_N[205] ;
 wire \ConfigBits_N[206] ;
 wire \ConfigBits_N[207] ;
 wire \ConfigBits_N[208] ;
 wire \ConfigBits_N[209] ;
 wire \ConfigBits_N[20] ;
 wire \ConfigBits_N[210] ;
 wire \ConfigBits_N[211] ;
 wire \ConfigBits_N[212] ;
 wire \ConfigBits_N[213] ;
 wire \ConfigBits_N[214] ;
 wire \ConfigBits_N[215] ;
 wire \ConfigBits_N[216] ;
 wire \ConfigBits_N[217] ;
 wire \ConfigBits_N[218] ;
 wire \ConfigBits_N[219] ;
 wire \ConfigBits_N[21] ;
 wire \ConfigBits_N[220] ;
 wire \ConfigBits_N[221] ;
 wire \ConfigBits_N[222] ;
 wire \ConfigBits_N[223] ;
 wire \ConfigBits_N[224] ;
 wire \ConfigBits_N[225] ;
 wire \ConfigBits_N[226] ;
 wire \ConfigBits_N[227] ;
 wire \ConfigBits_N[228] ;
 wire \ConfigBits_N[229] ;
 wire \ConfigBits_N[22] ;
 wire \ConfigBits_N[230] ;
 wire \ConfigBits_N[231] ;
 wire \ConfigBits_N[232] ;
 wire \ConfigBits_N[233] ;
 wire \ConfigBits_N[234] ;
 wire \ConfigBits_N[235] ;
 wire \ConfigBits_N[236] ;
 wire \ConfigBits_N[237] ;
 wire \ConfigBits_N[238] ;
 wire \ConfigBits_N[239] ;
 wire \ConfigBits_N[23] ;
 wire \ConfigBits_N[240] ;
 wire \ConfigBits_N[241] ;
 wire \ConfigBits_N[242] ;
 wire \ConfigBits_N[243] ;
 wire \ConfigBits_N[244] ;
 wire \ConfigBits_N[245] ;
 wire \ConfigBits_N[246] ;
 wire \ConfigBits_N[247] ;
 wire \ConfigBits_N[248] ;
 wire \ConfigBits_N[249] ;
 wire \ConfigBits_N[24] ;
 wire \ConfigBits_N[250] ;
 wire \ConfigBits_N[251] ;
 wire \ConfigBits_N[252] ;
 wire \ConfigBits_N[253] ;
 wire \ConfigBits_N[254] ;
 wire \ConfigBits_N[255] ;
 wire \ConfigBits_N[256] ;
 wire \ConfigBits_N[257] ;
 wire \ConfigBits_N[258] ;
 wire \ConfigBits_N[259] ;
 wire \ConfigBits_N[25] ;
 wire \ConfigBits_N[260] ;
 wire \ConfigBits_N[261] ;
 wire \ConfigBits_N[262] ;
 wire \ConfigBits_N[263] ;
 wire \ConfigBits_N[264] ;
 wire \ConfigBits_N[265] ;
 wire \ConfigBits_N[266] ;
 wire \ConfigBits_N[267] ;
 wire \ConfigBits_N[268] ;
 wire \ConfigBits_N[269] ;
 wire \ConfigBits_N[26] ;
 wire \ConfigBits_N[270] ;
 wire \ConfigBits_N[271] ;
 wire \ConfigBits_N[272] ;
 wire \ConfigBits_N[273] ;
 wire \ConfigBits_N[274] ;
 wire \ConfigBits_N[275] ;
 wire \ConfigBits_N[276] ;
 wire \ConfigBits_N[277] ;
 wire \ConfigBits_N[278] ;
 wire \ConfigBits_N[279] ;
 wire \ConfigBits_N[27] ;
 wire \ConfigBits_N[280] ;
 wire \ConfigBits_N[281] ;
 wire \ConfigBits_N[282] ;
 wire \ConfigBits_N[283] ;
 wire \ConfigBits_N[284] ;
 wire \ConfigBits_N[285] ;
 wire \ConfigBits_N[286] ;
 wire \ConfigBits_N[287] ;
 wire \ConfigBits_N[288] ;
 wire \ConfigBits_N[289] ;
 wire \ConfigBits_N[28] ;
 wire \ConfigBits_N[290] ;
 wire \ConfigBits_N[291] ;
 wire \ConfigBits_N[292] ;
 wire \ConfigBits_N[293] ;
 wire \ConfigBits_N[294] ;
 wire \ConfigBits_N[295] ;
 wire \ConfigBits_N[296] ;
 wire \ConfigBits_N[297] ;
 wire \ConfigBits_N[298] ;
 wire \ConfigBits_N[299] ;
 wire \ConfigBits_N[29] ;
 wire \ConfigBits_N[2] ;
 wire \ConfigBits_N[300] ;
 wire \ConfigBits_N[301] ;
 wire \ConfigBits_N[302] ;
 wire \ConfigBits_N[303] ;
 wire \ConfigBits_N[304] ;
 wire \ConfigBits_N[305] ;
 wire \ConfigBits_N[306] ;
 wire \ConfigBits_N[307] ;
 wire \ConfigBits_N[308] ;
 wire \ConfigBits_N[309] ;
 wire \ConfigBits_N[30] ;
 wire \ConfigBits_N[310] ;
 wire \ConfigBits_N[311] ;
 wire \ConfigBits_N[312] ;
 wire \ConfigBits_N[313] ;
 wire \ConfigBits_N[314] ;
 wire \ConfigBits_N[315] ;
 wire \ConfigBits_N[316] ;
 wire \ConfigBits_N[317] ;
 wire \ConfigBits_N[318] ;
 wire \ConfigBits_N[319] ;
 wire \ConfigBits_N[31] ;
 wire \ConfigBits_N[320] ;
 wire \ConfigBits_N[321] ;
 wire \ConfigBits_N[322] ;
 wire \ConfigBits_N[323] ;
 wire \ConfigBits_N[324] ;
 wire \ConfigBits_N[325] ;
 wire \ConfigBits_N[326] ;
 wire \ConfigBits_N[327] ;
 wire \ConfigBits_N[328] ;
 wire \ConfigBits_N[329] ;
 wire \ConfigBits_N[32] ;
 wire \ConfigBits_N[330] ;
 wire \ConfigBits_N[331] ;
 wire \ConfigBits_N[332] ;
 wire \ConfigBits_N[333] ;
 wire \ConfigBits_N[334] ;
 wire \ConfigBits_N[335] ;
 wire \ConfigBits_N[336] ;
 wire \ConfigBits_N[337] ;
 wire \ConfigBits_N[338] ;
 wire \ConfigBits_N[339] ;
 wire \ConfigBits_N[33] ;
 wire \ConfigBits_N[340] ;
 wire \ConfigBits_N[341] ;
 wire \ConfigBits_N[342] ;
 wire \ConfigBits_N[343] ;
 wire \ConfigBits_N[344] ;
 wire \ConfigBits_N[345] ;
 wire \ConfigBits_N[346] ;
 wire \ConfigBits_N[347] ;
 wire \ConfigBits_N[348] ;
 wire \ConfigBits_N[349] ;
 wire \ConfigBits_N[34] ;
 wire \ConfigBits_N[350] ;
 wire \ConfigBits_N[351] ;
 wire \ConfigBits_N[352] ;
 wire \ConfigBits_N[353] ;
 wire \ConfigBits_N[354] ;
 wire \ConfigBits_N[355] ;
 wire \ConfigBits_N[356] ;
 wire \ConfigBits_N[357] ;
 wire \ConfigBits_N[358] ;
 wire \ConfigBits_N[359] ;
 wire \ConfigBits_N[35] ;
 wire \ConfigBits_N[360] ;
 wire \ConfigBits_N[361] ;
 wire \ConfigBits_N[362] ;
 wire \ConfigBits_N[363] ;
 wire \ConfigBits_N[364] ;
 wire \ConfigBits_N[365] ;
 wire \ConfigBits_N[366] ;
 wire \ConfigBits_N[367] ;
 wire \ConfigBits_N[368] ;
 wire \ConfigBits_N[369] ;
 wire \ConfigBits_N[36] ;
 wire \ConfigBits_N[370] ;
 wire \ConfigBits_N[371] ;
 wire \ConfigBits_N[372] ;
 wire \ConfigBits_N[373] ;
 wire \ConfigBits_N[374] ;
 wire \ConfigBits_N[375] ;
 wire \ConfigBits_N[376] ;
 wire \ConfigBits_N[377] ;
 wire \ConfigBits_N[378] ;
 wire \ConfigBits_N[379] ;
 wire \ConfigBits_N[37] ;
 wire \ConfigBits_N[380] ;
 wire \ConfigBits_N[381] ;
 wire \ConfigBits_N[382] ;
 wire \ConfigBits_N[383] ;
 wire \ConfigBits_N[384] ;
 wire \ConfigBits_N[385] ;
 wire \ConfigBits_N[386] ;
 wire \ConfigBits_N[387] ;
 wire \ConfigBits_N[388] ;
 wire \ConfigBits_N[389] ;
 wire \ConfigBits_N[38] ;
 wire \ConfigBits_N[390] ;
 wire \ConfigBits_N[391] ;
 wire \ConfigBits_N[392] ;
 wire \ConfigBits_N[393] ;
 wire \ConfigBits_N[394] ;
 wire \ConfigBits_N[395] ;
 wire \ConfigBits_N[396] ;
 wire \ConfigBits_N[397] ;
 wire \ConfigBits_N[398] ;
 wire \ConfigBits_N[399] ;
 wire \ConfigBits_N[39] ;
 wire \ConfigBits_N[3] ;
 wire \ConfigBits_N[400] ;
 wire \ConfigBits_N[401] ;
 wire \ConfigBits_N[402] ;
 wire \ConfigBits_N[403] ;
 wire \ConfigBits_N[404] ;
 wire \ConfigBits_N[405] ;
 wire \ConfigBits_N[406] ;
 wire \ConfigBits_N[407] ;
 wire \ConfigBits_N[408] ;
 wire \ConfigBits_N[409] ;
 wire \ConfigBits_N[40] ;
 wire \ConfigBits_N[410] ;
 wire \ConfigBits_N[411] ;
 wire \ConfigBits_N[412] ;
 wire \ConfigBits_N[413] ;
 wire \ConfigBits_N[414] ;
 wire \ConfigBits_N[415] ;
 wire \ConfigBits_N[416] ;
 wire \ConfigBits_N[417] ;
 wire \ConfigBits_N[418] ;
 wire \ConfigBits_N[419] ;
 wire \ConfigBits_N[41] ;
 wire \ConfigBits_N[420] ;
 wire \ConfigBits_N[421] ;
 wire \ConfigBits_N[422] ;
 wire \ConfigBits_N[423] ;
 wire \ConfigBits_N[424] ;
 wire \ConfigBits_N[425] ;
 wire \ConfigBits_N[426] ;
 wire \ConfigBits_N[427] ;
 wire \ConfigBits_N[428] ;
 wire \ConfigBits_N[429] ;
 wire \ConfigBits_N[42] ;
 wire \ConfigBits_N[430] ;
 wire \ConfigBits_N[431] ;
 wire \ConfigBits_N[432] ;
 wire \ConfigBits_N[433] ;
 wire \ConfigBits_N[434] ;
 wire \ConfigBits_N[435] ;
 wire \ConfigBits_N[436] ;
 wire \ConfigBits_N[437] ;
 wire \ConfigBits_N[438] ;
 wire \ConfigBits_N[439] ;
 wire \ConfigBits_N[43] ;
 wire \ConfigBits_N[440] ;
 wire \ConfigBits_N[441] ;
 wire \ConfigBits_N[442] ;
 wire \ConfigBits_N[443] ;
 wire \ConfigBits_N[444] ;
 wire \ConfigBits_N[445] ;
 wire \ConfigBits_N[446] ;
 wire \ConfigBits_N[447] ;
 wire \ConfigBits_N[448] ;
 wire \ConfigBits_N[449] ;
 wire \ConfigBits_N[44] ;
 wire \ConfigBits_N[450] ;
 wire \ConfigBits_N[451] ;
 wire \ConfigBits_N[452] ;
 wire \ConfigBits_N[453] ;
 wire \ConfigBits_N[454] ;
 wire \ConfigBits_N[455] ;
 wire \ConfigBits_N[456] ;
 wire \ConfigBits_N[457] ;
 wire \ConfigBits_N[458] ;
 wire \ConfigBits_N[459] ;
 wire \ConfigBits_N[45] ;
 wire \ConfigBits_N[460] ;
 wire \ConfigBits_N[461] ;
 wire \ConfigBits_N[462] ;
 wire \ConfigBits_N[463] ;
 wire \ConfigBits_N[464] ;
 wire \ConfigBits_N[465] ;
 wire \ConfigBits_N[466] ;
 wire \ConfigBits_N[467] ;
 wire \ConfigBits_N[468] ;
 wire \ConfigBits_N[469] ;
 wire \ConfigBits_N[46] ;
 wire \ConfigBits_N[470] ;
 wire \ConfigBits_N[471] ;
 wire \ConfigBits_N[472] ;
 wire \ConfigBits_N[473] ;
 wire \ConfigBits_N[474] ;
 wire \ConfigBits_N[475] ;
 wire \ConfigBits_N[476] ;
 wire \ConfigBits_N[477] ;
 wire \ConfigBits_N[478] ;
 wire \ConfigBits_N[479] ;
 wire \ConfigBits_N[47] ;
 wire \ConfigBits_N[480] ;
 wire \ConfigBits_N[481] ;
 wire \ConfigBits_N[482] ;
 wire \ConfigBits_N[483] ;
 wire \ConfigBits_N[484] ;
 wire \ConfigBits_N[485] ;
 wire \ConfigBits_N[486] ;
 wire \ConfigBits_N[487] ;
 wire \ConfigBits_N[488] ;
 wire \ConfigBits_N[489] ;
 wire \ConfigBits_N[48] ;
 wire \ConfigBits_N[490] ;
 wire \ConfigBits_N[491] ;
 wire \ConfigBits_N[492] ;
 wire \ConfigBits_N[493] ;
 wire \ConfigBits_N[494] ;
 wire \ConfigBits_N[495] ;
 wire \ConfigBits_N[496] ;
 wire \ConfigBits_N[497] ;
 wire \ConfigBits_N[498] ;
 wire \ConfigBits_N[499] ;
 wire \ConfigBits_N[49] ;
 wire \ConfigBits_N[4] ;
 wire \ConfigBits_N[500] ;
 wire \ConfigBits_N[501] ;
 wire \ConfigBits_N[502] ;
 wire \ConfigBits_N[503] ;
 wire \ConfigBits_N[504] ;
 wire \ConfigBits_N[505] ;
 wire \ConfigBits_N[506] ;
 wire \ConfigBits_N[507] ;
 wire \ConfigBits_N[508] ;
 wire \ConfigBits_N[509] ;
 wire \ConfigBits_N[50] ;
 wire \ConfigBits_N[510] ;
 wire \ConfigBits_N[511] ;
 wire \ConfigBits_N[512] ;
 wire \ConfigBits_N[513] ;
 wire \ConfigBits_N[514] ;
 wire \ConfigBits_N[515] ;
 wire \ConfigBits_N[516] ;
 wire \ConfigBits_N[517] ;
 wire \ConfigBits_N[518] ;
 wire \ConfigBits_N[519] ;
 wire \ConfigBits_N[51] ;
 wire \ConfigBits_N[520] ;
 wire \ConfigBits_N[521] ;
 wire \ConfigBits_N[522] ;
 wire \ConfigBits_N[523] ;
 wire \ConfigBits_N[524] ;
 wire \ConfigBits_N[525] ;
 wire \ConfigBits_N[526] ;
 wire \ConfigBits_N[527] ;
 wire \ConfigBits_N[528] ;
 wire \ConfigBits_N[529] ;
 wire \ConfigBits_N[52] ;
 wire \ConfigBits_N[530] ;
 wire \ConfigBits_N[531] ;
 wire \ConfigBits_N[532] ;
 wire \ConfigBits_N[533] ;
 wire \ConfigBits_N[534] ;
 wire \ConfigBits_N[535] ;
 wire \ConfigBits_N[536] ;
 wire \ConfigBits_N[537] ;
 wire \ConfigBits_N[538] ;
 wire \ConfigBits_N[539] ;
 wire \ConfigBits_N[53] ;
 wire \ConfigBits_N[540] ;
 wire \ConfigBits_N[541] ;
 wire \ConfigBits_N[542] ;
 wire \ConfigBits_N[543] ;
 wire \ConfigBits_N[544] ;
 wire \ConfigBits_N[545] ;
 wire \ConfigBits_N[546] ;
 wire \ConfigBits_N[547] ;
 wire \ConfigBits_N[548] ;
 wire \ConfigBits_N[549] ;
 wire \ConfigBits_N[54] ;
 wire \ConfigBits_N[550] ;
 wire \ConfigBits_N[551] ;
 wire \ConfigBits_N[552] ;
 wire \ConfigBits_N[553] ;
 wire \ConfigBits_N[554] ;
 wire \ConfigBits_N[555] ;
 wire \ConfigBits_N[556] ;
 wire \ConfigBits_N[557] ;
 wire \ConfigBits_N[558] ;
 wire \ConfigBits_N[559] ;
 wire \ConfigBits_N[55] ;
 wire \ConfigBits_N[560] ;
 wire \ConfigBits_N[561] ;
 wire \ConfigBits_N[562] ;
 wire \ConfigBits_N[563] ;
 wire \ConfigBits_N[564] ;
 wire \ConfigBits_N[565] ;
 wire \ConfigBits_N[566] ;
 wire \ConfigBits_N[567] ;
 wire \ConfigBits_N[568] ;
 wire \ConfigBits_N[569] ;
 wire \ConfigBits_N[56] ;
 wire \ConfigBits_N[570] ;
 wire \ConfigBits_N[571] ;
 wire \ConfigBits_N[572] ;
 wire \ConfigBits_N[573] ;
 wire \ConfigBits_N[574] ;
 wire \ConfigBits_N[575] ;
 wire \ConfigBits_N[576] ;
 wire \ConfigBits_N[577] ;
 wire \ConfigBits_N[578] ;
 wire \ConfigBits_N[579] ;
 wire \ConfigBits_N[57] ;
 wire \ConfigBits_N[580] ;
 wire \ConfigBits_N[581] ;
 wire \ConfigBits_N[582] ;
 wire \ConfigBits_N[583] ;
 wire \ConfigBits_N[584] ;
 wire \ConfigBits_N[585] ;
 wire \ConfigBits_N[586] ;
 wire \ConfigBits_N[587] ;
 wire \ConfigBits_N[588] ;
 wire \ConfigBits_N[589] ;
 wire \ConfigBits_N[58] ;
 wire \ConfigBits_N[590] ;
 wire \ConfigBits_N[591] ;
 wire \ConfigBits_N[592] ;
 wire \ConfigBits_N[593] ;
 wire \ConfigBits_N[594] ;
 wire \ConfigBits_N[595] ;
 wire \ConfigBits_N[596] ;
 wire \ConfigBits_N[597] ;
 wire \ConfigBits_N[598] ;
 wire \ConfigBits_N[599] ;
 wire \ConfigBits_N[59] ;
 wire \ConfigBits_N[5] ;
 wire \ConfigBits_N[600] ;
 wire \ConfigBits_N[601] ;
 wire \ConfigBits_N[602] ;
 wire \ConfigBits_N[603] ;
 wire \ConfigBits_N[604] ;
 wire \ConfigBits_N[605] ;
 wire \ConfigBits_N[606] ;
 wire \ConfigBits_N[607] ;
 wire \ConfigBits_N[608] ;
 wire \ConfigBits_N[609] ;
 wire \ConfigBits_N[60] ;
 wire \ConfigBits_N[610] ;
 wire \ConfigBits_N[611] ;
 wire \ConfigBits_N[612] ;
 wire \ConfigBits_N[613] ;
 wire \ConfigBits_N[614] ;
 wire \ConfigBits_N[615] ;
 wire \ConfigBits_N[61] ;
 wire \ConfigBits_N[62] ;
 wire \ConfigBits_N[63] ;
 wire \ConfigBits_N[64] ;
 wire \ConfigBits_N[65] ;
 wire \ConfigBits_N[66] ;
 wire \ConfigBits_N[67] ;
 wire \ConfigBits_N[68] ;
 wire \ConfigBits_N[69] ;
 wire \ConfigBits_N[6] ;
 wire \ConfigBits_N[70] ;
 wire \ConfigBits_N[71] ;
 wire \ConfigBits_N[72] ;
 wire \ConfigBits_N[73] ;
 wire \ConfigBits_N[74] ;
 wire \ConfigBits_N[75] ;
 wire \ConfigBits_N[76] ;
 wire \ConfigBits_N[77] ;
 wire \ConfigBits_N[78] ;
 wire \ConfigBits_N[79] ;
 wire \ConfigBits_N[7] ;
 wire \ConfigBits_N[80] ;
 wire \ConfigBits_N[81] ;
 wire \ConfigBits_N[82] ;
 wire \ConfigBits_N[83] ;
 wire \ConfigBits_N[84] ;
 wire \ConfigBits_N[85] ;
 wire \ConfigBits_N[86] ;
 wire \ConfigBits_N[87] ;
 wire \ConfigBits_N[88] ;
 wire \ConfigBits_N[89] ;
 wire \ConfigBits_N[8] ;
 wire \ConfigBits_N[90] ;
 wire \ConfigBits_N[91] ;
 wire \ConfigBits_N[92] ;
 wire \ConfigBits_N[93] ;
 wire \ConfigBits_N[94] ;
 wire \ConfigBits_N[95] ;
 wire \ConfigBits_N[96] ;
 wire \ConfigBits_N[97] ;
 wire \ConfigBits_N[98] ;
 wire \ConfigBits_N[99] ;
 wire \ConfigBits_N[9] ;
 wire D;
 wire E;
 wire \E6BEG_i[0] ;
 wire \E6BEG_i[1] ;
 wire \E6BEG_i[2] ;
 wire \E6BEG_i[3] ;
 wire \E6BEG_i[4] ;
 wire \E6BEG_i[5] ;
 wire \E6BEG_i[6] ;
 wire \E6BEG_i[7] ;
 wire \E6BEG_i[8] ;
 wire \E6BEG_i[9] ;
 wire \EE4BEG_i[0] ;
 wire \EE4BEG_i[10] ;
 wire \EE4BEG_i[11] ;
 wire \EE4BEG_i[1] ;
 wire \EE4BEG_i[2] ;
 wire \EE4BEG_i[3] ;
 wire \EE4BEG_i[4] ;
 wire \EE4BEG_i[5] ;
 wire \EE4BEG_i[6] ;
 wire \EE4BEG_i[7] ;
 wire \EE4BEG_i[8] ;
 wire \EE4BEG_i[9] ;
 wire F;
 wire \FrameData_O_i[0] ;
 wire \FrameData_O_i[10] ;
 wire \FrameData_O_i[11] ;
 wire \FrameData_O_i[12] ;
 wire \FrameData_O_i[13] ;
 wire \FrameData_O_i[14] ;
 wire \FrameData_O_i[15] ;
 wire \FrameData_O_i[16] ;
 wire \FrameData_O_i[17] ;
 wire \FrameData_O_i[18] ;
 wire \FrameData_O_i[19] ;
 wire \FrameData_O_i[1] ;
 wire \FrameData_O_i[20] ;
 wire \FrameData_O_i[21] ;
 wire \FrameData_O_i[22] ;
 wire \FrameData_O_i[23] ;
 wire \FrameData_O_i[24] ;
 wire \FrameData_O_i[25] ;
 wire \FrameData_O_i[26] ;
 wire \FrameData_O_i[27] ;
 wire \FrameData_O_i[28] ;
 wire \FrameData_O_i[29] ;
 wire \FrameData_O_i[2] ;
 wire \FrameData_O_i[30] ;
 wire \FrameData_O_i[31] ;
 wire \FrameData_O_i[3] ;
 wire \FrameData_O_i[4] ;
 wire \FrameData_O_i[5] ;
 wire \FrameData_O_i[6] ;
 wire \FrameData_O_i[7] ;
 wire \FrameData_O_i[8] ;
 wire \FrameData_O_i[9] ;
 wire \FrameStrobe_O_i[0] ;
 wire \FrameStrobe_O_i[10] ;
 wire \FrameStrobe_O_i[11] ;
 wire \FrameStrobe_O_i[12] ;
 wire \FrameStrobe_O_i[13] ;
 wire \FrameStrobe_O_i[14] ;
 wire \FrameStrobe_O_i[15] ;
 wire \FrameStrobe_O_i[16] ;
 wire \FrameStrobe_O_i[17] ;
 wire \FrameStrobe_O_i[18] ;
 wire \FrameStrobe_O_i[19] ;
 wire \FrameStrobe_O_i[1] ;
 wire \FrameStrobe_O_i[2] ;
 wire \FrameStrobe_O_i[3] ;
 wire \FrameStrobe_O_i[4] ;
 wire \FrameStrobe_O_i[5] ;
 wire \FrameStrobe_O_i[6] ;
 wire \FrameStrobe_O_i[7] ;
 wire \FrameStrobe_O_i[8] ;
 wire \FrameStrobe_O_i[9] ;
 wire G;
 wire H;
 wire \Inst_LA_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/I0mux ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/LUT_flop ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/LUT_out ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_00_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_01_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_02_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_03_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_04_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_05_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/_06_ ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ;
 wire \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_MUX8LUT_frame_config_mux/AD ;
 wire \Inst_MUX8LUT_frame_config_mux/AH ;
 wire \Inst_MUX8LUT_frame_config_mux/CD ;
 wire \Inst_MUX8LUT_frame_config_mux/EH ;
 wire \Inst_MUX8LUT_frame_config_mux/EH_GH ;
 wire \Inst_MUX8LUT_frame_config_mux/GH ;
 wire \Inst_MUX8LUT_frame_config_mux/sCD ;
 wire \Inst_MUX8LUT_frame_config_mux/sEF ;
 wire \Inst_MUX8LUT_frame_config_mux/sEH ;
 wire \Inst_MUX8LUT_frame_config_mux/sGH ;
 wire \J2END_AB_BEG[0] ;
 wire \J2END_AB_BEG[1] ;
 wire \J2END_AB_BEG[2] ;
 wire \J2END_AB_BEG[3] ;
 wire \J2END_CD_BEG[0] ;
 wire \J2END_CD_BEG[1] ;
 wire \J2END_CD_BEG[2] ;
 wire \J2END_CD_BEG[3] ;
 wire \J2END_EF_BEG[0] ;
 wire \J2END_EF_BEG[1] ;
 wire \J2END_EF_BEG[2] ;
 wire \J2END_EF_BEG[3] ;
 wire \J2END_GH_BEG[0] ;
 wire \J2END_GH_BEG[1] ;
 wire \J2END_GH_BEG[2] ;
 wire \J2END_GH_BEG[3] ;
 wire \J2MID_ABa_BEG[0] ;
 wire \J2MID_ABa_BEG[1] ;
 wire \J2MID_ABa_BEG[2] ;
 wire \J2MID_ABa_BEG[3] ;
 wire \J2MID_ABb_BEG[0] ;
 wire \J2MID_ABb_BEG[1] ;
 wire \J2MID_ABb_BEG[2] ;
 wire \J2MID_ABb_BEG[3] ;
 wire \J2MID_CDa_BEG[0] ;
 wire \J2MID_CDa_BEG[1] ;
 wire \J2MID_CDa_BEG[2] ;
 wire \J2MID_CDa_BEG[3] ;
 wire \J2MID_CDb_BEG[0] ;
 wire \J2MID_CDb_BEG[1] ;
 wire \J2MID_CDb_BEG[2] ;
 wire \J2MID_CDb_BEG[3] ;
 wire \J2MID_EFa_BEG[0] ;
 wire \J2MID_EFa_BEG[1] ;
 wire \J2MID_EFa_BEG[2] ;
 wire \J2MID_EFa_BEG[3] ;
 wire \J2MID_EFb_BEG[0] ;
 wire \J2MID_EFb_BEG[1] ;
 wire \J2MID_EFb_BEG[2] ;
 wire \J2MID_EFb_BEG[3] ;
 wire \J2MID_GHa_BEG[0] ;
 wire \J2MID_GHa_BEG[1] ;
 wire \J2MID_GHa_BEG[2] ;
 wire \J2MID_GHa_BEG[3] ;
 wire \J2MID_GHb_BEG[0] ;
 wire \J2MID_GHb_BEG[1] ;
 wire \J2MID_GHb_BEG[2] ;
 wire \J2MID_GHb_BEG[3] ;
 wire \JE2BEG[0] ;
 wire \JE2BEG[1] ;
 wire \JE2BEG[2] ;
 wire \JE2BEG[3] ;
 wire \JE2BEG[4] ;
 wire \JE2BEG[5] ;
 wire \JE2BEG[6] ;
 wire \JE2BEG[7] ;
 wire \JN2BEG[0] ;
 wire \JN2BEG[1] ;
 wire \JN2BEG[2] ;
 wire \JN2BEG[3] ;
 wire \JN2BEG[4] ;
 wire \JN2BEG[5] ;
 wire \JN2BEG[6] ;
 wire \JN2BEG[7] ;
 wire \JS2BEG[0] ;
 wire \JS2BEG[1] ;
 wire \JS2BEG[2] ;
 wire \JS2BEG[3] ;
 wire \JS2BEG[4] ;
 wire \JS2BEG[5] ;
 wire \JS2BEG[6] ;
 wire \JS2BEG[7] ;
 wire \JW2BEG[0] ;
 wire \JW2BEG[1] ;
 wire \JW2BEG[2] ;
 wire \JW2BEG[3] ;
 wire \JW2BEG[4] ;
 wire \JW2BEG[5] ;
 wire \JW2BEG[6] ;
 wire \JW2BEG[7] ;
 wire J_EN_BEG;
 wire J_SR_BEG;
 wire \J_l_AB_BEG[0] ;
 wire \J_l_AB_BEG[1] ;
 wire \J_l_AB_BEG[2] ;
 wire \J_l_AB_BEG[3] ;
 wire \J_l_CD_BEG[0] ;
 wire \J_l_CD_BEG[1] ;
 wire \J_l_CD_BEG[2] ;
 wire \J_l_CD_BEG[3] ;
 wire \J_l_EF_BEG[0] ;
 wire \J_l_EF_BEG[1] ;
 wire \J_l_EF_BEG[2] ;
 wire \J_l_EF_BEG[3] ;
 wire \J_l_GH_BEG[0] ;
 wire \J_l_GH_BEG[1] ;
 wire \J_l_GH_BEG[2] ;
 wire \J_l_GH_BEG[3] ;
 wire LA_Ci;
 wire LA_Co;
 wire LA_EN;
 wire LA_I0;
 wire LA_I1;
 wire LA_I2;
 wire LA_I3;
 wire LA_O;
 wire LA_SR;
 wire LB_Ci;
 wire LB_Co;
 wire LB_EN;
 wire LB_I0;
 wire LB_I1;
 wire LB_I2;
 wire LB_I3;
 wire LB_O;
 wire LB_SR;
 wire LC_Ci;
 wire LC_Co;
 wire LC_EN;
 wire LC_I0;
 wire LC_I1;
 wire LC_I2;
 wire LC_I3;
 wire LC_O;
 wire LC_SR;
 wire LD_Ci;
 wire LD_Co;
 wire LD_EN;
 wire LD_I0;
 wire LD_I1;
 wire LD_I2;
 wire LD_I3;
 wire LD_O;
 wire LD_SR;
 wire LE_Ci;
 wire LE_Co;
 wire LE_EN;
 wire LE_I0;
 wire LE_I1;
 wire LE_I2;
 wire LE_I3;
 wire LE_O;
 wire LE_SR;
 wire LF_Ci;
 wire LF_Co;
 wire LF_EN;
 wire LF_I0;
 wire LF_I1;
 wire LF_I2;
 wire LF_I3;
 wire LF_O;
 wire LF_SR;
 wire LG_Ci;
 wire LG_Co;
 wire LG_EN;
 wire LG_I0;
 wire LG_I1;
 wire LG_I2;
 wire LG_I3;
 wire LG_O;
 wire LG_SR;
 wire LH_Ci;
 wire LH_Co;
 wire LH_EN;
 wire LH_I0;
 wire LH_I1;
 wire LH_I2;
 wire LH_I3;
 wire LH_O;
 wire LH_SR;
 wire M_AB;
 wire M_AD;
 wire M_AH;
 wire M_EF;
 wire \N4BEG_i[0] ;
 wire \N4BEG_i[10] ;
 wire \N4BEG_i[11] ;
 wire \N4BEG_i[1] ;
 wire \N4BEG_i[2] ;
 wire \N4BEG_i[3] ;
 wire \N4BEG_i[4] ;
 wire \N4BEG_i[5] ;
 wire \N4BEG_i[6] ;
 wire \N4BEG_i[7] ;
 wire \N4BEG_i[8] ;
 wire \N4BEG_i[9] ;
 wire \NN4BEG_i[0] ;
 wire \NN4BEG_i[10] ;
 wire \NN4BEG_i[11] ;
 wire \NN4BEG_i[1] ;
 wire \NN4BEG_i[2] ;
 wire \NN4BEG_i[3] ;
 wire \NN4BEG_i[4] ;
 wire \NN4BEG_i[5] ;
 wire \NN4BEG_i[6] ;
 wire \NN4BEG_i[7] ;
 wire \NN4BEG_i[8] ;
 wire \NN4BEG_i[9] ;
 wire S0;
 wire S1;
 wire S2;
 wire S3;
 wire \S4BEG_i[0] ;
 wire \S4BEG_i[10] ;
 wire \S4BEG_i[11] ;
 wire \S4BEG_i[1] ;
 wire \S4BEG_i[2] ;
 wire \S4BEG_i[3] ;
 wire \S4BEG_i[4] ;
 wire \S4BEG_i[5] ;
 wire \S4BEG_i[6] ;
 wire \S4BEG_i[7] ;
 wire \S4BEG_i[8] ;
 wire \S4BEG_i[9] ;
 wire \SS4BEG_i[0] ;
 wire \SS4BEG_i[10] ;
 wire \SS4BEG_i[11] ;
 wire \SS4BEG_i[1] ;
 wire \SS4BEG_i[2] ;
 wire \SS4BEG_i[3] ;
 wire \SS4BEG_i[4] ;
 wire \SS4BEG_i[5] ;
 wire \SS4BEG_i[6] ;
 wire \SS4BEG_i[7] ;
 wire \SS4BEG_i[8] ;
 wire \SS4BEG_i[9] ;
 wire \W6BEG_i[0] ;
 wire \W6BEG_i[1] ;
 wire \W6BEG_i[2] ;
 wire \W6BEG_i[3] ;
 wire \W6BEG_i[4] ;
 wire \W6BEG_i[5] ;
 wire \W6BEG_i[6] ;
 wire \W6BEG_i[7] ;
 wire \W6BEG_i[8] ;
 wire \W6BEG_i[9] ;
 wire \WW4BEG_i[0] ;
 wire \WW4BEG_i[10] ;
 wire \WW4BEG_i[11] ;
 wire \WW4BEG_i[1] ;
 wire \WW4BEG_i[2] ;
 wire \WW4BEG_i[3] ;
 wire \WW4BEG_i[4] ;
 wire \WW4BEG_i[5] ;
 wire \WW4BEG_i[6] ;
 wire \WW4BEG_i[7] ;
 wire \WW4BEG_i[8] ;
 wire \WW4BEG_i[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\JS2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\WW4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\WW4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\S4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\W6BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_0/_0__A  (.DIODE(\E6BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_1/_0__A  (.DIODE(\E6BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_2/_0__A  (.DIODE(\E6BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_3/_0__A  (.DIODE(\E6BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_4/_0__A  (.DIODE(\E6BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_5/_0__A  (.DIODE(\E6BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_6/_0__A  (.DIODE(\E6BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_7/_0__A  (.DIODE(\E6BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_8/_0__A  (.DIODE(\E6BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_E6BEG_outbuf_9/_0__A  (.DIODE(\E6BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_0/_0__A  (.DIODE(\EE4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_1/_0__A  (.DIODE(\EE4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_10/_0__A  (.DIODE(\EE4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_11/_0__A  (.DIODE(\EE4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_2/_0__A  (.DIODE(\EE4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_3/_0__A  (.DIODE(\EE4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_4/_0__A  (.DIODE(\EE4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_5/_0__A  (.DIODE(\EE4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_6/_0__A  (.DIODE(\EE4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_7/_0__A  (.DIODE(\EE4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_8/_0__A  (.DIODE(\EE4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_EE4BEG_outbuf_9/_0__A  (.DIODE(\EE4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LE_LUT4c_frame_config_dffesr/_10__A  (.DIODE(LE_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S1  (.DIODE(LE_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LF_LUT4c_frame_config_dffesr/_10__A  (.DIODE(LF_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S1  (.DIODE(LF_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/_09__A  (.DIODE(LG_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/_10__A  (.DIODE(LG_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/_11__A1  (.DIODE(LG_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/_12__A1  (.DIODE(LG_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S0  (.DIODE(LG_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S1  (.DIODE(LG_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/_09__A  (.DIODE(LH_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/_10__A  (.DIODE(LH_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/_11__A1  (.DIODE(LH_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/_12__A1  (.DIODE(LH_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S0  (.DIODE(LH_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4_S1  (.DIODE(LH_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit0_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit10_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit11_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit12_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit13_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit14_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit15_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit16_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit17_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit18_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit19_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit1_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit20_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit21_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit22_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit23_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit24_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit3_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit4_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit5_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit6_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit7_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit8_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame0_bit9_GATE  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit0_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit10_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit11_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit12_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit13_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit14_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit15_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit16_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit17_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit18_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit19_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit1_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit20_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit21_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit22_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit23_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit24_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit25_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit26_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit27_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit28_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit29_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit2_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit30_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit31_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit3_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit4_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit5_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit6_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit7_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit8_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame10_bit9_GATE  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit0_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit10_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit11_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit12_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit13_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit14_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit15_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit16_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit17_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit18_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit19_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit1_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit20_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit21_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit22_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit23_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit24_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit25_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit26_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit27_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit28_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit29_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit2_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit30_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit31_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit3_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit4_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit5_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit6_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit7_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit8_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame11_bit9_GATE  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit0_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit10_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit11_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit12_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit13_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit14_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit15_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit16_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit17_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit18_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit19_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit1_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit20_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit21_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit22_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit23_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit24_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit25_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit26_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit27_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit28_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit29_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit2_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit30_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit31_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit3_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit4_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit5_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit6_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit7_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit8_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame12_bit9_GATE  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit0_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit10_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit11_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit12_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit13_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit14_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit15_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit16_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit17_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit18_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit19_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit1_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit20_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit21_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit22_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit23_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit24_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit25_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit26_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit27_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit28_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit29_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit2_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit30_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit31_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit3_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit4_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit5_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit6_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit7_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit8_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame13_bit9_GATE  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit0_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit10_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit11_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit12_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit13_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit14_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit15_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit16_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit17_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit18_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit19_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit1_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit20_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit21_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit22_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit23_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit24_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit25_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit26_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit27_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit28_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit29_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit2_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit30_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit31_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit3_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit4_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit5_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit6_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit7_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit8_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame14_bit9_GATE  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit0_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit10_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit11_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit12_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit13_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit14_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit15_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit16_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit17_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit18_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit19_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit1_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit20_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit21_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit22_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit23_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit24_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit25_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit26_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit27_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit28_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit29_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit2_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit30_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit31_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit3_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit4_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit5_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit6_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit7_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit8_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame15_bit9_GATE  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit0_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit10_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit11_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit12_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit13_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit14_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit15_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit16_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit17_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit18_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit19_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit1_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit20_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit21_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit22_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit23_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit24_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit25_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit26_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit27_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit28_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit29_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit2_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit30_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit31_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit3_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit4_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit5_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit6_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit7_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit8_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame16_bit9_GATE  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit0_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit10_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit11_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit12_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit13_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit14_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit15_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit16_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit17_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit18_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit19_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit1_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit20_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit21_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit22_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit23_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit24_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit25_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit26_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit27_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit28_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit29_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit2_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit30_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit31_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit3_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit4_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit5_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit6_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit7_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit8_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame17_bit9_GATE  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit0_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit10_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit11_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit12_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit13_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit14_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit15_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit16_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit17_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit18_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit19_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit1_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit20_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit21_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit22_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit23_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit24_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit25_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit26_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit27_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit28_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit29_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit2_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit30_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit31_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit3_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit4_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit5_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit6_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit7_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit8_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame18_bit9_GATE  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit10_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit11_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit12_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit13_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit14_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit15_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit16_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit17_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit18_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit19_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit20_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit21_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit22_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit23_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit24_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit25_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit2_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit3_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit4_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit5_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit6_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit7_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit8_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame19_bit9_GATE  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit10_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit11_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit12_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit13_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit14_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit15_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit16_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit17_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit18_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit19_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit20_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit21_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit22_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit23_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit24_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit25_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit26_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit27_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit28_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit29_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit2_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit30_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit31_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit3_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit4_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit5_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit7_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit8_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame1_bit9_GATE  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit10_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit11_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit12_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit13_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit14_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit15_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit16_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit17_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit18_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit19_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit1_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit20_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit21_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit22_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit23_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit24_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit25_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit26_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit27_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit28_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit30_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit31_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit4_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit5_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit6_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit7_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit8_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame2_bit9_GATE  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit10_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit11_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit12_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit13_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit14_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit15_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit16_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit17_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit18_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit19_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit1_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit20_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit21_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit22_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit23_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit24_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit25_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit26_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit27_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit28_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit29_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit2_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit30_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit31_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit3_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit4_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit5_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit6_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit7_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit8_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame3_bit9_GATE  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit0_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit10_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit11_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit12_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit13_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit14_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit15_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit16_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit17_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit18_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit19_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit1_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit20_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit21_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit22_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit23_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit24_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit25_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit26_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit27_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit28_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit29_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit2_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit30_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit31_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit3_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit4_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit5_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit6_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit7_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit8_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame4_bit9_GATE  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit0_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit10_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit11_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit12_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit13_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit14_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit15_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit16_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit17_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit18_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit19_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit1_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit20_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit21_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit22_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit23_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit24_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit25_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit26_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit27_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit28_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit29_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit2_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit30_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit31_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit3_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit4_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit5_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit6_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit7_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit8_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame5_bit9_GATE  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit0_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit10_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit11_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit12_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit13_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit14_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit15_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit16_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit17_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit18_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit19_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit1_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit20_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit21_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit22_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit23_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit24_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit25_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit26_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit27_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit28_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit29_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit2_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit30_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit31_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit3_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit4_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit5_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit6_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit7_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit8_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame6_bit9_GATE  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit0_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit10_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit11_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit12_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit13_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit14_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit15_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit16_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit17_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit18_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit19_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit1_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit20_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit21_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit22_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit23_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit24_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit25_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit26_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit27_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit28_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit29_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit2_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit30_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit31_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit3_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit4_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit5_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit6_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit7_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit8_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame7_bit9_GATE  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit0_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit10_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit11_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit12_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit13_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit14_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit15_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit16_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit17_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit18_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit19_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit1_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit20_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit21_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit22_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit23_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit24_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit25_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit26_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit27_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit28_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit29_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit2_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit30_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit31_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit3_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit4_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit5_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit6_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit7_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit8_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame8_bit9_GATE  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit0_D  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit0_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit10_D  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit10_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit11_D  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit11_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit12_D  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit12_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit13_D  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit13_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit14_D  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit14_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit15_D  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit15_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit16_D  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit16_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit17_D  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit17_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit18_D  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit18_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit19_D  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit19_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit1_D  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit1_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit20_D  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit20_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit21_D  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit21_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit22_D  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit22_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit23_D  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit23_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit24_D  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit24_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit25_D  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit25_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit26_D  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit26_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit27_D  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit27_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit28_D  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit28_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit29_D  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit29_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit2_D  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit2_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit30_D  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit30_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit31_D  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit31_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit3_D  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit3_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit4_D  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit4_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit5_D  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit5_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit6_D  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit6_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit7_D  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit7_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit8_D  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit8_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit9_D  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_ConfigMem/Inst_Frame9_bit9_GATE  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_032__A  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_033__A  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_034__A  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_036__A  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_037__A  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_038__A  (.DIODE(\JE2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_039__A  (.DIODE(\JE2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_040__A  (.DIODE(\JE2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_041__A  (.DIODE(\JE2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_042__A  (.DIODE(\JE2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_043__A  (.DIODE(\JE2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_044__A  (.DIODE(\JE2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_045__A  (.DIODE(\JE2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_046__A  (.DIODE(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_047__A  (.DIODE(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_048__A  (.DIODE(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_049__A  (.DIODE(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_050__A  (.DIODE(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_051__A  (.DIODE(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_052__A  (.DIODE(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_053__A  (.DIODE(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_054__A  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_055__A  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_056__A  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_065__A  (.DIODE(\JN2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_066__A  (.DIODE(\JN2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_067__A  (.DIODE(\JN2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_068__A  (.DIODE(\JN2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_069__A  (.DIODE(\JN2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_071__A  (.DIODE(\JN2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_072__A  (.DIODE(\JN2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_073__A  (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_074__A  (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_075__A  (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_076__A  (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_077__A  (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_078__A  (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_079__A  (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_080__A  (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_081__A  (.DIODE(\JS2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_082__A  (.DIODE(\JS2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_083__A  (.DIODE(\JS2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_084__A  (.DIODE(\JS2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_085__A  (.DIODE(\JS2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_086__A  (.DIODE(\JS2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_087__A  (.DIODE(\JS2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_089__A  (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_090__A  (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_091__A  (.DIODE(net168),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_092__A  (.DIODE(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_093__A  (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_094__A  (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_095__A  (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_096__A  (.DIODE(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_098__A  (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_099__A  (.DIODE(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_100__A  (.DIODE(\JW2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_101__A  (.DIODE(\JW2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_102__A  (.DIODE(\JW2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_103__A  (.DIODE(\JW2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_104__A  (.DIODE(\JW2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_105__A  (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_106__A  (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_107__A  (.DIODE(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_108__A  (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_109__A  (.DIODE(net222),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_110__A  (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_111__A  (.DIODE(net224),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/_112__A  (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0_A2  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1_A1  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1_A2  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2_A2  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3_A0  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3_A1  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3_A2  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3_A3  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0_A2  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1_A1  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1_A2  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2_A2  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3_A0  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3_A1  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3_A2  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3_A3  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0_A3  (.DIODE(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1_A1  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1_A2  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0_A3  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1_A0  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1_A1  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1_A2  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1_A3  (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0_A3  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1_A1  (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1_A2  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0_A3  (.DIODE(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1_A0  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1_A1  (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1_A2  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1_A3  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0_A1  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0_A2  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0_A3  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1_A1  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1_A2  (.DIODE(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1_A3  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0_A1  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0_A2  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0_A3  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1_A1  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1_A2  (.DIODE(net164),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0_A1  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0_A2  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0_A3  (.DIODE(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1_A1  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1_A2  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0_A1  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0_A2  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0_A3  (.DIODE(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1_A1  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1_A2  (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1_A3  (.DIODE(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3_A2  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0_A3  (.DIODE(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1_A1  (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1_A2  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0_A3  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1_A0  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1_A1  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1_A2  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1_A3  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0_A3  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1_A1  (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1_A2  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1_A3  (.DIODE(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0_A3  (.DIODE(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1_A0  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1_A1  (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1_A2  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1_A3  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0_A1  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0_A2  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0_A3  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1_A1  (.DIODE(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0_A1  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0_A2  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0_A3  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1_A0  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1_A1  (.DIODE(net164),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0_A1  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0_A2  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0_A3  (.DIODE(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1_A0  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1_A1  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0_A1  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0_A2  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0_A3  (.DIODE(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1_A1  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3_A2  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0_A3  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1_A0  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1_A1  (.DIODE(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1_A2  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0_A3  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1_A0  (.DIODE(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1_A1  (.DIODE(net198),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1_A2  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1_A3  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0_A3  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1_A0  (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1_A1  (.DIODE(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1_A2  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0_A3  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1_A0  (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1_A1  (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1_A2  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1_A3  (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0_A1  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0_A2  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0_A3  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1_A1  (.DIODE(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0_A1  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0_A2  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0_A3  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1_A0  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1_A1  (.DIODE(net164),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0_A1  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0_A2  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0_A3  (.DIODE(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1_A0  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1_A1  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0_A1  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0_A2  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0_A3  (.DIODE(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1_A1  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3_A2  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0_A3  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1_A0  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1_A1  (.DIODE(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1_A2  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0_A3  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1_A0  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1_A1  (.DIODE(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1_A2  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1_A3  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0_A3  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1_A0  (.DIODE(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1_A1  (.DIODE(net199),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1_A2  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1_A3  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2_A2  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0_A3  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1_A0  (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1_A1  (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1_A2  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1_A3  (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0_A1  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0_A2  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0_A3  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1_A1  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1_A2  (.DIODE(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1_A3  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3_A3  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0_A1  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0_A2  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0_A3  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1_A1  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1_A2  (.DIODE(net164),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1_A3  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3_A1  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0_A1  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0_A2  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0_A3  (.DIODE(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1_A0  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1_A1  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1_A2  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1_A3  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3_A2  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0_A1  (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0_A2  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0_A3  (.DIODE(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1_A0  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1_A1  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1_A2  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1_A3  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2_A1  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2_A2  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3_A1  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3_A2  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3_A3  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0_A2  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1_A1  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1_A2  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2_A1  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2_A2  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2_A3  (.DIODE(M_AH),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3_A0  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3_A1  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3_A2  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3_A3  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0_A2  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1_A1  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1_A2  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2_A1  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2_A2  (.DIODE(M_AD),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2_A3  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3_A0  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3_A1  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3_A2  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3_A3  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_EN/_0__A1  (.DIODE(J_EN_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_SR/_0__A1  (.DIODE(J_SR_BEG),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG0_A0  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG0_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG0_A2  (.DIODE(\JN2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG0_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG1_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG1_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG1_A2  (.DIODE(\JN2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG1_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG2_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG2_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG2_A2  (.DIODE(\JN2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG2_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG3_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG3_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG3_A2  (.DIODE(\JN2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG3_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0_A0  (.DIODE(net112),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0_A1  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0_A2  (.DIODE(net199),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0_A3  (.DIODE(net216),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1_A0  (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1_A1  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1_A2  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1_A3  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2_A1  (.DIODE(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2_A2  (.DIODE(net162),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2_A3  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3_A0  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3_A1  (.DIODE(net6),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3_A2  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3_A3  (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0_A0  (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0_A1  (.DIODE(net12),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0_A2  (.DIODE(net164),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0_A3  (.DIODE(net216),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1_A0  (.DIODE(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1_A1  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1_A2  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1_A3  (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2_A1  (.DIODE(net10),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2_A2  (.DIODE(net198),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2_A3  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3_A0  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3_A1  (.DIODE(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3_A2  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3_A3  (.DIODE(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0_A0  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0_A1  (.DIODE(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0_A2  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0_A3  (.DIODE(net217),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1_A0  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1_A1  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1_A2  (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1_A3  (.DIODE(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2_A0  (.DIODE(net111),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2_A1  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2_A2  (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2_A3  (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3_A1  (.DIODE(net7),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3_A2  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3_A3  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0_A0  (.DIODE(net113),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0_A1  (.DIODE(net13),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0_A2  (.DIODE(net165),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0_A3  (.DIODE(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1_A0  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1_A1  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1_A2  (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1_A3  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2_A1  (.DIODE(net11),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2_A2  (.DIODE(net163),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2_A3  (.DIODE(net215),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3_A0  (.DIODE(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3_A1  (.DIODE(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3_A2  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3_A3  (.DIODE(net211),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0_A0  (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0_A1  (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0_A2  (.DIODE(net224),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0_A3  (.DIODE(\JN2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1_A0  (.DIODE(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1_A1  (.DIODE(net168),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1_A2  (.DIODE(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1_A3  (.DIODE(\JE2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2_A0  (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2_A1  (.DIODE(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2_A2  (.DIODE(net222),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2_A3  (.DIODE(\JS2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3_A0  (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3_A1  (.DIODE(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3_A2  (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3_A3  (.DIODE(\JW2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0_A0  (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0_A1  (.DIODE(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0_A2  (.DIODE(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0_A3  (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1_A0  (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1_A1  (.DIODE(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1_A2  (.DIODE(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1_A3  (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2_A0  (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2_A1  (.DIODE(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2_A2  (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2_A3  (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3_A0  (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3_A1  (.DIODE(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3_A2  (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3_A3  (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0_A0  (.DIODE(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0_A1  (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0_A2  (.DIODE(net224),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0_A3  (.DIODE(\JN2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1_A0  (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1_A1  (.DIODE(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1_A2  (.DIODE(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1_A3  (.DIODE(\JE2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2_A0  (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2_A1  (.DIODE(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2_A2  (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2_A3  (.DIODE(\JS2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3_A0  (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3_A1  (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3_A2  (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3_A3  (.DIODE(\JW2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0_A0  (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0_A1  (.DIODE(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0_A2  (.DIODE(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0_A3  (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1_A0  (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1_A1  (.DIODE(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1_A2  (.DIODE(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1_A3  (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2_A0  (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2_A1  (.DIODE(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2_A2  (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2_A3  (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3_A0  (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3_A1  (.DIODE(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3_A2  (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3_A3  (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0_A0  (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0_A1  (.DIODE(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0_A2  (.DIODE(net224),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1_A0  (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1_A1  (.DIODE(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1_A2  (.DIODE(net168),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1_A3  (.DIODE(\JE2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2_A0  (.DIODE(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2_A1  (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2_A2  (.DIODE(net222),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2_A3  (.DIODE(\JS2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3_A0  (.DIODE(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3_A1  (.DIODE(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3_A2  (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3_A3  (.DIODE(\JW2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0_A0  (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0_A1  (.DIODE(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0_A2  (.DIODE(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0_A3  (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1_A0  (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1_A1  (.DIODE(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1_A2  (.DIODE(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1_A3  (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2_A0  (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2_A1  (.DIODE(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2_A2  (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2_A3  (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3_A0  (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3_A1  (.DIODE(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3_A2  (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3_A3  (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0_A0  (.DIODE(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0_A1  (.DIODE(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0_A2  (.DIODE(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0_A3  (.DIODE(\JN2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1_A0  (.DIODE(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1_A1  (.DIODE(net168),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1_A2  (.DIODE(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1_A3  (.DIODE(\JE2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2_A0  (.DIODE(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2_A1  (.DIODE(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2_A2  (.DIODE(net222),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2_A3  (.DIODE(\JS2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3_A0  (.DIODE(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3_A1  (.DIODE(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3_A2  (.DIODE(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3_A3  (.DIODE(\JW2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0_A0  (.DIODE(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0_A1  (.DIODE(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0_A2  (.DIODE(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0_A3  (.DIODE(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1_A0  (.DIODE(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1_A1  (.DIODE(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1_A2  (.DIODE(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1_A3  (.DIODE(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2_A0  (.DIODE(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2_A1  (.DIODE(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2_A2  (.DIODE(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2_A3  (.DIODE(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3_A0  (.DIODE(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3_A1  (.DIODE(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3_A2  (.DIODE(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3_A3  (.DIODE(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0_A0  (.DIODE(net147),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0_A1  (.DIODE(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0_A2  (.DIODE(net238),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0_A3  (.DIODE(\JN2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1_A0  (.DIODE(net42),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1_A1  (.DIODE(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1_A2  (.DIODE(net217),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1_A3  (.DIODE(\JE2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2_A0  (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2_A1  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2_A2  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2_A3  (.DIODE(\JS2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3_A0  (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3_A1  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3_A2  (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3_A3  (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0_A0  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0_A1  (.DIODE(net199),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0_A2  (.DIODE(net246),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0_A3  (.DIODE(\JN2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1_A0  (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1_A1  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1_A2  (.DIODE(net217),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1_A3  (.DIODE(\JE2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2_A1  (.DIODE(net41),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2_A2  (.DIODE(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2_A3  (.DIODE(\JS2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3_A0  (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3_A1  (.DIODE(net190),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3_A2  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3_A3  (.DIODE(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0_A0  (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0_A1  (.DIODE(net9),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0_A2  (.DIODE(net213),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0_A3  (.DIODE(\JN2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1_A1  (.DIODE(net8),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1_A2  (.DIODE(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1_A3  (.DIODE(\JE2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2_A0  (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2_A1  (.DIODE(net197),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2_A2  (.DIODE(net214),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2_A3  (.DIODE(\JS2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3_A0  (.DIODE(net43),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3_A1  (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3_A2  (.DIODE(net245),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3_A3  (.DIODE(\JW2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0_A0  (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0_A1  (.DIODE(net34),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0_A2  (.DIODE(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0_A3  (.DIODE(\JN2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1_A0  (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1_A1  (.DIODE(net198),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1_A2  (.DIODE(net212),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1_A3  (.DIODE(\JE2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2_A1  (.DIODE(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2_A2  (.DIODE(net247),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2_A3  (.DIODE(\JS2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3_A0  (.DIODE(net138),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3_A1  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3_A2  (.DIODE(net210),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3_A3  (.DIODE(\JW2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I0_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I1_A2  (.DIODE(\J2END_AB_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I2_A0  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I2_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I2_A2  (.DIODE(\J2END_AB_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I0_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I1_A2  (.DIODE(\J2END_AB_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I2_A0  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I2_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I2_A2  (.DIODE(\J2END_AB_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I1_A1  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I1_A2  (.DIODE(\J2END_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I1_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I2_A0  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I2_A2  (.DIODE(\J2END_CD_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I3_A0  (.DIODE(\J2MID_CDa_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I3_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I3_A2  (.DIODE(\J2END_CD_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I1_A1  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I1_A2  (.DIODE(\J2END_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I1_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I2_A0  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I2_A2  (.DIODE(\J2END_CD_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I3_A0  (.DIODE(\J2MID_CDa_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I3_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I3_A2  (.DIODE(\J2END_CD_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I0_A0  (.DIODE(\J2MID_EFa_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I0_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I1_A2  (.DIODE(\J2END_EF_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I2_A0  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I2_A2  (.DIODE(\J2END_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I2_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I0_A0  (.DIODE(\J2MID_EFa_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I0_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I1_A2  (.DIODE(\J2END_EF_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I2_A0  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I2_A2  (.DIODE(\J2END_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I2_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I1_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I2_A0  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I2_A2  (.DIODE(\J2END_GH_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I3_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I1_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I2_A0  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I2_A2  (.DIODE(\J2END_GH_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I3_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG0_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG0_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG0_A2  (.DIODE(\JW2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG0_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG1_A0  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG1_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG1_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG2_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG2_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG2_A2  (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG2_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG3_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG3_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG3_A2  (.DIODE(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG3_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG0_A0  (.DIODE(net108),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG0_A1  (.DIODE(net129),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG0_A2  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG0_A3  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG1_A0  (.DIODE(net109),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG1_A1  (.DIODE(net130),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG1_A2  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG1_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG2_A0  (.DIODE(net106),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG2_A1  (.DIODE(net131),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG2_A2  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG2_A3  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG3_A0  (.DIODE(net107),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG3_A1  (.DIODE(net122),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG3_A2  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG3_A3  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S0_A0  (.DIODE(\JN2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S0_A1  (.DIODE(\JE2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S0_A2  (.DIODE(\JS2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S0_A3  (.DIODE(\JW2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG0_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG0_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG0_A2  (.DIODE(\JE2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG0_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG1_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG1_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG1_A2  (.DIODE(\JE2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG1_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG2_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG2_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG2_A2  (.DIODE(\JE2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG2_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG3_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG3_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG3_A2  (.DIODE(\JE2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG3_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1_A1  (.DIODE(\JE2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1_A2  (.DIODE(\JS2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1_A3  (.DIODE(\JW2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S2_A0  (.DIODE(\JN2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S2_A1  (.DIODE(\JE2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S2_A2  (.DIODE(\JS2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S2_A3  (.DIODE(\JW2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S3_A0  (.DIODE(\JN2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S3_A1  (.DIODE(\JE2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S3_A3  (.DIODE(\JW2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG0_A0  (.DIODE(net25),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG0_A1  (.DIODE(net160),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG0_A2  (.DIODE(net181),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG0_A3  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG1_A0  (.DIODE(net22),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG1_A1  (.DIODE(net161),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG1_A2  (.DIODE(net182),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG1_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG2_A0  (.DIODE(net158),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG2_A1  (.DIODE(net183),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG2_A2  (.DIODE(net229),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG2_A3  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG3_A0  (.DIODE(net159),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG3_A1  (.DIODE(net174),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG3_A2  (.DIODE(net226),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG3_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG0_A0  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG0_A1  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG0_A2  (.DIODE(\JS2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG0_A3  (.DIODE(\J_l_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG1_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG1_A1  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG1_A2  (.DIODE(\JS2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG1_A3  (.DIODE(\J_l_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG2_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG2_A1  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG2_A2  (.DIODE(\JS2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG2_A3  (.DIODE(\J_l_GH_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG3_A0  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG3_A1  (.DIODE(\J2MID_ABb_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG3_A2  (.DIODE(\JS2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG3_A3  (.DIODE(\J_l_AB_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst0_A2  (.DIODE(\J2MID_CDb_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst1_A0  (.DIODE(\JN2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\JE2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\JS2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst1_A3  (.DIODE(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst0_A3  (.DIODE(\J2MID_EFb_BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst1_A0  (.DIODE(\JN2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\JE2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\JS2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst1_A3  (.DIODE(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_EF_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_CD_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_AB_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net4),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net5),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_CD_BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0_A0  (.DIODE(net104),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0_A1  (.DIODE(net156),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0_A2  (.DIODE(net208),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0_A3  (.DIODE(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1_A0  (.DIODE(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_GH_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0_A0  (.DIODE(net105),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0_A1  (.DIODE(net157),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0_A2  (.DIODE(net209),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0_A3  (.DIODE(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1_A0  (.DIODE(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_ABa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_CDa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_EF_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0_A0  (.DIODE(net102),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0_A1  (.DIODE(net154),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0_A2  (.DIODE(net206),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0_A3  (.DIODE(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1_A0  (.DIODE(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHb_BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_CD_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0_A0  (.DIODE(net103),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0_A1  (.DIODE(net155),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0_A2  (.DIODE(net207),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0_A3  (.DIODE(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1_A0  (.DIODE(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1_A1  (.DIODE(\J2MID_EFa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1_A2  (.DIODE(\J2MID_GHa_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1_A3  (.DIODE(\J2END_AB_BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_MUX8LUT_frame_config_mux/cus_mux21_AD/_0__A0  (.DIODE(M_AB),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_Inst_MUX8LUT_frame_config_mux/cus_mux21_EH/_0__A0  (.DIODE(M_EF),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_0/_0__A  (.DIODE(\N4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_1/_0__A  (.DIODE(\N4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_10/_0__A  (.DIODE(\N4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_11/_0__A  (.DIODE(\N4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_2/_0__A  (.DIODE(\N4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_3/_0__A  (.DIODE(\N4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_4/_0__A  (.DIODE(\N4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_5/_0__A  (.DIODE(\N4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_6/_0__A  (.DIODE(\N4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_7/_0__A  (.DIODE(\N4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_8/_0__A  (.DIODE(\N4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_N4BEG_outbuf_9/_0__A  (.DIODE(\N4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_0/_0__A  (.DIODE(\NN4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_1/_0__A  (.DIODE(\NN4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_10/_0__A  (.DIODE(\NN4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_11/_0__A  (.DIODE(\NN4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_2/_0__A  (.DIODE(\NN4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_3/_0__A  (.DIODE(\NN4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_4/_0__A  (.DIODE(\NN4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_5/_0__A  (.DIODE(\NN4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_6/_0__A  (.DIODE(\NN4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_7/_0__A  (.DIODE(\NN4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_8/_0__A  (.DIODE(\NN4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_NN4BEG_outbuf_9/_0__A  (.DIODE(\NN4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_0/_0__A  (.DIODE(\S4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_1/_0__A  (.DIODE(\S4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_10/_0__A  (.DIODE(\S4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_11/_0__A  (.DIODE(\S4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_2/_0__A  (.DIODE(\S4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_3/_0__A  (.DIODE(\S4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_4/_0__A  (.DIODE(\S4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_5/_0__A  (.DIODE(\S4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_6/_0__A  (.DIODE(\S4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_7/_0__A  (.DIODE(\S4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_8/_0__A  (.DIODE(\S4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_S4BEG_outbuf_9/_0__A  (.DIODE(\S4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_0/_0__A  (.DIODE(\SS4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_1/_0__A  (.DIODE(\SS4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_10/_0__A  (.DIODE(\SS4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_11/_0__A  (.DIODE(\SS4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_2/_0__A  (.DIODE(\SS4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_3/_0__A  (.DIODE(\SS4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_4/_0__A  (.DIODE(\SS4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_5/_0__A  (.DIODE(\SS4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_6/_0__A  (.DIODE(\SS4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_7/_0__A  (.DIODE(\SS4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_8/_0__A  (.DIODE(\SS4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_SS4BEG_outbuf_9/_0__A  (.DIODE(\SS4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_0/_0__A  (.DIODE(\W6BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_1/_0__A  (.DIODE(\W6BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_2/_0__A  (.DIODE(\W6BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_3/_0__A  (.DIODE(\W6BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_4/_0__A  (.DIODE(\W6BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_5/_0__A  (.DIODE(\W6BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_6/_0__A  (.DIODE(\W6BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_7/_0__A  (.DIODE(\W6BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_8/_0__A  (.DIODE(\W6BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_W6BEG_outbuf_9/_0__A  (.DIODE(\W6BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_0/_0__A  (.DIODE(\WW4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_1/_0__A  (.DIODE(\WW4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_10/_0__A  (.DIODE(\WW4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_11/_0__A  (.DIODE(\WW4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_2/_0__A  (.DIODE(\WW4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_3/_0__A  (.DIODE(\WW4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_4/_0__A  (.DIODE(\WW4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_5/_0__A  (.DIODE(\WW4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_6/_0__A  (.DIODE(\WW4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_7/_0__A  (.DIODE(\WW4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_8/_0__A  (.DIODE(\WW4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_WW4BEG_outbuf_9/_0__A  (.DIODE(\WW4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_0/_0__A  (.DIODE(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_1/_0__A  (.DIODE(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_10/_0__A  (.DIODE(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_11/_0__A  (.DIODE(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_12/_0__A  (.DIODE(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_13/_0__A  (.DIODE(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_14/_0__A  (.DIODE(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_15/_0__A  (.DIODE(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_16/_0__A  (.DIODE(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_17/_0__A  (.DIODE(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_18/_0__A  (.DIODE(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_19/_0__A  (.DIODE(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_2/_0__A  (.DIODE(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_20/_0__A  (.DIODE(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_21/_0__A  (.DIODE(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_22/_0__A  (.DIODE(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_23/_0__A  (.DIODE(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_24/_0__A  (.DIODE(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_25/_0__A  (.DIODE(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_26/_0__A  (.DIODE(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_27/_0__A  (.DIODE(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_28/_0__A  (.DIODE(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_29/_0__A  (.DIODE(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_3/_0__A  (.DIODE(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_30/_0__A  (.DIODE(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_31/_0__A  (.DIODE(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_4/_0__A  (.DIODE(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_5/_0__A  (.DIODE(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_6/_0__A  (.DIODE(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_7/_0__A  (.DIODE(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_8/_0__A  (.DIODE(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data_inbuf_9/_0__A  (.DIODE(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output277_A (.DIODE(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output356_A (.DIODE(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_A (.DIODE(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output473_A (.DIODE(net473),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_A (.DIODE(net477),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_0/_0__A  (.DIODE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_1/_0__A  (.DIODE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_10/_0__A  (.DIODE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_11/_0__A  (.DIODE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_12/_0__A  (.DIODE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_13/_0__A  (.DIODE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_14/_0__A  (.DIODE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_15/_0__A  (.DIODE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_16/_0__A  (.DIODE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_17/_0__A  (.DIODE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_18/_0__A  (.DIODE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_19/_0__A  (.DIODE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_2/_0__A  (.DIODE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_3/_0__A  (.DIODE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_4/_0__A  (.DIODE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_5/_0__A  (.DIODE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_6/_0__A  (.DIODE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_7/_0__A  (.DIODE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_8/_0__A  (.DIODE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__diode_2 \ANTENNA_strobe_inbuf_9/_0__A  (.DIODE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_0/_0_  (.A(\E6BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_1/_0_  (.A(\E6BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_2/_0_  (.A(\E6BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_3/_0_  (.A(\E6BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_4/_0_  (.A(\E6BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_5/_0_  (.A(\E6BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_6/_0_  (.A(\E6BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_7/_0_  (.A(\E6BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_8/_0_  (.A(\E6BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 \E6BEG_outbuf_9/_0_  (.A(\E6BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_0/_0_  (.A(net26),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_1/_0_  (.A(net27),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_2/_0_  (.A(net28),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_3/_0_  (.A(net29),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_4/_0_  (.A(net30),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_5/_0_  (.A(net31),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_6/_0_  (.A(net32),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_7/_0_  (.A(net33),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_8/_0_  (.A(net23),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \E6END_inbuf_9/_0_  (.A(net24),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\E6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_0/_0_  (.A(\EE4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_1/_0_  (.A(\EE4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_10/_0_  (.A(\EE4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_11/_0_  (.A(\EE4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_2/_0_  (.A(\EE4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_3/_0_  (.A(\EE4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_4/_0_  (.A(\EE4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_5/_0_  (.A(\EE4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_6/_0_  (.A(\EE4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_7/_0_  (.A(\EE4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_8/_0_  (.A(\EE4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 \EE4BEG_outbuf_9/_0_  (.A(\EE4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_0/_0_  (.A(net44),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_1/_0_  (.A(net45),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_10/_0_  (.A(net39),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_11/_0_  (.A(net40),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_2/_0_  (.A(net46),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_3/_0_  (.A(net47),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_4/_0_  (.A(net48),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_5/_0_  (.A(net49),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_6/_0_  (.A(net35),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_7/_0_  (.A(net36),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_8/_0_  (.A(net37),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \EE4END_inbuf_9/_0_  (.A(net38),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\EE4BEG_i[9] ));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_422 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_347 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_366 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_339 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_462 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_398 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_470 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_339 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_394 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_398 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_364 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_312 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_336 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_376 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_466 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_32_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_398 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_34_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_426 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_34_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_34_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_34_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_290 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_35_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_35_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_35_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_36_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_36_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_343 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_36_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_36_463 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_36_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_36_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_252 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_37_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_372 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_37_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_37_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_37_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_38_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_38_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_38_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_38_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_38_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_39_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_39_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_39_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_40_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_40_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_379 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_40_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_40_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_40_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_308 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_312 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_41_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_41_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_41_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_41_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_41_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_41_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_224 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_42_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_42_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_42_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_42_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_42_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_42_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_43_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_423 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_43_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_43_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_43_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_44_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_44_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_314 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_44_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_433 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_44_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_44_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_44_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_45_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_312 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_45_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_45_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_45_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_46_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_46_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_46_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_46_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_46_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_47_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_367 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_47_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_47_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_47_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_47_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_47_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_48_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_48_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_48_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_48_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_48_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_49_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_49_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_49_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_49_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_211 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_267 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_283 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_371 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_404 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_50_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_50_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_50_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_51_366 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_51_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_51_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_51_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_51_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_223 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_52_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_52_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_52_459 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_310 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_407 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_53_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_53_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_53_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_54_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_54_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_54_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_54_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_157 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_55_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_426 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_55_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_55_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_55_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_185 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_56_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_227 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_275 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_294 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_298 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_56_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_56_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_56_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_56_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_177 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_198 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_57_405 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_423 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_57_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_57_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_57_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_318 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_322 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_58_375 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_58_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_58_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_296 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_59_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_59_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_59_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_59_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_208 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_291 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_303 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_364 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_370 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_261 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_60_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_305 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_60_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_60_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_60_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_182 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_246 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_61_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_61_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_61_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_61_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_62_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_424 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_62_467 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_62_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_174 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_245 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_289 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_297 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_356 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_366 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_420 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_63_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_63_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_63_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_64_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_64_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_346 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_429 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_64_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_64_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_64_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_64_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_162 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_237 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_256 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_65_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_65_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_65_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_65_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_192 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_209 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_217 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_66_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_66_236 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_282 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_352 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_66_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_66_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_451 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_66_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_66_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_238 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_260 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_293 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_316 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_320 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_354 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_67_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_67_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_67_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_67_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_67_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_67_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_168 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_280 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_68_338 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_68_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_392 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_68_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_455 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_68_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_68_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_68_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_68_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_241 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_69_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_288 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_292 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_384 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_69_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_441 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_69_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_69_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_69_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_193 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_214 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_243 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_247 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_257 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_340 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_426 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_430 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_434 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_448 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_464 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_472 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_159 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_163 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_380 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_70_403 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_411 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_432 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_70_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_70_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_70_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_70_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_204 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_216 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_229 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_235 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_239 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_258 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_262 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_266 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_408 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_412 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_71_416 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_428 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_474 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_71_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_71_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_71_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_71_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_176 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_180 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_212 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_234 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_72_242 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_265 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_269 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_302 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_306 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_313 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_321 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_333 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_351 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_388 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_409 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_415 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_439 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_443 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_450 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_454 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_458 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_468 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_72_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_72_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_72_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_178 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_190 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_202 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_210 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_215 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_263 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_271 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_373 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_386 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_396 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_73_400 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_73_425 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_73_437 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_73_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_73_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_158 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_161 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_165 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_171 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_179 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_184 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_188 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_201 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_249 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_328 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_344 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_348 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_355 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_359 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_368 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_402 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_406 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_410 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_427 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_431 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_74_435 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_447 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_74_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_74_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_74_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_74_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_172 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_196 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_200 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_203 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_207 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_219 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_273 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_285 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_295 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_301 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_438 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_75_442 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_8 FILLER_0_75_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_75_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_75_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_75_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_75_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_186 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_206 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_76_220 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_362 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_377 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_76_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_76_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_173 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_197 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_231 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_299 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_307 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_324 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_350 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_77_381 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_77_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_77_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_77_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_156 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_160 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_169 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_175 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_181 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_213 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_264 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_268 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_272 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_276 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_311 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_315 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_319 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_323 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_327 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_331 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_358 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_414 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_418 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_422 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_426 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_436 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_440 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_465 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_469 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_473 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_167 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_183 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_189 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_218 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_222 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_226 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_230 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_233 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_270 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_274 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_278 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_284 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_325 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_329 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_369 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_374 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_378 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_382 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_399 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_421 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_452 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_456 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_460 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_187 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_191 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_195 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_199 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_205 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_240 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_244 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_248 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_251 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_255 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_259 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_287 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_326 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_330 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_337 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_341 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_345 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_349 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_353 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_357 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_361 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_365 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_383 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_387 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_397 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_401 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_453 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_457 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_461 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr/_08_  (.A(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr/_09_  (.A(LA_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LA_LUT4c_frame_config_dffesr/_10_  (.A(LA_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LA_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LA_LUT4c_frame_config_dffesr/_11_  (.A1(LA_I2),
    .A2(LA_Ci),
    .B1(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LA_LUT4c_frame_config_dffesr/_12_  (.A1(LA_I2),
    .A2(LA_Ci),
    .B1(\Inst_LA_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LA_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LA_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[18] ),
    .S(LA_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LA_LUT4c_frame_config_dffesr/_14_  (.A0(net531),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr/_06_ ),
    .S(LA_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LA_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LA_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LA_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LA_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LA_I0),
    .A1(LA_Ci),
    .S(\ConfigBits[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LA_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LA_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[0] ),
    .A1(\ConfigBits[1] ),
    .A2(\ConfigBits[2] ),
    .A3(\ConfigBits[3] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[4] ),
    .A1(\ConfigBits[5] ),
    .A2(\ConfigBits[6] ),
    .A3(\ConfigBits[7] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[8] ),
    .A1(\ConfigBits[9] ),
    .A2(\ConfigBits[10] ),
    .A3(\ConfigBits[11] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[12] ),
    .A1(\ConfigBits[13] ),
    .A2(\ConfigBits[14] ),
    .A3(\ConfigBits[15] ),
    .S0(\Inst_LA_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LA_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LA_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LA_I2),
    .S1(LA_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LA_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr/_08_  (.A(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr/_09_  (.A(LB_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LB_LUT4c_frame_config_dffesr/_10_  (.A(LB_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LB_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LB_LUT4c_frame_config_dffesr/_11_  (.A1(LB_I2),
    .A2(LB_Ci),
    .B1(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LB_LUT4c_frame_config_dffesr/_12_  (.A1(LB_I2),
    .A2(LB_Ci),
    .B1(\Inst_LB_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LB_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LB_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[37] ),
    .S(LB_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LB_LUT4c_frame_config_dffesr/_14_  (.A0(net526),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr/_06_ ),
    .S(LB_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LB_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LB_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LB_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LB_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LB_I0),
    .A1(LB_Ci),
    .S(\ConfigBits[36] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LB_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LB_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[35] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[19] ),
    .A1(\ConfigBits[20] ),
    .A2(\ConfigBits[21] ),
    .A3(\ConfigBits[22] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[23] ),
    .A1(\ConfigBits[24] ),
    .A2(\ConfigBits[25] ),
    .A3(\ConfigBits[26] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[27] ),
    .A1(\ConfigBits[28] ),
    .A2(\ConfigBits[29] ),
    .A3(\ConfigBits[30] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[31] ),
    .A1(\ConfigBits[32] ),
    .A2(\ConfigBits[33] ),
    .A3(\ConfigBits[34] ),
    .S0(\Inst_LB_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LB_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LB_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LB_I2),
    .S1(LB_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LB_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr/_08_  (.A(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr/_09_  (.A(LC_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LC_LUT4c_frame_config_dffesr/_10_  (.A(LC_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LC_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LC_LUT4c_frame_config_dffesr/_11_  (.A1(LC_I2),
    .A2(LC_Ci),
    .B1(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LC_LUT4c_frame_config_dffesr/_12_  (.A1(LC_I2),
    .A2(LC_Ci),
    .B1(\Inst_LC_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LC_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LC_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[56] ),
    .S(LC_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LC_LUT4c_frame_config_dffesr/_14_  (.A0(net529),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr/_06_ ),
    .S(LC_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LC_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LC_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LC_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LC_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LC_I0),
    .A1(LC_Ci),
    .S(\ConfigBits[55] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LC_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LC_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[54] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[38] ),
    .A1(\ConfigBits[39] ),
    .A2(\ConfigBits[40] ),
    .A3(\ConfigBits[41] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[42] ),
    .A1(\ConfigBits[43] ),
    .A2(\ConfigBits[44] ),
    .A3(\ConfigBits[45] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[46] ),
    .A1(\ConfigBits[47] ),
    .A2(\ConfigBits[48] ),
    .A3(\ConfigBits[49] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[50] ),
    .A1(\ConfigBits[51] ),
    .A2(\ConfigBits[52] ),
    .A3(\ConfigBits[53] ),
    .S0(\Inst_LC_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LC_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LC_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LC_I2),
    .S1(LC_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LC_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr/_08_  (.A(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr/_09_  (.A(LD_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LD_LUT4c_frame_config_dffesr/_10_  (.A(LD_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LD_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LD_LUT4c_frame_config_dffesr/_11_  (.A1(LD_I2),
    .A2(LD_Ci),
    .B1(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LD_LUT4c_frame_config_dffesr/_12_  (.A1(LD_I2),
    .A2(LD_Ci),
    .B1(\Inst_LD_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LD_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LD_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[75] ),
    .S(LD_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LD_LUT4c_frame_config_dffesr/_14_  (.A0(net530),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr/_06_ ),
    .S(LD_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LD_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LD_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LD_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LD_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LD_I0),
    .A1(LD_Ci),
    .S(\ConfigBits[74] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LD_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LD_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[73] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[57] ),
    .A1(\ConfigBits[58] ),
    .A2(\ConfigBits[59] ),
    .A3(\ConfigBits[60] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[61] ),
    .A1(\ConfigBits[62] ),
    .A2(\ConfigBits[63] ),
    .A3(\ConfigBits[64] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[65] ),
    .A1(\ConfigBits[66] ),
    .A2(\ConfigBits[67] ),
    .A3(\ConfigBits[68] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[69] ),
    .A1(\ConfigBits[70] ),
    .A2(\ConfigBits[71] ),
    .A3(\ConfigBits[72] ),
    .S0(\Inst_LD_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LD_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LD_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LD_I2),
    .S1(LD_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LD_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr/_08_  (.A(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr/_09_  (.A(LE_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LE_LUT4c_frame_config_dffesr/_10_  (.A(LE_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LE_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LE_LUT4c_frame_config_dffesr/_11_  (.A1(LE_I2),
    .A2(LE_Ci),
    .B1(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LE_LUT4c_frame_config_dffesr/_12_  (.A1(LE_I2),
    .A2(LE_Ci),
    .B1(\Inst_LE_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LE_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LE_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[94] ),
    .S(LE_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LE_LUT4c_frame_config_dffesr/_14_  (.A0(net524),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr/_06_ ),
    .S(LE_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LE_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LE_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LE_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LE_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LE_I0),
    .A1(LE_Ci),
    .S(\ConfigBits[93] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LE_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LE_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[92] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[76] ),
    .A1(\ConfigBits[77] ),
    .A2(\ConfigBits[78] ),
    .A3(\ConfigBits[79] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[80] ),
    .A1(\ConfigBits[81] ),
    .A2(\ConfigBits[82] ),
    .A3(\ConfigBits[83] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[84] ),
    .A1(\ConfigBits[85] ),
    .A2(\ConfigBits[86] ),
    .A3(\ConfigBits[87] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[88] ),
    .A1(\ConfigBits[89] ),
    .A2(\ConfigBits[90] ),
    .A3(\ConfigBits[91] ),
    .S0(\Inst_LE_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LE_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LE_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LE_I2),
    .S1(LE_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LE_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr/_08_  (.A(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr/_09_  (.A(LF_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LF_LUT4c_frame_config_dffesr/_10_  (.A(LF_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LF_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LF_LUT4c_frame_config_dffesr/_11_  (.A1(LF_I2),
    .A2(LF_Ci),
    .B1(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LF_LUT4c_frame_config_dffesr/_12_  (.A1(LF_I2),
    .A2(LF_Ci),
    .B1(\Inst_LF_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LF_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LF_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[113] ),
    .S(LF_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LF_LUT4c_frame_config_dffesr/_14_  (.A0(net528),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr/_06_ ),
    .S(LF_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LF_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LF_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LF_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LF_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LF_I0),
    .A1(LF_Ci),
    .S(\ConfigBits[112] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LF_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LF_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[111] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[95] ),
    .A1(\ConfigBits[96] ),
    .A2(\ConfigBits[97] ),
    .A3(\ConfigBits[98] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[99] ),
    .A1(\ConfigBits[100] ),
    .A2(\ConfigBits[101] ),
    .A3(\ConfigBits[102] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[103] ),
    .A1(\ConfigBits[104] ),
    .A2(\ConfigBits[105] ),
    .A3(\ConfigBits[106] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[107] ),
    .A1(\ConfigBits[108] ),
    .A2(\ConfigBits[109] ),
    .A3(\ConfigBits[110] ),
    .S0(\Inst_LF_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LF_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LF_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LF_I2),
    .S1(LF_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LF_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr/_08_  (.A(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr/_09_  (.A(LG_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LG_LUT4c_frame_config_dffesr/_10_  (.A(LG_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LG_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LG_LUT4c_frame_config_dffesr/_11_  (.A1(LG_I2),
    .A2(LG_Ci),
    .B1(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LG_LUT4c_frame_config_dffesr/_12_  (.A1(LG_I2),
    .A2(LG_Ci),
    .B1(\Inst_LG_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LG_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LG_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[132] ),
    .S(LG_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LG_LUT4c_frame_config_dffesr/_14_  (.A0(net527),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr/_06_ ),
    .S(LG_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LG_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LG_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LG_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LG_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LG_I0),
    .A1(LG_Ci),
    .S(\ConfigBits[131] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LG_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LG_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[130] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[114] ),
    .A1(\ConfigBits[115] ),
    .A2(\ConfigBits[116] ),
    .A3(\ConfigBits[117] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[118] ),
    .A1(\ConfigBits[119] ),
    .A2(\ConfigBits[120] ),
    .A3(\ConfigBits[121] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[122] ),
    .A1(\ConfigBits[123] ),
    .A2(\ConfigBits[124] ),
    .A3(\ConfigBits[125] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[126] ),
    .A1(\ConfigBits[127] ),
    .A2(\ConfigBits[128] ),
    .A3(\ConfigBits[129] ),
    .S0(\Inst_LG_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LG_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LG_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LG_I2),
    .S1(LG_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LG_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr/_07_  (.A(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr/_00_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr/_08_  (.A(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr/_01_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr/_09_  (.A(LH_I2),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr/_02_ ));
 sky130_fd_sc_hd__inv_2 \Inst_LH_LUT4c_frame_config_dffesr/_10_  (.A(LH_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Y(\Inst_LH_LUT4c_frame_config_dffesr/_03_ ));
 sky130_fd_sc_hd__o21a_1 \Inst_LH_LUT4c_frame_config_dffesr/_11_  (.A1(LH_I2),
    .A2(LH_Ci),
    .B1(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/_05_ ));
 sky130_fd_sc_hd__a21o_1 \Inst_LH_LUT4c_frame_config_dffesr/_12_  (.A1(LH_I2),
    .A2(LH_Ci),
    .B1(\Inst_LH_LUT4c_frame_config_dffesr/_05_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_Co));
 sky130_fd_sc_hd__mux2_1 \Inst_LH_LUT4c_frame_config_dffesr/_13_  (.A0(\Inst_LH_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\ConfigBits[151] ),
    .S(LH_SR),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/_06_ ));
 sky130_fd_sc_hd__mux2_1 \Inst_LH_LUT4c_frame_config_dffesr/_14_  (.A0(net525),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr/_06_ ),
    .S(LH_EN),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/_04_ ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_LH_LUT4c_frame_config_dffesr/_15_  (.CLK(UserCLK),
    .D(\Inst_LH_LUT4c_frame_config_dffesr/_04_ ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\Inst_LH_LUT4c_frame_config_dffesr/LUT_flop ));
 sky130_fd_sc_hd__mux2_2 \Inst_LH_LUT4c_frame_config_dffesr/cus_mux21_I0mux/_0_  (.A0(LH_I0),
    .A1(LH_Ci),
    .S(\ConfigBits[150] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ));
 sky130_fd_sc_hd__mux2_8 \Inst_LH_LUT4c_frame_config_dffesr/cus_mux21_O/_0_  (.A0(\Inst_LH_LUT4c_frame_config_dffesr/LUT_out ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr/LUT_flop ),
    .S(\ConfigBits[149] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_O));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst0  (.A0(\ConfigBits[133] ),
    .A1(\ConfigBits[134] ),
    .A2(\ConfigBits[135] ),
    .A3(\ConfigBits[136] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst1  (.A0(\ConfigBits[137] ),
    .A1(\ConfigBits[138] ),
    .A2(\ConfigBits[139] ),
    .A3(\ConfigBits[140] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst2  (.A0(\ConfigBits[141] ),
    .A1(\ConfigBits[142] ),
    .A2(\ConfigBits[143] ),
    .A3(\ConfigBits[144] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst3  (.A0(\ConfigBits[145] ),
    .A1(\ConfigBits[146] ),
    .A2(\ConfigBits[147] ),
    .A3(\ConfigBits[148] ),
    .S0(\Inst_LH_LUT4c_frame_config_dffesr/I0mux ),
    .S1(LH_I1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_inst4  (.A0(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out0 ),
    .A1(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out1 ),
    .A2(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out2 ),
    .A3(\Inst_LH_LUT4c_frame_config_dffesr/inst_cus_mux161_buf/cus_mux41_buf_out3 ),
    .S0(LH_I2),
    .S1(LH_I3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LH_LUT4c_frame_config_dffesr/LUT_out ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit0  (.D(net50),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[389] ),
    .Q_N(\ConfigBits_N[389] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit1  (.D(net61),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[397] ),
    .Q_N(\ConfigBits_N[397] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit10  (.D(net51),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[577] ),
    .Q_N(\ConfigBits_N[577] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit11  (.D(net52),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[576] ),
    .Q_N(\ConfigBits_N[576] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit12  (.D(net53),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[568] ),
    .Q_N(\ConfigBits_N[568] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit13  (.D(net54),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[159] ),
    .Q_N(\ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit14  (.D(net55),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[158] ),
    .Q_N(\ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit15  (.D(net56),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[157] ),
    .Q_N(\ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit16  (.D(net57),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[241] ),
    .Q_N(\ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit17  (.D(net58),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[240] ),
    .Q_N(\ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit18  (.D(net59),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[263] ),
    .Q_N(\ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit19  (.D(net60),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[261] ),
    .Q_N(\ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit20  (.D(net62),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[259] ),
    .Q_N(\ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit21  (.D(net63),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[248] ),
    .Q_N(\ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit22  (.D(net64),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[247] ),
    .Q_N(\ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit23  (.D(net65),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[243] ),
    .Q_N(\ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit24  (.D(net66),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[242] ),
    .Q_N(\ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit3  (.D(net75),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[413] ),
    .Q_N(\ConfigBits_N[413] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit4  (.D(net76),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[462] ),
    .Q_N(\ConfigBits_N[462] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit5  (.D(net77),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[481] ),
    .Q_N(\ConfigBits_N[481] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit6  (.D(net78),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[473] ),
    .Q_N(\ConfigBits_N[473] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit7  (.D(net79),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[472] ),
    .Q_N(\ConfigBits_N[472] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit8  (.D(net80),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[502] ),
    .Q_N(\ConfigBits_N[502] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame0_bit9  (.D(net81),
    .GATE(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[558] ),
    .Q_N(\ConfigBits_N[558] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit0  (.D(net50),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[330] ),
    .Q_N(\ConfigBits_N[330] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit1  (.D(net61),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[338] ),
    .Q_N(\ConfigBits_N[338] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit10  (.D(net51),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[395] ),
    .Q_N(\ConfigBits_N[395] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit11  (.D(net52),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[411] ),
    .Q_N(\ConfigBits_N[411] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit12  (.D(net53),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[557] ),
    .Q_N(\ConfigBits_N[557] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit13  (.D(net54),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[581] ),
    .Q_N(\ConfigBits_N[581] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit14  (.D(net55),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[63] ),
    .Q_N(\ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit15  (.D(net56),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[133] ),
    .Q_N(\ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit16  (.D(net57),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[127] ),
    .Q_N(\ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit17  (.D(net58),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[118] ),
    .Q_N(\ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit18  (.D(net59),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[117] ),
    .Q_N(\ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit19  (.D(net60),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[115] ),
    .Q_N(\ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit2  (.D(net72),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[391] ),
    .Q_N(\ConfigBits_N[391] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit20  (.D(net62),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[139] ),
    .Q_N(\ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit21  (.D(net63),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[199] ),
    .Q_N(\ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit22  (.D(net64),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[196] ),
    .Q_N(\ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit23  (.D(net65),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[222] ),
    .Q_N(\ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit24  (.D(net66),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[221] ),
    .Q_N(\ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit25  (.D(net67),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[220] ),
    .Q_N(\ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit26  (.D(net68),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[200] ),
    .Q_N(\ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit27  (.D(net69),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[232] ),
    .Q_N(\ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit28  (.D(net70),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[271] ),
    .Q_N(\ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit29  (.D(net71),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[270] ),
    .Q_N(\ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit3  (.D(net75),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[390] ),
    .Q_N(\ConfigBits_N[390] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit30  (.D(net73),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[615] ),
    .Q_N(\ConfigBits_N[615] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit31  (.D(net74),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[601] ),
    .Q_N(\ConfigBits_N[601] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit4  (.D(net76),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[381] ),
    .Q_N(\ConfigBits_N[381] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit5  (.D(net77),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[380] ),
    .Q_N(\ConfigBits_N[380] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit6  (.D(net78),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[377] ),
    .Q_N(\ConfigBits_N[377] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit7  (.D(net79),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[376] ),
    .Q_N(\ConfigBits_N[376] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit8  (.D(net80),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[360] ),
    .Q_N(\ConfigBits_N[360] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame10_bit9  (.D(net81),
    .GATE(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[398] ),
    .Q_N(\ConfigBits_N[398] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit0  (.D(net50),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[322] ),
    .Q_N(\ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit1  (.D(net61),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[318] ),
    .Q_N(\ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit10  (.D(net51),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[416] ),
    .Q_N(\ConfigBits_N[416] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit11  (.D(net52),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[394] ),
    .Q_N(\ConfigBits_N[394] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit12  (.D(net53),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[410] ),
    .Q_N(\ConfigBits_N[410] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit13  (.D(net54),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[403] ),
    .Q_N(\ConfigBits_N[403] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit14  (.D(net55),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[521] ),
    .Q_N(\ConfigBits_N[521] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit15  (.D(net56),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[134] ),
    .Q_N(\ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit16  (.D(net57),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[128] ),
    .Q_N(\ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit17  (.D(net58),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[120] ),
    .Q_N(\ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit18  (.D(net59),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[114] ),
    .Q_N(\ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit19  (.D(net60),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[140] ),
    .Q_N(\ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit2  (.D(net72),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[296] ),
    .Q_N(\ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit20  (.D(net62),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[138] ),
    .Q_N(\ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit21  (.D(net63),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[151] ),
    .Q_N(\ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit22  (.D(net64),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[198] ),
    .Q_N(\ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit23  (.D(net65),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[188] ),
    .Q_N(\ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit24  (.D(net66),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[187] ),
    .Q_N(\ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit25  (.D(net67),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[201] ),
    .Q_N(\ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit26  (.D(net68),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[234] ),
    .Q_N(\ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit27  (.D(net69),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[233] ),
    .Q_N(\ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit28  (.D(net70),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[610] ),
    .Q_N(\ConfigBits_N[610] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit29  (.D(net71),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[602] ),
    .Q_N(\ConfigBits_N[602] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit3  (.D(net75),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[332] ),
    .Q_N(\ConfigBits_N[332] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit30  (.D(net73),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[585] ),
    .Q_N(\ConfigBits_N[585] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit31  (.D(net74),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[584] ),
    .Q_N(\ConfigBits_N[584] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit4  (.D(net76),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[331] ),
    .Q_N(\ConfigBits_N[331] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit5  (.D(net77),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[355] ),
    .Q_N(\ConfigBits_N[355] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit6  (.D(net78),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[339] ),
    .Q_N(\ConfigBits_N[339] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit7  (.D(net79),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[387] ),
    .Q_N(\ConfigBits_N[387] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit8  (.D(net80),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[400] ),
    .Q_N(\ConfigBits_N[400] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame11_bit9  (.D(net81),
    .GATE(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[417] ),
    .Q_N(\ConfigBits_N[417] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit0  (.D(net50),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[327] ),
    .Q_N(\ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit1  (.D(net61),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[297] ),
    .Q_N(\ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit10  (.D(net51),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[39] ),
    .Q_N(\ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit11  (.D(net52),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[28] ),
    .Q_N(\ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit12  (.D(net53),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[135] ),
    .Q_N(\ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit13  (.D(net54),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[131] ),
    .Q_N(\ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit14  (.D(net55),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[123] ),
    .Q_N(\ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit15  (.D(net56),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[122] ),
    .Q_N(\ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit16  (.D(net57),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[116] ),
    .Q_N(\ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit17  (.D(net58),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[143] ),
    .Q_N(\ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit18  (.D(net59),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[150] ),
    .Q_N(\ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit19  (.D(net60),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[148] ),
    .Q_N(\ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit2  (.D(net72),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[337] ),
    .Q_N(\ConfigBits_N[337] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit20  (.D(net62),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[191] ),
    .Q_N(\ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit21  (.D(net63),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[227] ),
    .Q_N(\ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit22  (.D(net64),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[225] ),
    .Q_N(\ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit23  (.D(net65),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[224] ),
    .Q_N(\ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit24  (.D(net66),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[223] ),
    .Q_N(\ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit25  (.D(net67),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[269] ),
    .Q_N(\ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit26  (.D(net68),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[266] ),
    .Q_N(\ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit27  (.D(net69),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[593] ),
    .Q_N(\ConfigBits_N[593] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit28  (.D(net70),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[587] ),
    .Q_N(\ConfigBits_N[587] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit29  (.D(net71),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[612] ),
    .Q_N(\ConfigBits_N[612] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit3  (.D(net75),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[333] ),
    .Q_N(\ConfigBits_N[333] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit30  (.D(net73),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[586] ),
    .Q_N(\ConfigBits_N[586] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit31  (.D(net74),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[594] ),
    .Q_N(\ConfigBits_N[594] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit4  (.D(net76),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[342] ),
    .Q_N(\ConfigBits_N[342] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit5  (.D(net77),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[362] ),
    .Q_N(\ConfigBits_N[362] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit6  (.D(net78),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[372] ),
    .Q_N(\ConfigBits_N[372] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit7  (.D(net79),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[401] ),
    .Q_N(\ConfigBits_N[401] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit8  (.D(net80),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[408] ),
    .Q_N(\ConfigBits_N[408] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame12_bit9  (.D(net81),
    .GATE(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[392] ),
    .Q_N(\ConfigBits_N[392] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit0  (.D(net50),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[302] ),
    .Q_N(\ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit1  (.D(net61),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[326] ),
    .Q_N(\ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit10  (.D(net51),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[406] ),
    .Q_N(\ConfigBits_N[406] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit11  (.D(net52),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[393] ),
    .Q_N(\ConfigBits_N[393] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit12  (.D(net53),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[26] ),
    .Q_N(\ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit13  (.D(net54),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[55] ),
    .Q_N(\ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit14  (.D(net55),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[125] ),
    .Q_N(\ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit15  (.D(net56),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[124] ),
    .Q_N(\ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit16  (.D(net57),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[145] ),
    .Q_N(\ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit17  (.D(net58),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[142] ),
    .Q_N(\ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit18  (.D(net59),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[141] ),
    .Q_N(\ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit19  (.D(net60),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[149] ),
    .Q_N(\ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit2  (.D(net72),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[321] ),
    .Q_N(\ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit20  (.D(net62),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[190] ),
    .Q_N(\ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit21  (.D(net63),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[189] ),
    .Q_N(\ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit22  (.D(net64),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[226] ),
    .Q_N(\ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit23  (.D(net65),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[267] ),
    .Q_N(\ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit24  (.D(net66),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[288] ),
    .Q_N(\ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit25  (.D(net67),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[287] ),
    .Q_N(\ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit26  (.D(net68),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[277] ),
    .Q_N(\ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit27  (.D(net69),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[276] ),
    .Q_N(\ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit28  (.D(net70),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[592] ),
    .Q_N(\ConfigBits_N[592] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit29  (.D(net71),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[613] ),
    .Q_N(\ConfigBits_N[613] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit3  (.D(net75),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[313] ),
    .Q_N(\ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit30  (.D(net73),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[611] ),
    .Q_N(\ConfigBits_N[611] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit31  (.D(net74),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[595] ),
    .Q_N(\ConfigBits_N[595] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit4  (.D(net76),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[306] ),
    .Q_N(\ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit5  (.D(net77),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[343] ),
    .Q_N(\ConfigBits_N[343] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit6  (.D(net78),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[365] ),
    .Q_N(\ConfigBits_N[365] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit7  (.D(net79),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[373] ),
    .Q_N(\ConfigBits_N[373] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit8  (.D(net80),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[409] ),
    .Q_N(\ConfigBits_N[409] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame13_bit9  (.D(net81),
    .GATE(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[407] ),
    .Q_N(\ConfigBits_N[407] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit0  (.D(net50),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[305] ),
    .Q_N(\ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit1  (.D(net61),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[303] ),
    .Q_N(\ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit10  (.D(net51),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[357] ),
    .Q_N(\ConfigBits_N[357] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit11  (.D(net52),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[356] ),
    .Q_N(\ConfigBits_N[356] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit12  (.D(net53),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[344] ),
    .Q_N(\ConfigBits_N[344] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit13  (.D(net54),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[364] ),
    .Q_N(\ConfigBits_N[364] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit14  (.D(net55),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[399] ),
    .Q_N(\ConfigBits_N[399] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit15  (.D(net56),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[7] ),
    .Q_N(\ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit16  (.D(net57),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[65] ),
    .Q_N(\ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit17  (.D(net58),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[62] ),
    .Q_N(\ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit18  (.D(net59),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[100] ),
    .Q_N(\ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit19  (.D(net60),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[107] ),
    .Q_N(\ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit2  (.D(net72),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[323] ),
    .Q_N(\ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit20  (.D(net62),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[130] ),
    .Q_N(\ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit21  (.D(net63),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[144] ),
    .Q_N(\ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit22  (.D(net64),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[147] ),
    .Q_N(\ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit23  (.D(net65),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[192] ),
    .Q_N(\ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit24  (.D(net66),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[183] ),
    .Q_N(\ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit25  (.D(net67),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[182] ),
    .Q_N(\ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit26  (.D(net68),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[228] ),
    .Q_N(\ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit27  (.D(net69),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[272] ),
    .Q_N(\ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit28  (.D(net70),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[293] ),
    .Q_N(\ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit29  (.D(net71),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[291] ),
    .Q_N(\ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit3  (.D(net75),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[320] ),
    .Q_N(\ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit30  (.D(net73),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[278] ),
    .Q_N(\ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit31  (.D(net74),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[614] ),
    .Q_N(\ConfigBits_N[614] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit4  (.D(net76),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[316] ),
    .Q_N(\ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit5  (.D(net77),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[312] ),
    .Q_N(\ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit6  (.D(net78),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[310] ),
    .Q_N(\ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit7  (.D(net79),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[308] ),
    .Q_N(\ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit8  (.D(net80),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[307] ),
    .Q_N(\ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame14_bit9  (.D(net81),
    .GATE(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[334] ),
    .Q_N(\ConfigBits_N[334] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit0  (.D(net50),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[301] ),
    .Q_N(\ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit1  (.D(net61),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[300] ),
    .Q_N(\ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit10  (.D(net51),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[25] ),
    .Q_N(\ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit11  (.D(net52),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[24] ),
    .Q_N(\ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit12  (.D(net53),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[23] ),
    .Q_N(\ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit13  (.D(net54),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[68] ),
    .Q_N(\ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit14  (.D(net55),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[64] ),
    .Q_N(\ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit15  (.D(net56),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[61] ),
    .Q_N(\ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit16  (.D(net57),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[81] ),
    .Q_N(\ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit17  (.D(net58),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[102] ),
    .Q_N(\ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit18  (.D(net59),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[101] ),
    .Q_N(\ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit19  (.D(net60),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[99] ),
    .Q_N(\ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit2  (.D(net72),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[319] ),
    .Q_N(\ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit20  (.D(net62),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[95] ),
    .Q_N(\ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit21  (.D(net63),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[74] ),
    .Q_N(\ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit22  (.D(net64),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[112] ),
    .Q_N(\ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit23  (.D(net65),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[110] ),
    .Q_N(\ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit24  (.D(net66),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[108] ),
    .Q_N(\ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit25  (.D(net67),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[132] ),
    .Q_N(\ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit26  (.D(net68),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[273] ),
    .Q_N(\ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit27  (.D(net69),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[268] ),
    .Q_N(\ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit28  (.D(net70),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[289] ),
    .Q_N(\ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit29  (.D(net71),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[282] ),
    .Q_N(\ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit3  (.D(net75),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[317] ),
    .Q_N(\ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit30  (.D(net73),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[279] ),
    .Q_N(\ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit31  (.D(net74),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[275] ),
    .Q_N(\ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit4  (.D(net76),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[298] ),
    .Q_N(\ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit5  (.D(net77),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[309] ),
    .Q_N(\ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit6  (.D(net78),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[3] ),
    .Q_N(\ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit7  (.D(net79),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[16] ),
    .Q_N(\ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit8  (.D(net80),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[38] ),
    .Q_N(\ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame15_bit9  (.D(net81),
    .GATE(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[36] ),
    .Q_N(\ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit0  (.D(net50),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[335] ),
    .Q_N(\ConfigBits_N[335] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit1  (.D(net61),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[345] ),
    .Q_N(\ConfigBits_N[345] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit10  (.D(net51),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[19] ),
    .Q_N(\ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit11  (.D(net52),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[18] ),
    .Q_N(\ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit12  (.D(net53),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[71] ),
    .Q_N(\ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit13  (.D(net54),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[43] ),
    .Q_N(\ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit14  (.D(net55),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[69] ),
    .Q_N(\ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit15  (.D(net56),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[66] ),
    .Q_N(\ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit16  (.D(net57),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[42] ),
    .Q_N(\ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit17  (.D(net58),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[58] ),
    .Q_N(\ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit18  (.D(net59),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[57] ),
    .Q_N(\ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit19  (.D(net60),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[40] ),
    .Q_N(\ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit2  (.D(net72),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[6] ),
    .Q_N(\ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit20  (.D(net62),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[80] ),
    .Q_N(\ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit21  (.D(net63),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[76] ),
    .Q_N(\ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit22  (.D(net64),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[103] ),
    .Q_N(\ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit23  (.D(net65),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[98] ),
    .Q_N(\ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit24  (.D(net66),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[96] ),
    .Q_N(\ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit25  (.D(net67),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[93] ),
    .Q_N(\ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit26  (.D(net68),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[72] ),
    .Q_N(\ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit27  (.D(net69),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[111] ),
    .Q_N(\ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit28  (.D(net70),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[109] ),
    .Q_N(\ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit29  (.D(net71),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[104] ),
    .Q_N(\ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit3  (.D(net75),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[17] ),
    .Q_N(\ConfigBits_N[17] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit30  (.D(net73),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[283] ),
    .Q_N(\ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit31  (.D(net74),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[274] ),
    .Q_N(\ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit4  (.D(net76),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[35] ),
    .Q_N(\ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit5  (.D(net77),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[32] ),
    .Q_N(\ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit6  (.D(net78),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[31] ),
    .Q_N(\ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit7  (.D(net79),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[29] ),
    .Q_N(\ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit8  (.D(net80),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[27] ),
    .Q_N(\ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame16_bit9  (.D(net81),
    .GATE(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[20] ),
    .Q_N(\ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit0  (.D(net50),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[304] ),
    .Q_N(\ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit1  (.D(net61),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[299] ),
    .Q_N(\ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit10  (.D(net51),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[22] ),
    .Q_N(\ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit11  (.D(net52),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[21] ),
    .Q_N(\ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit12  (.D(net53),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[48] ),
    .Q_N(\ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit13  (.D(net54),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[45] ),
    .Q_N(\ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit14  (.D(net55),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[44] ),
    .Q_N(\ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit15  (.D(net56),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[60] ),
    .Q_N(\ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit16  (.D(net57),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[59] ),
    .Q_N(\ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit17  (.D(net58),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[56] ),
    .Q_N(\ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit18  (.D(net59),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[50] ),
    .Q_N(\ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit19  (.D(net60),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[41] ),
    .Q_N(\ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit2  (.D(net72),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[325] ),
    .Q_N(\ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit20  (.D(net62),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[79] ),
    .Q_N(\ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit21  (.D(net63),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[78] ),
    .Q_N(\ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit22  (.D(net64),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[77] ),
    .Q_N(\ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit23  (.D(net65),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[97] ),
    .Q_N(\ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit24  (.D(net66),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[92] ),
    .Q_N(\ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit25  (.D(net67),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[83] ),
    .Q_N(\ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit26  (.D(net68),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[82] ),
    .Q_N(\ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit27  (.D(net69),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[113] ),
    .Q_N(\ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit28  (.D(net70),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[106] ),
    .Q_N(\ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit29  (.D(net71),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[105] ),
    .Q_N(\ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit3  (.D(net75),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[5] ),
    .Q_N(\ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit30  (.D(net73),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[295] ),
    .Q_N(\ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit31  (.D(net74),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[285] ),
    .Q_N(\ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit4  (.D(net76),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[4] ),
    .Q_N(\ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit5  (.D(net77),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[2] ),
    .Q_N(\ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit6  (.D(net78),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[1] ),
    .Q_N(\ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit7  (.D(net79),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[0] ),
    .Q_N(\ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit8  (.D(net80),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[34] ),
    .Q_N(\ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame17_bit9  (.D(net81),
    .GATE(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[33] ),
    .Q_N(\ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit0  (.D(net50),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[324] ),
    .Q_N(\ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit1  (.D(net61),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[315] ),
    .Q_N(\ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit10  (.D(net51),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[9] ),
    .Q_N(\ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit11  (.D(net52),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[8] ),
    .Q_N(\ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit12  (.D(net53),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[49] ),
    .Q_N(\ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit13  (.D(net54),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[47] ),
    .Q_N(\ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit14  (.D(net55),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[46] ),
    .Q_N(\ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit15  (.D(net56),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[54] ),
    .Q_N(\ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit16  (.D(net57),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[53] ),
    .Q_N(\ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit17  (.D(net58),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[52] ),
    .Q_N(\ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit18  (.D(net59),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[51] ),
    .Q_N(\ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit19  (.D(net60),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[75] ),
    .Q_N(\ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit2  (.D(net72),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[314] ),
    .Q_N(\ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit20  (.D(net62),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[94] ),
    .Q_N(\ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit21  (.D(net63),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[91] ),
    .Q_N(\ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit22  (.D(net64),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[90] ),
    .Q_N(\ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit23  (.D(net65),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[89] ),
    .Q_N(\ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit24  (.D(net66),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[88] ),
    .Q_N(\ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit25  (.D(net67),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[87] ),
    .Q_N(\ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit26  (.D(net68),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[86] ),
    .Q_N(\ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit27  (.D(net69),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[85] ),
    .Q_N(\ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit28  (.D(net70),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[84] ),
    .Q_N(\ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit29  (.D(net71),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[73] ),
    .Q_N(\ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit3  (.D(net75),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[15] ),
    .Q_N(\ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit30  (.D(net73),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[294] ),
    .Q_N(\ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit31  (.D(net74),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[284] ),
    .Q_N(\ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit4  (.D(net76),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[14] ),
    .Q_N(\ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit5  (.D(net77),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[13] ),
    .Q_N(\ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit6  (.D(net78),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[12] ),
    .Q_N(\ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit7  (.D(net79),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[11] ),
    .Q_N(\ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit8  (.D(net80),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[37] ),
    .Q_N(\ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame18_bit9  (.D(net81),
    .GATE(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[10] ),
    .Q_N(\ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit10  (.D(net51),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[467] ),
    .Q_N(\ConfigBits_N[467] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit11  (.D(net52),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[575] ),
    .Q_N(\ConfigBits_N[575] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit12  (.D(net53),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[574] ),
    .Q_N(\ConfigBits_N[574] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit13  (.D(net54),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[567] ),
    .Q_N(\ConfigBits_N[567] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit14  (.D(net55),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[566] ),
    .Q_N(\ConfigBits_N[566] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit15  (.D(net56),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[562] ),
    .Q_N(\ConfigBits_N[562] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit16  (.D(net57),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[156] ),
    .Q_N(\ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit17  (.D(net58),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[155] ),
    .Q_N(\ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit18  (.D(net59),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[154] ),
    .Q_N(\ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit19  (.D(net60),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[239] ),
    .Q_N(\ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit2  (.D(net72),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[396] ),
    .Q_N(\ConfigBits_N[396] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit20  (.D(net62),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[238] ),
    .Q_N(\ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit21  (.D(net63),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[258] ),
    .Q_N(\ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit22  (.D(net64),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[254] ),
    .Q_N(\ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit23  (.D(net65),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[253] ),
    .Q_N(\ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit24  (.D(net66),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[252] ),
    .Q_N(\ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit25  (.D(net67),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[246] ),
    .Q_N(\ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit3  (.D(net75),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[412] ),
    .Q_N(\ConfigBits_N[412] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit4  (.D(net76),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[405] ),
    .Q_N(\ConfigBits_N[405] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit5  (.D(net77),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[404] ),
    .Q_N(\ConfigBits_N[404] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit6  (.D(net78),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[479] ),
    .Q_N(\ConfigBits_N[479] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit7  (.D(net79),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[478] ),
    .Q_N(\ConfigBits_N[478] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit8  (.D(net80),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[471] ),
    .Q_N(\ConfigBits_N[471] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame19_bit9  (.D(net81),
    .GATE(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[470] ),
    .Q_N(\ConfigBits_N[470] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit10  (.D(net51),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[526] ),
    .Q_N(\ConfigBits_N[526] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit11  (.D(net52),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[543] ),
    .Q_N(\ConfigBits_N[543] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit12  (.D(net53),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[542] ),
    .Q_N(\ConfigBits_N[542] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit13  (.D(net54),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[537] ),
    .Q_N(\ConfigBits_N[537] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit14  (.D(net55),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[534] ),
    .Q_N(\ConfigBits_N[534] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit15  (.D(net56),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[530] ),
    .Q_N(\ConfigBits_N[530] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit16  (.D(net57),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[560] ),
    .Q_N(\ConfigBits_N[560] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit17  (.D(net58),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[559] ),
    .Q_N(\ConfigBits_N[559] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit18  (.D(net59),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[578] ),
    .Q_N(\ConfigBits_N[578] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit19  (.D(net60),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[573] ),
    .Q_N(\ConfigBits_N[573] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit2  (.D(net72),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[388] ),
    .Q_N(\ConfigBits_N[388] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit20  (.D(net62),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[572] ),
    .Q_N(\ConfigBits_N[572] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit21  (.D(net63),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[571] ),
    .Q_N(\ConfigBits_N[571] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit22  (.D(net64),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[570] ),
    .Q_N(\ConfigBits_N[570] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit23  (.D(net65),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[569] ),
    .Q_N(\ConfigBits_N[569] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit24  (.D(net66),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[565] ),
    .Q_N(\ConfigBits_N[565] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit25  (.D(net67),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[563] ),
    .Q_N(\ConfigBits_N[563] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit26  (.D(net68),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[262] ),
    .Q_N(\ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit27  (.D(net69),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[260] ),
    .Q_N(\ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit28  (.D(net70),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[256] ),
    .Q_N(\ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit29  (.D(net71),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[255] ),
    .Q_N(\ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit3  (.D(net75),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[386] ),
    .Q_N(\ConfigBits_N[386] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit30  (.D(net73),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[250] ),
    .Q_N(\ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit31  (.D(net74),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[249] ),
    .Q_N(\ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit4  (.D(net76),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[422] ),
    .Q_N(\ConfigBits_N[422] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit5  (.D(net77),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[463] ),
    .Q_N(\ConfigBits_N[463] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit7  (.D(net79),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[480] ),
    .Q_N(\ConfigBits_N[480] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit8  (.D(net80),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[504] ),
    .Q_N(\ConfigBits_N[504] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame1_bit9  (.D(net81),
    .GATE(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[527] ),
    .Q_N(\ConfigBits_N[527] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit1  (.D(net61),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[348] ),
    .Q_N(\ConfigBits_N[348] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit10  (.D(net51),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[483] ),
    .Q_N(\ConfigBits_N[483] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit11  (.D(net52),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[475] ),
    .Q_N(\ConfigBits_N[475] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit12  (.D(net53),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[474] ),
    .Q_N(\ConfigBits_N[474] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit13  (.D(net54),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[494] ),
    .Q_N(\ConfigBits_N[494] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit14  (.D(net55),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[503] ),
    .Q_N(\ConfigBits_N[503] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit15  (.D(net56),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[499] ),
    .Q_N(\ConfigBits_N[499] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit16  (.D(net57),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[498] ),
    .Q_N(\ConfigBits_N[498] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit17  (.D(net58),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[529] ),
    .Q_N(\ConfigBits_N[529] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit18  (.D(net59),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[528] ),
    .Q_N(\ConfigBits_N[528] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit19  (.D(net60),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[544] ),
    .Q_N(\ConfigBits_N[544] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit20  (.D(net62),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[536] ),
    .Q_N(\ConfigBits_N[536] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit21  (.D(net63),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[535] ),
    .Q_N(\ConfigBits_N[535] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit22  (.D(net64),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[531] ),
    .Q_N(\ConfigBits_N[531] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit23  (.D(net65),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[561] ),
    .Q_N(\ConfigBits_N[561] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit24  (.D(net66),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[564] ),
    .Q_N(\ConfigBits_N[564] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit25  (.D(net67),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[167] ),
    .Q_N(\ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit26  (.D(net68),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[163] ),
    .Q_N(\ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit27  (.D(net69),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[257] ),
    .Q_N(\ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit28  (.D(net70),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[251] ),
    .Q_N(\ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit30  (.D(net73),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[265] ),
    .Q_N(\ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit31  (.D(net74),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[264] ),
    .Q_N(\ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit4  (.D(net76),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[366] ),
    .Q_N(\ConfigBits_N[366] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit5  (.D(net77),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[374] ),
    .Q_N(\ConfigBits_N[374] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit6  (.D(net78),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[423] ),
    .Q_N(\ConfigBits_N[423] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit7  (.D(net79),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[439] ),
    .Q_N(\ConfigBits_N[439] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit8  (.D(net80),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[464] ),
    .Q_N(\ConfigBits_N[464] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame2_bit9  (.D(net81),
    .GATE(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[461] ),
    .Q_N(\ConfigBits_N[461] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit1  (.D(net61),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[336] ),
    .Q_N(\ConfigBits_N[336] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit10  (.D(net51),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[438] ),
    .Q_N(\ConfigBits_N[438] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit11  (.D(net52),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[465] ),
    .Q_N(\ConfigBits_N[465] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit12  (.D(net53),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[477] ),
    .Q_N(\ConfigBits_N[477] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit13  (.D(net54),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[476] ),
    .Q_N(\ConfigBits_N[476] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit14  (.D(net55),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[497] ),
    .Q_N(\ConfigBits_N[497] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit15  (.D(net56),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[496] ),
    .Q_N(\ConfigBits_N[496] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit16  (.D(net57),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[495] ),
    .Q_N(\ConfigBits_N[495] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit17  (.D(net58),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[491] ),
    .Q_N(\ConfigBits_N[491] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit18  (.D(net59),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[505] ),
    .Q_N(\ConfigBits_N[505] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit19  (.D(net60),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[501] ),
    .Q_N(\ConfigBits_N[501] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit2  (.D(net72),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[353] ),
    .Q_N(\ConfigBits_N[353] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit20  (.D(net62),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[500] ),
    .Q_N(\ConfigBits_N[500] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit21  (.D(net63),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[547] ),
    .Q_N(\ConfigBits_N[547] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit22  (.D(net64),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[546] ),
    .Q_N(\ConfigBits_N[546] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit23  (.D(net65),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[545] ),
    .Q_N(\ConfigBits_N[545] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit24  (.D(net66),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[533] ),
    .Q_N(\ConfigBits_N[533] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit25  (.D(net67),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[67] ),
    .Q_N(\ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit26  (.D(net68),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[166] ),
    .Q_N(\ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit27  (.D(net69),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[164] ),
    .Q_N(\ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit28  (.D(net70),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[162] ),
    .Q_N(\ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit29  (.D(net71),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[153] ),
    .Q_N(\ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit3  (.D(net75),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[349] ),
    .Q_N(\ConfigBits_N[349] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit30  (.D(net73),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[186] ),
    .Q_N(\ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit31  (.D(net74),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[168] ),
    .Q_N(\ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit4  (.D(net76),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[367] ),
    .Q_N(\ConfigBits_N[367] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit5  (.D(net77),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[431] ),
    .Q_N(\ConfigBits_N[431] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit6  (.D(net78),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[430] ),
    .Q_N(\ConfigBits_N[430] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit7  (.D(net79),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[451] ),
    .Q_N(\ConfigBits_N[451] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit8  (.D(net80),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[450] ),
    .Q_N(\ConfigBits_N[450] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame3_bit9  (.D(net81),
    .GATE(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[446] ),
    .Q_N(\ConfigBits_N[446] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit0  (.D(net50),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[358] ),
    .Q_N(\ConfigBits_N[358] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit1  (.D(net61),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[352] ),
    .Q_N(\ConfigBits_N[352] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit10  (.D(net51),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[486] ),
    .Q_N(\ConfigBits_N[486] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit11  (.D(net52),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[482] ),
    .Q_N(\ConfigBits_N[482] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit12  (.D(net53),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[469] ),
    .Q_N(\ConfigBits_N[469] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit13  (.D(net54),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[468] ),
    .Q_N(\ConfigBits_N[468] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit14  (.D(net55),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[466] ),
    .Q_N(\ConfigBits_N[466] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit15  (.D(net56),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[517] ),
    .Q_N(\ConfigBits_N[517] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit16  (.D(net57),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[515] ),
    .Q_N(\ConfigBits_N[515] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit17  (.D(net58),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[514] ),
    .Q_N(\ConfigBits_N[514] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit18  (.D(net59),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[509] ),
    .Q_N(\ConfigBits_N[509] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit19  (.D(net60),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[489] ),
    .Q_N(\ConfigBits_N[489] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit2  (.D(net72),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[363] ),
    .Q_N(\ConfigBits_N[363] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit20  (.D(net62),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[550] ),
    .Q_N(\ConfigBits_N[550] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit21  (.D(net63),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[549] ),
    .Q_N(\ConfigBits_N[549] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit22  (.D(net64),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[532] ),
    .Q_N(\ConfigBits_N[532] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit23  (.D(net65),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[165] ),
    .Q_N(\ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit24  (.D(net66),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[152] ),
    .Q_N(\ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit25  (.D(net67),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[176] ),
    .Q_N(\ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit26  (.D(net68),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[184] ),
    .Q_N(\ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit27  (.D(net69),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[179] ),
    .Q_N(\ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit28  (.D(net70),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[169] ),
    .Q_N(\ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit29  (.D(net71),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[203] ),
    .Q_N(\ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit3  (.D(net75),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[375] ),
    .Q_N(\ConfigBits_N[375] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit30  (.D(net73),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[216] ),
    .Q_N(\ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit31  (.D(net74),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[604] ),
    .Q_N(\ConfigBits_N[604] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit4  (.D(net76),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[371] ),
    .Q_N(\ConfigBits_N[371] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit5  (.D(net77),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[370] ),
    .Q_N(\ConfigBits_N[370] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit6  (.D(net78),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[428] ),
    .Q_N(\ConfigBits_N[428] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit7  (.D(net79),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[455] ),
    .Q_N(\ConfigBits_N[455] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit8  (.D(net80),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[452] ),
    .Q_N(\ConfigBits_N[452] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame4_bit9  (.D(net81),
    .GATE(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[447] ),
    .Q_N(\ConfigBits_N[447] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit0  (.D(net50),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[359] ),
    .Q_N(\ConfigBits_N[359] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit1  (.D(net61),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[346] ),
    .Q_N(\ConfigBits_N[346] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit10  (.D(net51),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[437] ),
    .Q_N(\ConfigBits_N[437] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit11  (.D(net52),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[436] ),
    .Q_N(\ConfigBits_N[436] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit12  (.D(net53),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[458] ),
    .Q_N(\ConfigBits_N[458] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit13  (.D(net54),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[457] ),
    .Q_N(\ConfigBits_N[457] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit14  (.D(net55),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[516] ),
    .Q_N(\ConfigBits_N[516] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit15  (.D(net56),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[511] ),
    .Q_N(\ConfigBits_N[511] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit16  (.D(net57),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[510] ),
    .Q_N(\ConfigBits_N[510] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit17  (.D(net58),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[506] ),
    .Q_N(\ConfigBits_N[506] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit18  (.D(net59),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[551] ),
    .Q_N(\ConfigBits_N[551] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit19  (.D(net60),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[548] ),
    .Q_N(\ConfigBits_N[548] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit2  (.D(net72),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[421] ),
    .Q_N(\ConfigBits_N[421] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit20  (.D(net62),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[126] ),
    .Q_N(\ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit21  (.D(net63),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[177] ),
    .Q_N(\ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit22  (.D(net64),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[175] ),
    .Q_N(\ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit23  (.D(net65),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[174] ),
    .Q_N(\ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit24  (.D(net66),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[173] ),
    .Q_N(\ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit25  (.D(net67),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[185] ),
    .Q_N(\ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit26  (.D(net68),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[178] ),
    .Q_N(\ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit27  (.D(net69),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[205] ),
    .Q_N(\ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit28  (.D(net70),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[229] ),
    .Q_N(\ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit29  (.D(net71),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[202] ),
    .Q_N(\ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit3  (.D(net75),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[429] ),
    .Q_N(\ConfigBits_N[429] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit30  (.D(net73),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[210] ),
    .Q_N(\ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit31  (.D(net74),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[589] ),
    .Q_N(\ConfigBits_N[589] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit4  (.D(net76),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[454] ),
    .Q_N(\ConfigBits_N[454] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit5  (.D(net77),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[453] ),
    .Q_N(\ConfigBits_N[453] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit6  (.D(net78),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[448] ),
    .Q_N(\ConfigBits_N[448] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit7  (.D(net79),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[444] ),
    .Q_N(\ConfigBits_N[444] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit8  (.D(net80),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[441] ),
    .Q_N(\ConfigBits_N[441] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame5_bit9  (.D(net81),
    .GATE(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[440] ),
    .Q_N(\ConfigBits_N[440] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit0  (.D(net50),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[311] ),
    .Q_N(\ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit1  (.D(net61),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[347] ),
    .Q_N(\ConfigBits_N[347] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit10  (.D(net51),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[484] ),
    .Q_N(\ConfigBits_N[484] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit11  (.D(net52),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[456] ),
    .Q_N(\ConfigBits_N[456] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit12  (.D(net53),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[492] ),
    .Q_N(\ConfigBits_N[492] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit13  (.D(net54),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[513] ),
    .Q_N(\ConfigBits_N[513] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit14  (.D(net55),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[490] ),
    .Q_N(\ConfigBits_N[490] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit15  (.D(net56),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[507] ),
    .Q_N(\ConfigBits_N[507] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit16  (.D(net57),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[553] ),
    .Q_N(\ConfigBits_N[553] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit17  (.D(net58),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[30] ),
    .Q_N(\ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit18  (.D(net59),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[70] ),
    .Q_N(\ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit19  (.D(net60),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[119] ),
    .Q_N(\ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit2  (.D(net72),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[420] ),
    .Q_N(\ConfigBits_N[420] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit20  (.D(net62),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[170] ),
    .Q_N(\ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit21  (.D(net63),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[181] ),
    .Q_N(\ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit22  (.D(net64),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[208] ),
    .Q_N(\ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit23  (.D(net65),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[206] ),
    .Q_N(\ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit24  (.D(net66),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[204] ),
    .Q_N(\ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit25  (.D(net67),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[231] ),
    .Q_N(\ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit26  (.D(net68),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[214] ),
    .Q_N(\ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit27  (.D(net69),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[213] ),
    .Q_N(\ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit28  (.D(net70),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[212] ),
    .Q_N(\ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit29  (.D(net71),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[211] ),
    .Q_N(\ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit3  (.D(net75),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[433] ),
    .Q_N(\ConfigBits_N[433] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit30  (.D(net73),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[606] ),
    .Q_N(\ConfigBits_N[606] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit31  (.D(net74),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[605] ),
    .Q_N(\ConfigBits_N[605] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit4  (.D(net76),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[449] ),
    .Q_N(\ConfigBits_N[449] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit5  (.D(net77),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[425] ),
    .Q_N(\ConfigBits_N[425] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit6  (.D(net78),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[424] ),
    .Q_N(\ConfigBits_N[424] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit7  (.D(net79),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[487] ),
    .Q_N(\ConfigBits_N[487] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit8  (.D(net80),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[459] ),
    .Q_N(\ConfigBits_N[459] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame6_bit9  (.D(net81),
    .GATE(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[485] ),
    .Q_N(\ConfigBits_N[485] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit0  (.D(net50),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[340] ),
    .Q_N(\ConfigBits_N[340] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit1  (.D(net61),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[385] ),
    .Q_N(\ConfigBits_N[385] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit10  (.D(net51),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[512] ),
    .Q_N(\ConfigBits_N[512] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit11  (.D(net52),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[508] ),
    .Q_N(\ConfigBits_N[508] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit12  (.D(net53),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[488] ),
    .Q_N(\ConfigBits_N[488] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit13  (.D(net54),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[540] ),
    .Q_N(\ConfigBits_N[540] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit14  (.D(net55),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[522] ),
    .Q_N(\ConfigBits_N[522] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit15  (.D(net56),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[582] ),
    .Q_N(\ConfigBits_N[582] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit16  (.D(net57),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[555] ),
    .Q_N(\ConfigBits_N[555] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit17  (.D(net58),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[552] ),
    .Q_N(\ConfigBits_N[552] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit18  (.D(net59),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[121] ),
    .Q_N(\ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit19  (.D(net60),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[160] ),
    .Q_N(\ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit2  (.D(net72),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[415] ),
    .Q_N(\ConfigBits_N[415] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit20  (.D(net62),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[146] ),
    .Q_N(\ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit21  (.D(net63),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[172] ),
    .Q_N(\ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit22  (.D(net64),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[171] ),
    .Q_N(\ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit23  (.D(net65),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[180] ),
    .Q_N(\ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit24  (.D(net66),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[217] ),
    .Q_N(\ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit25  (.D(net67),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[236] ),
    .Q_N(\ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit26  (.D(net68),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[280] ),
    .Q_N(\ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit27  (.D(net69),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[590] ),
    .Q_N(\ConfigBits_N[590] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit28  (.D(net70),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[588] ),
    .Q_N(\ConfigBits_N[588] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit29  (.D(net71),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[609] ),
    .Q_N(\ConfigBits_N[609] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit3  (.D(net75),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[402] ),
    .Q_N(\ConfigBits_N[402] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit30  (.D(net73),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[608] ),
    .Q_N(\ConfigBits_N[608] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit31  (.D(net74),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[596] ),
    .Q_N(\ConfigBits_N[596] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit4  (.D(net76),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[442] ),
    .Q_N(\ConfigBits_N[442] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit5  (.D(net77),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[435] ),
    .Q_N(\ConfigBits_N[435] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit6  (.D(net78),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[434] ),
    .Q_N(\ConfigBits_N[434] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit7  (.D(net79),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[460] ),
    .Q_N(\ConfigBits_N[460] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit8  (.D(net80),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[493] ),
    .Q_N(\ConfigBits_N[493] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame7_bit9  (.D(net81),
    .GATE(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[519] ),
    .Q_N(\ConfigBits_N[519] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit0  (.D(net50),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[351] ),
    .Q_N(\ConfigBits_N[351] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit1  (.D(net61),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[329] ),
    .Q_N(\ConfigBits_N[329] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit10  (.D(net51),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[538] ),
    .Q_N(\ConfigBits_N[538] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit11  (.D(net52),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[520] ),
    .Q_N(\ConfigBits_N[520] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit12  (.D(net53),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[580] ),
    .Q_N(\ConfigBits_N[580] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit13  (.D(net54),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[554] ),
    .Q_N(\ConfigBits_N[554] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit14  (.D(net55),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[129] ),
    .Q_N(\ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit15  (.D(net56),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[161] ),
    .Q_N(\ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit16  (.D(net57),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[137] ),
    .Q_N(\ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit17  (.D(net58),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[194] ),
    .Q_N(\ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit18  (.D(net59),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[193] ),
    .Q_N(\ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit19  (.D(net60),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[209] ),
    .Q_N(\ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit2  (.D(net72),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[369] ),
    .Q_N(\ConfigBits_N[369] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit20  (.D(net62),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[207] ),
    .Q_N(\ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit21  (.D(net63),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[230] ),
    .Q_N(\ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit22  (.D(net64),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[219] ),
    .Q_N(\ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit23  (.D(net65),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[215] ),
    .Q_N(\ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit24  (.D(net66),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[235] ),
    .Q_N(\ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit25  (.D(net67),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[244] ),
    .Q_N(\ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit26  (.D(net68),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[290] ),
    .Q_N(\ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit27  (.D(net69),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[286] ),
    .Q_N(\ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit28  (.D(net70),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[607] ),
    .Q_N(\ConfigBits_N[607] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit29  (.D(net71),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[600] ),
    .Q_N(\ConfigBits_N[600] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit3  (.D(net75),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[432] ),
    .Q_N(\ConfigBits_N[432] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit30  (.D(net73),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[598] ),
    .Q_N(\ConfigBits_N[598] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit31  (.D(net74),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[597] ),
    .Q_N(\ConfigBits_N[597] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit4  (.D(net76),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[427] ),
    .Q_N(\ConfigBits_N[427] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit5  (.D(net77),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[426] ),
    .Q_N(\ConfigBits_N[426] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit6  (.D(net78),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[443] ),
    .Q_N(\ConfigBits_N[443] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit7  (.D(net79),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[518] ),
    .Q_N(\ConfigBits_N[518] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit8  (.D(net80),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[523] ),
    .Q_N(\ConfigBits_N[523] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame8_bit9  (.D(net81),
    .GATE(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[539] ),
    .Q_N(\ConfigBits_N[539] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit0  (.D(net50),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[354] ),
    .Q_N(\ConfigBits_N[354] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit1  (.D(net61),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[350] ),
    .Q_N(\ConfigBits_N[350] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit10  (.D(net51),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[361] ),
    .Q_N(\ConfigBits_N[361] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit11  (.D(net52),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[419] ),
    .Q_N(\ConfigBits_N[419] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit12  (.D(net53),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[418] ),
    .Q_N(\ConfigBits_N[418] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit13  (.D(net54),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[414] ),
    .Q_N(\ConfigBits_N[414] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit14  (.D(net55),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[445] ),
    .Q_N(\ConfigBits_N[445] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit15  (.D(net56),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[525] ),
    .Q_N(\ConfigBits_N[525] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit16  (.D(net57),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[524] ),
    .Q_N(\ConfigBits_N[524] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit17  (.D(net58),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[541] ),
    .Q_N(\ConfigBits_N[541] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit18  (.D(net59),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[556] ),
    .Q_N(\ConfigBits_N[556] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit19  (.D(net60),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[583] ),
    .Q_N(\ConfigBits_N[583] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit2  (.D(net72),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[341] ),
    .Q_N(\ConfigBits_N[341] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit20  (.D(net62),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[579] ),
    .Q_N(\ConfigBits_N[579] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit21  (.D(net63),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[136] ),
    .Q_N(\ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit22  (.D(net64),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[197] ),
    .Q_N(\ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit23  (.D(net65),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[195] ),
    .Q_N(\ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit24  (.D(net66),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[218] ),
    .Q_N(\ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit25  (.D(net67),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[237] ),
    .Q_N(\ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit26  (.D(net68),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[245] ),
    .Q_N(\ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit27  (.D(net69),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[292] ),
    .Q_N(\ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit28  (.D(net70),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[281] ),
    .Q_N(\ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit29  (.D(net71),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[591] ),
    .Q_N(\ConfigBits_N[591] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit3  (.D(net75),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[328] ),
    .Q_N(\ConfigBits_N[328] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit30  (.D(net73),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[603] ),
    .Q_N(\ConfigBits_N[603] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit31  (.D(net74),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[599] ),
    .Q_N(\ConfigBits_N[599] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit4  (.D(net76),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[368] ),
    .Q_N(\ConfigBits_N[368] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit5  (.D(net77),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[384] ),
    .Q_N(\ConfigBits_N[384] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit6  (.D(net78),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[383] ),
    .Q_N(\ConfigBits_N[383] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit7  (.D(net79),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[382] ),
    .Q_N(\ConfigBits_N[382] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit8  (.D(net80),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[379] ),
    .Q_N(\ConfigBits_N[379] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_LUT4AB_ConfigMem/Inst_Frame9_bit9  (.D(net81),
    .GATE(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .Q(\ConfigBits[378] ),
    .Q_N(\ConfigBits_N[378] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_032_  (.A(LA_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(A));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_033_  (.A(LB_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(B));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_034_  (.A(LC_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(C));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_035_  (.A(LH_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_036_  (.A(LD_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(D));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_037_  (.A(LE_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_038_  (.A(\JE2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_039_  (.A(\JE2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net260));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_040_  (.A(\JE2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_041_  (.A(\JE2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_042_  (.A(\JE2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_043_  (.A(\JE2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net264));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_044_  (.A(\JE2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_045_  (.A(\JE2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_046_  (.A(net14),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_047_  (.A(net15),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_048_  (.A(net16),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_2 \Inst_LUT4AB_switch_matrix/_049_  (.A(net17),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_050_  (.A(net18),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_051_  (.A(net19),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_052_  (.A(net20),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_053_  (.A(net21),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_054_  (.A(LF_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(F));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_055_  (.A(LG_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(G));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_056_  (.A(LH_O),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(H));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_057_  (.A(net1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_058_  (.A(LA_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_059_  (.A(LB_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_060_  (.A(LC_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_061_  (.A(LD_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_062_  (.A(LE_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_063_  (.A(LF_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_Ci));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_064_  (.A(LG_Co),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_Ci));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_065_  (.A(\JN2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_066_  (.A(\JN2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net360));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_067_  (.A(\JN2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_068_  (.A(\JN2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_069_  (.A(\JN2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_070_  (.A(\JN2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_071_  (.A(\JN2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_072_  (.A(\JN2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_073_  (.A(net114),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_074_  (.A(net115),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_075_  (.A(net116),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_076_  (.A(net117),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_077_  (.A(net118),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_078_  (.A(net119),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_079_  (.A(net120),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_080_  (.A(net121),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_081_  (.A(\JS2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_082_  (.A(\JS2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_083_  (.A(\JS2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_084_  (.A(\JS2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_085_  (.A(\JS2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net415));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_086_  (.A(\JS2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net416));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_087_  (.A(\JS2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net417));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_088_  (.A(\JS2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_089_  (.A(net166),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_090_  (.A(net167),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_091_  (.A(net168),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net421));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_092_  (.A(net169),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_093_  (.A(net170),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_094_  (.A(net171),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_095_  (.A(net172),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_096_  (.A(net173),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_097_  (.A(\JW2BEG[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_098_  (.A(\JW2BEG[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_099_  (.A(\JW2BEG[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_100_  (.A(\JW2BEG[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_101_  (.A(\JW2BEG[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_102_  (.A(\JW2BEG[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net469));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_103_  (.A(\JW2BEG[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_104_  (.A(\JW2BEG[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_105_  (.A(net218),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net472));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_106_  (.A(net219),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_107_  (.A(net220),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_108_  (.A(net221),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_109_  (.A(net222),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net476));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_110_  (.A(net223),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_1 \Inst_LUT4AB_switch_matrix/_111_  (.A(net224),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net478));
 sky130_fd_sc_hd__buf_1 \Inst_LUT4AB_switch_matrix/_112_  (.A(net225),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net479));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst0  (.A0(net5),
    .A1(net209),
    .A2(LA_O),
    .A3(LB_O),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(LD_O),
    .A2(LE_O),
    .A3(LF_O),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst2  (.A0(LG_O),
    .A1(LH_O),
    .A2(M_AB),
    .A3(M_AH),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst3  (.A0(\J2MID_ABb_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2MID_EFb_BEG[1] ),
    .A3(\J2MID_GHb_BEG[1] ),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[204] ),
    .S1(\ConfigBits[205] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net276));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net208),
    .A2(LA_O),
    .A3(LB_O),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(LD_O),
    .A2(LE_O),
    .A3(LF_O),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst2  (.A0(LG_O),
    .A1(LH_O),
    .A2(M_AD),
    .A3(M_EF),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst3  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_CDa_BEG[2] ),
    .A2(\J2MID_EFa_BEG[2] ),
    .A3(\J2MID_GHa_BEG[2] ),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_E6BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[208] ),
    .S1(\ConfigBits[209] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net107),
    .A2(net129),
    .A3(net41),
    .S0(\ConfigBits[482] ),
    .S1(\ConfigBits[483] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst1  (.A0(net25),
    .A1(net159),
    .A2(net211),
    .A3(net229),
    .S0(\ConfigBits[482] ),
    .S1(\ConfigBits[483] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst2  (.A0(LB_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[482] ),
    .S1(\ConfigBits[483] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[482] ),
    .S1(\ConfigBits[483] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[484] ),
    .S1(\ConfigBits[485] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net130),
    .A3(net8),
    .S0(\ConfigBits[486] ),
    .S1(\ConfigBits[487] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst1  (.A0(net22),
    .A1(net160),
    .A2(net212),
    .A3(net247),
    .S0(\ConfigBits[486] ),
    .S1(\ConfigBits[487] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[486] ),
    .S1(\ConfigBits[487] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[486] ),
    .S1(\ConfigBits[487] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[488] ),
    .S1(\ConfigBits[489] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net131),
    .A3(net9),
    .S0(\ConfigBits[490] ),
    .S1(\ConfigBits[491] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst1  (.A0(net25),
    .A1(net161),
    .A2(net213),
    .A3(net229),
    .S0(\ConfigBits[490] ),
    .S1(\ConfigBits[491] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[490] ),
    .S1(\ConfigBits[491] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[490] ),
    .S1(\ConfigBits[491] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[492] ),
    .S1(\ConfigBits[493] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net110),
    .A2(net122),
    .A3(net10),
    .S0(\ConfigBits[494] ),
    .S1(\ConfigBits[495] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst1  (.A0(net22),
    .A1(net162),
    .A2(net214),
    .A3(net226),
    .S0(\ConfigBits[494] ),
    .S1(\ConfigBits[495] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LE_O),
    .S0(\ConfigBits[494] ),
    .S1(\ConfigBits[495] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[494] ),
    .S1(\ConfigBits[495] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[496] ),
    .S1(\ConfigBits[497] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[498] ),
    .S1(\ConfigBits[499] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net163),
    .A3(net207),
    .S0(\ConfigBits[498] ),
    .S1(\ConfigBits[499] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[498] ),
    .S1(\ConfigBits[499] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[498] ),
    .S1(\ConfigBits[499] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[500] ),
    .S1(\ConfigBits[501] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[502] ),
    .S1(\ConfigBits[503] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net164),
    .A3(net208),
    .S0(\ConfigBits[502] ),
    .S1(\ConfigBits[503] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[502] ),
    .S1(\ConfigBits[503] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[502] ),
    .S1(\ConfigBits[503] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[504] ),
    .S1(\ConfigBits[505] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\ConfigBits[506] ),
    .S1(\ConfigBits[507] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net165),
    .A3(net209),
    .S0(\ConfigBits[506] ),
    .S1(\ConfigBits[507] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[506] ),
    .S1(\ConfigBits[507] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[506] ),
    .S1(\ConfigBits[507] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[508] ),
    .S1(\ConfigBits[509] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net6),
    .S0(\ConfigBits[510] ),
    .S1(\ConfigBits[511] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net190),
    .A3(net238),
    .S0(\ConfigBits[510] ),
    .S1(\ConfigBits[511] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[510] ),
    .S1(\ConfigBits[511] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LG_O),
    .A3(M_AH),
    .S0(\ConfigBits[510] ),
    .S1(\ConfigBits[511] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JE2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[512] ),
    .S1(\ConfigBits[513] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JE2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst0  (.A0(net107),
    .A1(net129),
    .A2(net5),
    .A3(net7),
    .S0(\ConfigBits[450] ),
    .S1(\ConfigBits[451] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst1  (.A0(net25),
    .A1(net197),
    .A2(net211),
    .A3(net229),
    .S0(\ConfigBits[450] ),
    .S1(\ConfigBits[451] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst2  (.A0(LB_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[450] ),
    .S1(\ConfigBits[451] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[450] ),
    .S1(\ConfigBits[451] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[452] ),
    .S1(\ConfigBits[453] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst0  (.A0(net108),
    .A1(net130),
    .A2(net2),
    .A3(net8),
    .S0(\ConfigBits[454] ),
    .S1(\ConfigBits[455] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst1  (.A0(net22),
    .A1(net160),
    .A2(net212),
    .A3(net226),
    .S0(\ConfigBits[454] ),
    .S1(\ConfigBits[455] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[454] ),
    .S1(\ConfigBits[455] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[454] ),
    .S1(\ConfigBits[455] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[456] ),
    .S1(\ConfigBits[457] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst0  (.A0(net109),
    .A1(net131),
    .A2(net3),
    .A3(net9),
    .S0(\ConfigBits[458] ),
    .S1(\ConfigBits[459] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst1  (.A0(net25),
    .A1(net161),
    .A2(net213),
    .A3(net245),
    .S0(\ConfigBits[458] ),
    .S1(\ConfigBits[459] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[458] ),
    .S1(\ConfigBits[459] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[458] ),
    .S1(\ConfigBits[459] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[460] ),
    .S1(\ConfigBits[461] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst0  (.A0(net110),
    .A1(net122),
    .A2(net4),
    .A3(net10),
    .S0(\ConfigBits[462] ),
    .S1(\ConfigBits[463] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst1  (.A0(net22),
    .A1(net162),
    .A2(net214),
    .A3(net226),
    .S0(\ConfigBits[462] ),
    .S1(\ConfigBits[463] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LE_O),
    .S0(\ConfigBits[462] ),
    .S1(\ConfigBits[463] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[462] ),
    .S1(\ConfigBits[463] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[464] ),
    .S1(\ConfigBits[465] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[466] ),
    .S1(\ConfigBits[467] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net163),
    .A2(net207),
    .A3(net209),
    .S0(\ConfigBits[466] ),
    .S1(\ConfigBits[467] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[466] ),
    .S1(\ConfigBits[467] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[466] ),
    .S1(\ConfigBits[467] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[468] ),
    .S1(\ConfigBits[469] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[470] ),
    .S1(\ConfigBits[471] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst1  (.A0(net156),
    .A1(net164),
    .A2(net206),
    .A3(net208),
    .S0(\ConfigBits[470] ),
    .S1(\ConfigBits[471] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[470] ),
    .S1(\ConfigBits[471] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[470] ),
    .S1(\ConfigBits[471] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[472] ),
    .S1(\ConfigBits[473] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\ConfigBits[474] ),
    .S1(\ConfigBits[475] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst1  (.A0(net157),
    .A1(net165),
    .A2(net207),
    .A3(net209),
    .S0(\ConfigBits[474] ),
    .S1(\ConfigBits[475] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[474] ),
    .S1(\ConfigBits[475] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[474] ),
    .S1(\ConfigBits[475] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[476] ),
    .S1(\ConfigBits[477] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net34),
    .S0(\ConfigBits[478] ),
    .S1(\ConfigBits[479] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net158),
    .A2(net206),
    .A3(net208),
    .S0(\ConfigBits[478] ),
    .S1(\ConfigBits[479] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[478] ),
    .S1(\ConfigBits[479] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LG_O),
    .A3(M_EF),
    .S0(\ConfigBits[478] ),
    .S1(\ConfigBits[479] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JN2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[480] ),
    .S1(\ConfigBits[481] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JN2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst0  (.A0(net145),
    .A1(net5),
    .A2(net7),
    .A3(net25),
    .S0(\ConfigBits[514] ),
    .S1(\ConfigBits[515] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net211),
    .A3(net229),
    .S0(\ConfigBits[514] ),
    .S1(\ConfigBits[515] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst2  (.A0(LB_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[514] ),
    .S1(\ConfigBits[515] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[514] ),
    .S1(\ConfigBits[515] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[516] ),
    .S1(\ConfigBits[517] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst0  (.A0(net146),
    .A1(net2),
    .A2(net42),
    .A3(net22),
    .S0(\ConfigBits[518] ),
    .S1(\ConfigBits[519] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst1  (.A0(net182),
    .A1(net198),
    .A2(net212),
    .A3(net226),
    .S0(\ConfigBits[518] ),
    .S1(\ConfigBits[519] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[518] ),
    .S1(\ConfigBits[519] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[518] ),
    .S1(\ConfigBits[519] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[520] ),
    .S1(\ConfigBits[521] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst0  (.A0(net147),
    .A1(net3),
    .A2(net9),
    .A3(net25),
    .S0(\ConfigBits[522] ),
    .S1(\ConfigBits[523] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst1  (.A0(net161),
    .A1(net183),
    .A2(net213),
    .A3(net229),
    .S0(\ConfigBits[522] ),
    .S1(\ConfigBits[523] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[522] ),
    .S1(\ConfigBits[523] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[522] ),
    .S1(\ConfigBits[523] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[524] ),
    .S1(\ConfigBits[525] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst0  (.A0(net110),
    .A1(net4),
    .A2(net10),
    .A3(net22),
    .S0(\ConfigBits[526] ),
    .S1(\ConfigBits[527] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst1  (.A0(net162),
    .A1(net174),
    .A2(net214),
    .A3(net246),
    .S0(\ConfigBits[526] ),
    .S1(\ConfigBits[527] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LE_O),
    .S0(\ConfigBits[526] ),
    .S1(\ConfigBits[527] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[526] ),
    .S1(\ConfigBits[527] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[528] ),
    .S1(\ConfigBits[529] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[530] ),
    .S1(\ConfigBits[531] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net163),
    .A2(net207),
    .A3(net209),
    .S0(\ConfigBits[530] ),
    .S1(\ConfigBits[531] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[530] ),
    .S1(\ConfigBits[531] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[530] ),
    .S1(\ConfigBits[531] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[532] ),
    .S1(\ConfigBits[533] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[534] ),
    .S1(\ConfigBits[535] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst1  (.A0(net156),
    .A1(net164),
    .A2(net206),
    .A3(net208),
    .S0(\ConfigBits[534] ),
    .S1(\ConfigBits[535] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[534] ),
    .S1(\ConfigBits[535] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[534] ),
    .S1(\ConfigBits[535] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[536] ),
    .S1(\ConfigBits[537] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\ConfigBits[538] ),
    .S1(\ConfigBits[539] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst1  (.A0(net157),
    .A1(net165),
    .A2(net207),
    .A3(net209),
    .S0(\ConfigBits[538] ),
    .S1(\ConfigBits[539] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[538] ),
    .S1(\ConfigBits[539] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[538] ),
    .S1(\ConfigBits[539] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[540] ),
    .S1(\ConfigBits[541] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net106),
    .A2(net2),
    .A3(net6),
    .S0(\ConfigBits[542] ),
    .S1(\ConfigBits[543] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net158),
    .A2(net206),
    .A3(net208),
    .S0(\ConfigBits[542] ),
    .S1(\ConfigBits[543] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[542] ),
    .S1(\ConfigBits[543] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LG_O),
    .A3(M_AD),
    .S0(\ConfigBits[542] ),
    .S1(\ConfigBits[543] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JS2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[544] ),
    .S1(\ConfigBits[545] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JS2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net107),
    .A2(net7),
    .A3(net25),
    .S0(\ConfigBits[546] ),
    .S1(\ConfigBits[547] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst1  (.A0(net159),
    .A1(net181),
    .A2(net211),
    .A3(net229),
    .S0(\ConfigBits[546] ),
    .S1(\ConfigBits[547] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst2  (.A0(LB_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[546] ),
    .S1(\ConfigBits[547] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[546] ),
    .S1(\ConfigBits[547] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[548] ),
    .S1(\ConfigBits[549] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net108),
    .A2(net8),
    .A3(net22),
    .S0(\ConfigBits[550] ),
    .S1(\ConfigBits[551] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst1  (.A0(net160),
    .A1(net182),
    .A2(net212),
    .A3(net226),
    .S0(\ConfigBits[550] ),
    .S1(\ConfigBits[551] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LC_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[550] ),
    .S1(\ConfigBits[551] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[550] ),
    .S1(\ConfigBits[551] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[552] ),
    .S1(\ConfigBits[553] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net109),
    .A2(net43),
    .A3(net25),
    .S0(\ConfigBits[554] ),
    .S1(\ConfigBits[555] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst1  (.A0(net183),
    .A1(net199),
    .A2(net213),
    .A3(net229),
    .S0(\ConfigBits[554] ),
    .S1(\ConfigBits[555] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LD_O),
    .A3(LE_O),
    .S0(\ConfigBits[554] ),
    .S1(\ConfigBits[555] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[554] ),
    .S1(\ConfigBits[555] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG2/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[556] ),
    .S1(\ConfigBits[557] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net110),
    .A2(net10),
    .A3(net22),
    .S0(\ConfigBits[558] ),
    .S1(\ConfigBits[559] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst1  (.A0(net162),
    .A1(net174),
    .A2(net214),
    .A3(net246),
    .S0(\ConfigBits[558] ),
    .S1(\ConfigBits[559] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LE_O),
    .S0(\ConfigBits[558] ),
    .S1(\ConfigBits[559] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AB),
    .S0(\ConfigBits[558] ),
    .S1(\ConfigBits[559] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG3/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[560] ),
    .S1(\ConfigBits[561] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net111),
    .A2(net3),
    .A3(net11),
    .S0(\ConfigBits[562] ),
    .S1(\ConfigBits[563] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net163),
    .A3(net207),
    .S0(\ConfigBits[562] ),
    .S1(\ConfigBits[563] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[562] ),
    .S1(\ConfigBits[563] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst3  (.A0(LF_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AD),
    .S0(\ConfigBits[562] ),
    .S1(\ConfigBits[563] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG4/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[564] ),
    .S1(\ConfigBits[565] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[4] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net112),
    .A2(net4),
    .A3(net12),
    .S0(\ConfigBits[566] ),
    .S1(\ConfigBits[567] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net164),
    .A3(net208),
    .S0(\ConfigBits[566] ),
    .S1(\ConfigBits[567] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[566] ),
    .S1(\ConfigBits[567] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LG_O),
    .A2(LH_O),
    .A3(M_AH),
    .S0(\ConfigBits[566] ),
    .S1(\ConfigBits[567] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG5/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[568] ),
    .S1(\ConfigBits[569] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[5] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net113),
    .A2(net5),
    .A3(net13),
    .S0(\ConfigBits[570] ),
    .S1(\ConfigBits[571] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst1  (.A0(net155),
    .A1(net157),
    .A2(net165),
    .A3(net209),
    .S0(\ConfigBits[570] ),
    .S1(\ConfigBits[571] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[570] ),
    .S1(\ConfigBits[571] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LH_O),
    .A3(M_EF),
    .S0(\ConfigBits[570] ),
    .S1(\ConfigBits[571] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG6/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[572] ),
    .S1(\ConfigBits[573] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[6] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net138),
    .A2(net2),
    .A3(net6),
    .S0(\ConfigBits[574] ),
    .S1(\ConfigBits[575] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst1  (.A0(net154),
    .A1(net156),
    .A2(net158),
    .A3(net206),
    .S0(\ConfigBits[574] ),
    .S1(\ConfigBits[575] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst2  (.A0(LA_O),
    .A1(LB_O),
    .A2(LC_O),
    .A3(LD_O),
    .S0(\ConfigBits[574] ),
    .S1(\ConfigBits[575] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst3  (.A0(LE_O),
    .A1(LF_O),
    .A2(LG_O),
    .A3(M_AB),
    .S0(\ConfigBits[574] ),
    .S1(\ConfigBits[575] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_JW2BEG7/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[576] ),
    .S1(\ConfigBits[577] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\JW2BEG[7] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst0  (.A0(net5),
    .A1(net209),
    .A2(LA_O),
    .A3(LB_O),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(LD_O),
    .A2(LE_O),
    .A3(LF_O),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst2  (.A0(LG_O),
    .A1(LH_O),
    .A2(M_AB),
    .A3(M_AH),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst3  (.A0(\J2MID_ABb_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2MID_EFb_BEG[1] ),
    .A3(\J2MID_GHb_BEG[1] ),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG0/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[260] ),
    .S1(\ConfigBits[261] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net481));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net208),
    .A2(LA_O),
    .A3(LB_O),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(LD_O),
    .A2(LE_O),
    .A3(LF_O),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst2  (.A0(LG_O),
    .A1(LH_O),
    .A2(M_AD),
    .A3(M_EF),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst3  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_CDa_BEG[2] ),
    .A2(\J2MID_EFa_BEG[2] ),
    .A3(\J2MID_GHa_BEG[2] ),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_inst4  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out1 ),
    .A2(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out2 ),
    .A3(\Inst_LUT4AB_switch_matrix/inst_cus_mux161_buf_W6BEG1/cus_mux41_buf_out3 ),
    .S0(\ConfigBits[264] ),
    .S1(\ConfigBits[265] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net482));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_EN/_0_  (.A0(net516),
    .A1(J_EN_BEG),
    .S(\ConfigBits[266] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_EN/_0__516  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net516));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_SR/_0_  (.A0(net508),
    .A1(J_SR_BEG),
    .S(\ConfigBits[275] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LA_SR/_0__508  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net508));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_EN/_0_  (.A0(net517),
    .A1(J_EN_BEG),
    .S(\ConfigBits[276] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_EN/_0__517  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net517));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_SR/_0_  (.A0(net509),
    .A1(J_SR_BEG),
    .S(\ConfigBits[285] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LB_SR/_0__509  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net509));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_EN/_0_  (.A0(net518),
    .A1(J_EN_BEG),
    .S(\ConfigBits[286] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_EN/_0__518  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net518));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_SR/_0_  (.A0(net510),
    .A1(J_SR_BEG),
    .S(\ConfigBits[295] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LC_SR/_0__510  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net510));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_EN/_0_  (.A0(net519),
    .A1(J_EN_BEG),
    .S(\ConfigBits[296] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_EN/_0__519  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net519));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_SR/_0_  (.A0(net511),
    .A1(J_SR_BEG),
    .S(\ConfigBits[305] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LD_SR/_0__511  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net511));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_EN/_0_  (.A0(net520),
    .A1(J_EN_BEG),
    .S(\ConfigBits[306] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_EN/_0__520  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net520));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_SR/_0_  (.A0(net512),
    .A1(J_SR_BEG),
    .S(\ConfigBits[315] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LE_SR/_0__512  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net512));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_EN/_0_  (.A0(net521),
    .A1(J_EN_BEG),
    .S(\ConfigBits[316] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_EN/_0__521  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net521));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_SR/_0_  (.A0(net513),
    .A1(J_SR_BEG),
    .S(\ConfigBits[325] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LF_SR/_0__513  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net513));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_EN/_0_  (.A0(net522),
    .A1(J_EN_BEG),
    .S(\ConfigBits[326] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_EN/_0__522  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net522));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_SR/_0_  (.A0(net514),
    .A1(J_SR_BEG),
    .S(\ConfigBits[335] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LG_SR/_0__514  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net514));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_EN/_0_  (.A0(net523),
    .A1(J_EN_BEG),
    .S(\ConfigBits[336] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_EN));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_EN/_0__523  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .HI(net523));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_SR/_0_  (.A0(net515),
    .A1(J_SR_BEG),
    .S(\ConfigBits[345] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_SR));
 sky130_fd_sc_hd__conb_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux21_LH_SR/_0__515  (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .LO(net515));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG0  (.A0(LD_O),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JN2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[182] ),
    .S1(\ConfigBits[183] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net255));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG1  (.A0(LE_O),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JN2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[184] ),
    .S1(\ConfigBits[185] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net256));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG2  (.A0(LF_O),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JN2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[186] ),
    .S1(\ConfigBits[187] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net257));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_E1BEG3  (.A0(LG_O),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JN2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[188] ),
    .S1(\ConfigBits[189] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net258));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG0  (.A0(net112),
    .A1(net12),
    .A2(net199),
    .A3(net216),
    .S0(\ConfigBits[418] ),
    .S1(\ConfigBits[419] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG1  (.A0(net138),
    .A1(net8),
    .A2(net160),
    .A3(net212),
    .S0(\ConfigBits[420] ),
    .S1(\ConfigBits[421] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG2  (.A0(net110),
    .A1(net34),
    .A2(net162),
    .A3(net214),
    .S0(\ConfigBits[422] ),
    .S1(\ConfigBits[423] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_AB_BEG3  (.A0(net106),
    .A1(net6),
    .A2(net158),
    .A3(net247),
    .S0(\ConfigBits[424] ),
    .S1(\ConfigBits[425] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG0  (.A0(net147),
    .A1(net12),
    .A2(net164),
    .A3(net216),
    .S0(\ConfigBits[426] ),
    .S1(\ConfigBits[427] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG1  (.A0(net108),
    .A1(net8),
    .A2(net160),
    .A3(net246),
    .S0(\ConfigBits[428] ),
    .S1(\ConfigBits[429] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG2  (.A0(net110),
    .A1(net10),
    .A2(net198),
    .A3(net214),
    .S0(\ConfigBits[430] ),
    .S1(\ConfigBits[431] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_CD_BEG3  (.A0(net106),
    .A1(net41),
    .A2(net158),
    .A3(net210),
    .S0(\ConfigBits[432] ),
    .S1(\ConfigBits[433] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG0  (.A0(net113),
    .A1(net42),
    .A2(net165),
    .A3(net217),
    .S0(\ConfigBits[434] ),
    .S1(\ConfigBits[435] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG1  (.A0(net109),
    .A1(net9),
    .A2(net161),
    .A3(net245),
    .S0(\ConfigBits[436] ),
    .S1(\ConfigBits[437] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG2  (.A0(net111),
    .A1(net11),
    .A2(net197),
    .A3(net215),
    .S0(\ConfigBits[438] ),
    .S1(\ConfigBits[439] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_EF_BEG3  (.A0(net146),
    .A1(net7),
    .A2(net159),
    .A3(net211),
    .S0(\ConfigBits[440] ),
    .S1(\ConfigBits[441] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG0  (.A0(net113),
    .A1(net13),
    .A2(net165),
    .A3(net238),
    .S0(\ConfigBits[442] ),
    .S1(\ConfigBits[443] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG1  (.A0(net109),
    .A1(net9),
    .A2(net190),
    .A3(net213),
    .S0(\ConfigBits[444] ),
    .S1(\ConfigBits[445] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG2  (.A0(net145),
    .A1(net11),
    .A2(net163),
    .A3(net215),
    .S0(\ConfigBits[446] ),
    .S1(\ConfigBits[447] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2END_GH_BEG3  (.A0(net107),
    .A1(net43),
    .A2(net159),
    .A3(net211),
    .S0(\ConfigBits[448] ),
    .S1(\ConfigBits[449] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2END_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG0  (.A0(net120),
    .A1(net172),
    .A2(net224),
    .A3(\JN2BEG[3] ),
    .S0(\ConfigBits[354] ),
    .S1(\ConfigBits[355] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG1  (.A0(net16),
    .A1(net168),
    .A2(net220),
    .A3(\JE2BEG[3] ),
    .S0(\ConfigBits[356] ),
    .S1(\ConfigBits[357] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net222),
    .A3(\JS2BEG[3] ),
    .S0(\ConfigBits[358] ),
    .S1(\ConfigBits[359] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABa_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net166),
    .A3(\JW2BEG[3] ),
    .S0(\ConfigBits[360] ),
    .S1(\ConfigBits[361] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\ConfigBits[386] ),
    .S1(\ConfigBits[387] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\ConfigBits[388] ),
    .S1(\ConfigBits[389] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABb_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\ConfigBits[390] ),
    .S1(\ConfigBits[391] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_ABb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\ConfigBits[392] ),
    .S1(\ConfigBits[393] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_ABb_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG0  (.A0(net20),
    .A1(net172),
    .A2(net224),
    .A3(\JN2BEG[4] ),
    .S0(\ConfigBits[362] ),
    .S1(\ConfigBits[363] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net220),
    .A3(\JE2BEG[4] ),
    .S0(\ConfigBits[364] ),
    .S1(\ConfigBits[365] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG2  (.A0(net118),
    .A1(net18),
    .A2(net170),
    .A3(\JS2BEG[4] ),
    .S0(\ConfigBits[366] ),
    .S1(\ConfigBits[367] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDa_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDa_BEG3  (.A0(net114),
    .A1(net166),
    .A2(net218),
    .A3(\JW2BEG[4] ),
    .S0(\ConfigBits[368] ),
    .S1(\ConfigBits[369] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\ConfigBits[394] ),
    .S1(\ConfigBits[395] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\ConfigBits[396] ),
    .S1(\ConfigBits[397] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\ConfigBits[398] ),
    .S1(\ConfigBits[399] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_CDb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\ConfigBits[400] ),
    .S1(\ConfigBits[401] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_CDb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net224),
    .A3(\JN2BEG[5] ),
    .S0(\ConfigBits[370] ),
    .S1(\ConfigBits[371] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG1  (.A0(net116),
    .A1(net16),
    .A2(net168),
    .A3(\JE2BEG[5] ),
    .S0(\ConfigBits[372] ),
    .S1(\ConfigBits[373] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG2  (.A0(net118),
    .A1(net170),
    .A2(net222),
    .A3(\JS2BEG[5] ),
    .S0(\ConfigBits[374] ),
    .S1(\ConfigBits[375] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFa_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFa_BEG3  (.A0(net14),
    .A1(net166),
    .A2(net218),
    .A3(\JW2BEG[5] ),
    .S0(\ConfigBits[376] ),
    .S1(\ConfigBits[377] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFa_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\ConfigBits[402] ),
    .S1(\ConfigBits[403] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\ConfigBits[404] ),
    .S1(\ConfigBits[405] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\ConfigBits[406] ),
    .S1(\ConfigBits[407] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFb_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_EFb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\ConfigBits[408] ),
    .S1(\ConfigBits[409] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_EFb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG0  (.A0(net120),
    .A1(net20),
    .A2(net172),
    .A3(\JN2BEG[6] ),
    .S0(\ConfigBits[378] ),
    .S1(\ConfigBits[379] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHa_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG1  (.A0(net116),
    .A1(net168),
    .A2(net220),
    .A3(\JE2BEG[6] ),
    .S0(\ConfigBits[380] ),
    .S1(\ConfigBits[381] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHa_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG2  (.A0(net18),
    .A1(net170),
    .A2(net222),
    .A3(\JS2BEG[6] ),
    .S0(\ConfigBits[382] ),
    .S1(\ConfigBits[383] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHa_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHa_BEG3  (.A0(net114),
    .A1(net14),
    .A2(net218),
    .A3(\JW2BEG[6] ),
    .S0(\ConfigBits[384] ),
    .S1(\ConfigBits[385] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHa_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG0  (.A0(net121),
    .A1(net21),
    .A2(net173),
    .A3(net225),
    .S0(\ConfigBits[410] ),
    .S1(\ConfigBits[411] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHb_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG1  (.A0(net117),
    .A1(net17),
    .A2(net169),
    .A3(net221),
    .S0(\ConfigBits[412] ),
    .S1(\ConfigBits[413] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHb_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG2  (.A0(net119),
    .A1(net19),
    .A2(net171),
    .A3(net223),
    .S0(\ConfigBits[414] ),
    .S1(\ConfigBits[415] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHb_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J2MID_GHb_BEG3  (.A0(net115),
    .A1(net15),
    .A2(net167),
    .A3(net219),
    .S0(\ConfigBits[416] ),
    .S1(\ConfigBits[417] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J2MID_GHb_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG0  (.A0(net147),
    .A1(net183),
    .A2(net238),
    .A3(\JN2BEG[1] ),
    .S0(\ConfigBits[578] ),
    .S1(\ConfigBits[579] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_AB_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG1  (.A0(net42),
    .A1(net182),
    .A2(net217),
    .A3(\JE2BEG[1] ),
    .S0(\ConfigBits[580] ),
    .S1(\ConfigBits[581] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_AB_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG2  (.A0(net129),
    .A1(net25),
    .A2(net229),
    .A3(\JS2BEG[1] ),
    .S0(\ConfigBits[582] ),
    .S1(\ConfigBits[583] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_AB_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_AB_BEG3  (.A0(net122),
    .A1(net22),
    .A2(net174),
    .A3(\JW2BEG[1] ),
    .S0(\ConfigBits[584] ),
    .S1(\ConfigBits[585] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_AB_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG0  (.A0(net9),
    .A1(net199),
    .A2(net246),
    .A3(\JN2BEG[2] ),
    .S0(\ConfigBits[586] ),
    .S1(\ConfigBits[587] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_CD_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG1  (.A0(net130),
    .A1(net8),
    .A2(net217),
    .A3(\JE2BEG[2] ),
    .S0(\ConfigBits[588] ),
    .S1(\ConfigBits[589] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_CD_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG2  (.A0(net145),
    .A1(net41),
    .A2(net181),
    .A3(\JS2BEG[2] ),
    .S0(\ConfigBits[590] ),
    .S1(\ConfigBits[591] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_CD_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_CD_BEG3  (.A0(net122),
    .A1(net190),
    .A2(net226),
    .A3(\JW2BEG[2] ),
    .S0(\ConfigBits[592] ),
    .S1(\ConfigBits[593] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_CD_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG0  (.A0(net131),
    .A1(net9),
    .A2(net213),
    .A3(\JN2BEG[3] ),
    .S0(\ConfigBits[594] ),
    .S1(\ConfigBits[595] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_EF_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG1  (.A0(net146),
    .A1(net8),
    .A2(net182),
    .A3(\JE2BEG[3] ),
    .S0(\ConfigBits[596] ),
    .S1(\ConfigBits[597] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_EF_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG2  (.A0(net129),
    .A1(net197),
    .A2(net214),
    .A3(\JS2BEG[3] ),
    .S0(\ConfigBits[598] ),
    .S1(\ConfigBits[599] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_EF_BEG[2] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_EF_BEG3  (.A0(net43),
    .A1(net174),
    .A2(net245),
    .A3(\JW2BEG[3] ),
    .S0(\ConfigBits[600] ),
    .S1(\ConfigBits[601] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_EF_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG0  (.A0(net131),
    .A1(net34),
    .A2(net183),
    .A3(\JN2BEG[4] ),
    .S0(\ConfigBits[602] ),
    .S1(\ConfigBits[603] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_GH_BEG[0] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG1  (.A0(net130),
    .A1(net198),
    .A2(net212),
    .A3(\JE2BEG[4] ),
    .S0(\ConfigBits[604] ),
    .S1(\ConfigBits[605] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_GH_BEG[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG2  (.A0(net25),
    .A1(net181),
    .A2(net247),
    .A3(\JS2BEG[4] ),
    .S0(\ConfigBits[606] ),
    .S1(\ConfigBits[607] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_GH_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_J_l_GH_BEG3  (.A0(net138),
    .A1(net22),
    .A2(net210),
    .A3(\JW2BEG[4] ),
    .S0(\ConfigBits[608] ),
    .S1(\ConfigBits[609] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\J_l_GH_BEG[3] ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I0  (.A0(\J2MID_ABa_BEG[0] ),
    .A1(\J2MID_ABb_BEG[0] ),
    .A2(\J2END_AB_BEG[0] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[267] ),
    .S1(\ConfigBits[268] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I1  (.A0(\J2MID_ABa_BEG[1] ),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2END_AB_BEG[1] ),
    .A3(\J_l_AB_BEG[1] ),
    .S0(\ConfigBits[269] ),
    .S1(\ConfigBits[270] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I2  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\J2END_AB_BEG[2] ),
    .A3(\J_l_AB_BEG[2] ),
    .S0(\ConfigBits[271] ),
    .S1(\ConfigBits[272] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LA_I3  (.A0(\J2MID_ABa_BEG[3] ),
    .A1(\J2MID_ABb_BEG[3] ),
    .A2(\J2END_AB_BEG[3] ),
    .A3(\J_l_AB_BEG[3] ),
    .S0(\ConfigBits[273] ),
    .S1(\ConfigBits[274] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LA_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I0  (.A0(\J2MID_ABa_BEG[0] ),
    .A1(\J2MID_ABb_BEG[0] ),
    .A2(\J2END_AB_BEG[0] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[277] ),
    .S1(\ConfigBits[278] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I1  (.A0(\J2MID_ABa_BEG[1] ),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2END_AB_BEG[1] ),
    .A3(\J_l_AB_BEG[1] ),
    .S0(\ConfigBits[279] ),
    .S1(\ConfigBits[280] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I2  (.A0(\J2MID_ABa_BEG[2] ),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\J2END_AB_BEG[2] ),
    .A3(\J_l_AB_BEG[2] ),
    .S0(\ConfigBits[281] ),
    .S1(\ConfigBits[282] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LB_I3  (.A0(\J2MID_ABa_BEG[3] ),
    .A1(\J2MID_ABb_BEG[3] ),
    .A2(\J2END_AB_BEG[3] ),
    .A3(\J_l_AB_BEG[3] ),
    .S0(\ConfigBits[283] ),
    .S1(\ConfigBits[284] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LB_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I0  (.A0(\J2MID_CDa_BEG[0] ),
    .A1(\J2MID_CDb_BEG[0] ),
    .A2(\J2END_CD_BEG[0] ),
    .A3(\J_l_CD_BEG[0] ),
    .S0(\ConfigBits[287] ),
    .S1(\ConfigBits[288] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I1  (.A0(\J2MID_CDa_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2END_CD_BEG[1] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[289] ),
    .S1(\ConfigBits[290] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I2  (.A0(\J2MID_CDa_BEG[2] ),
    .A1(\J2MID_CDb_BEG[2] ),
    .A2(\J2END_CD_BEG[2] ),
    .A3(\J_l_CD_BEG[2] ),
    .S0(\ConfigBits[291] ),
    .S1(\ConfigBits[292] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LC_I3  (.A0(\J2MID_CDa_BEG[3] ),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\J2END_CD_BEG[3] ),
    .A3(\J_l_CD_BEG[3] ),
    .S0(\ConfigBits[293] ),
    .S1(\ConfigBits[294] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LC_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I0  (.A0(\J2MID_CDa_BEG[0] ),
    .A1(\J2MID_CDb_BEG[0] ),
    .A2(\J2END_CD_BEG[0] ),
    .A3(\J_l_CD_BEG[0] ),
    .S0(\ConfigBits[297] ),
    .S1(\ConfigBits[298] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I1  (.A0(\J2MID_CDa_BEG[1] ),
    .A1(\J2MID_CDb_BEG[1] ),
    .A2(\J2END_CD_BEG[1] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[299] ),
    .S1(\ConfigBits[300] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I2  (.A0(\J2MID_CDa_BEG[2] ),
    .A1(\J2MID_CDb_BEG[2] ),
    .A2(\J2END_CD_BEG[2] ),
    .A3(\J_l_CD_BEG[2] ),
    .S0(\ConfigBits[301] ),
    .S1(\ConfigBits[302] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LD_I3  (.A0(\J2MID_CDa_BEG[3] ),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\J2END_CD_BEG[3] ),
    .A3(\J_l_CD_BEG[3] ),
    .S0(\ConfigBits[303] ),
    .S1(\ConfigBits[304] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LD_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I0  (.A0(\J2MID_EFa_BEG[0] ),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\J2END_EF_BEG[0] ),
    .A3(\J_l_EF_BEG[0] ),
    .S0(\ConfigBits[307] ),
    .S1(\ConfigBits[308] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I1  (.A0(\J2MID_EFa_BEG[1] ),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2END_EF_BEG[1] ),
    .A3(\J_l_EF_BEG[1] ),
    .S0(\ConfigBits[309] ),
    .S1(\ConfigBits[310] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I2  (.A0(\J2MID_EFa_BEG[2] ),
    .A1(\J2MID_EFb_BEG[2] ),
    .A2(\J2END_EF_BEG[2] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[311] ),
    .S1(\ConfigBits[312] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LE_I3  (.A0(\J2MID_EFa_BEG[3] ),
    .A1(\J2MID_EFb_BEG[3] ),
    .A2(\J2END_EF_BEG[3] ),
    .A3(\J_l_EF_BEG[3] ),
    .S0(\ConfigBits[313] ),
    .S1(\ConfigBits[314] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LE_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I0  (.A0(\J2MID_EFa_BEG[0] ),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\J2END_EF_BEG[0] ),
    .A3(\J_l_EF_BEG[0] ),
    .S0(\ConfigBits[317] ),
    .S1(\ConfigBits[318] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I1  (.A0(\J2MID_EFa_BEG[1] ),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2END_EF_BEG[1] ),
    .A3(\J_l_EF_BEG[1] ),
    .S0(\ConfigBits[319] ),
    .S1(\ConfigBits[320] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I2  (.A0(\J2MID_EFa_BEG[2] ),
    .A1(\J2MID_EFb_BEG[2] ),
    .A2(\J2END_EF_BEG[2] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[321] ),
    .S1(\ConfigBits[322] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LF_I3  (.A0(\J2MID_EFa_BEG[3] ),
    .A1(\J2MID_EFb_BEG[3] ),
    .A2(\J2END_EF_BEG[3] ),
    .A3(\J_l_EF_BEG[3] ),
    .S0(\ConfigBits[323] ),
    .S1(\ConfigBits[324] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LF_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I0  (.A0(\J2MID_GHa_BEG[0] ),
    .A1(\J2MID_GHb_BEG[0] ),
    .A2(\J2END_GH_BEG[0] ),
    .A3(\J_l_GH_BEG[0] ),
    .S0(\ConfigBits[327] ),
    .S1(\ConfigBits[328] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I1  (.A0(\J2MID_GHa_BEG[1] ),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\J2END_GH_BEG[1] ),
    .A3(\J_l_GH_BEG[1] ),
    .S0(\ConfigBits[329] ),
    .S1(\ConfigBits[330] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I2  (.A0(\J2MID_GHa_BEG[2] ),
    .A1(\J2MID_GHb_BEG[2] ),
    .A2(\J2END_GH_BEG[2] ),
    .A3(\J_l_GH_BEG[2] ),
    .S0(\ConfigBits[331] ),
    .S1(\ConfigBits[332] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LG_I3  (.A0(\J2MID_GHa_BEG[3] ),
    .A1(\J2MID_GHb_BEG[3] ),
    .A2(\J2END_GH_BEG[3] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[333] ),
    .S1(\ConfigBits[334] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LG_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I0  (.A0(\J2MID_GHa_BEG[0] ),
    .A1(\J2MID_GHb_BEG[0] ),
    .A2(\J2END_GH_BEG[0] ),
    .A3(\J_l_GH_BEG[0] ),
    .S0(\ConfigBits[337] ),
    .S1(\ConfigBits[338] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I1  (.A0(\J2MID_GHa_BEG[1] ),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\J2END_GH_BEG[1] ),
    .A3(\J_l_GH_BEG[1] ),
    .S0(\ConfigBits[339] ),
    .S1(\ConfigBits[340] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I2  (.A0(\J2MID_GHa_BEG[2] ),
    .A1(\J2MID_GHb_BEG[2] ),
    .A2(\J2END_GH_BEG[2] ),
    .A3(\J_l_GH_BEG[2] ),
    .S0(\ConfigBits[341] ),
    .S1(\ConfigBits[342] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_I2));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_LH_I3  (.A0(\J2MID_GHa_BEG[3] ),
    .A1(\J2MID_GHb_BEG[3] ),
    .A2(\J2END_GH_BEG[3] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[343] ),
    .S1(\ConfigBits[344] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(LH_I3));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(LC_O),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JW2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[154] ),
    .S1(\ConfigBits[155] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net355));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(LD_O),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JW2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[156] ),
    .S1(\ConfigBits[157] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(LE_O),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JW2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[158] ),
    .S1(\ConfigBits[159] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net357));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(LF_O),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JW2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[160] ),
    .S1(\ConfigBits[161] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net358));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG0  (.A0(net108),
    .A1(net129),
    .A2(net25),
    .A3(LE_O),
    .S0(\ConfigBits[162] ),
    .S1(\ConfigBits[163] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG1  (.A0(net109),
    .A1(net130),
    .A2(net22),
    .A3(LF_O),
    .S0(\ConfigBits[164] ),
    .S1(\ConfigBits[165] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG2  (.A0(net106),
    .A1(net131),
    .A2(net229),
    .A3(LG_O),
    .S0(\ConfigBits[166] ),
    .S1(\ConfigBits[167] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net380));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_N4BEG3  (.A0(net107),
    .A1(net122),
    .A2(net226),
    .A3(LH_O),
    .S0(\ConfigBits[168] ),
    .S1(\ConfigBits[169] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net381));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S0  (.A0(\JN2BEG[4] ),
    .A1(\JE2BEG[4] ),
    .A2(\JS2BEG[4] ),
    .A3(\JW2BEG[4] ),
    .S0(\ConfigBits[346] ),
    .S1(\ConfigBits[347] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S0));
 sky130_fd_sc_hd__mux4_2 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1  (.A0(\JN2BEG[5] ),
    .A1(\JE2BEG[5] ),
    .A2(\JS2BEG[5] ),
    .A3(\JW2BEG[5] ),
    .S0(\ConfigBits[348] ),
    .S1(\ConfigBits[349] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S1));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(LE_O),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JE2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[210] ),
    .S1(\ConfigBits[211] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net407));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(LF_O),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JE2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[212] ),
    .S1(\ConfigBits[213] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net408));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(LG_O),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JE2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[214] ),
    .S1(\ConfigBits[215] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net409));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(LH_O),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JE2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[216] ),
    .S1(\ConfigBits[217] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net410));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S2  (.A0(\JN2BEG[6] ),
    .A1(\JE2BEG[6] ),
    .A2(\JS2BEG[6] ),
    .A3(\JW2BEG[6] ),
    .S0(\ConfigBits[350] ),
    .S1(\ConfigBits[351] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S3  (.A0(\JN2BEG[7] ),
    .A1(\JE2BEG[7] ),
    .A2(\JS2BEG[7] ),
    .A3(\JW2BEG[7] ),
    .S0(\ConfigBits[352] ),
    .S1(\ConfigBits[353] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S3));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG0  (.A0(net25),
    .A1(net160),
    .A2(net181),
    .A3(LA_O),
    .S0(\ConfigBits[218] ),
    .S1(\ConfigBits[219] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net430));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG1  (.A0(net22),
    .A1(net161),
    .A2(net182),
    .A3(LB_O),
    .S0(\ConfigBits[220] ),
    .S1(\ConfigBits[221] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net431));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG2  (.A0(net158),
    .A1(net183),
    .A2(net229),
    .A3(LC_O),
    .S0(\ConfigBits[222] ),
    .S1(\ConfigBits[223] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net432));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_S4BEG3  (.A0(net159),
    .A1(net174),
    .A2(net226),
    .A3(LD_O),
    .S0(\ConfigBits[224] ),
    .S1(\ConfigBits[225] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net433));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(LF_O),
    .A1(\J2MID_CDb_BEG[3] ),
    .A2(\JS2BEG[3] ),
    .A3(\J_l_CD_BEG[1] ),
    .S0(\ConfigBits[238] ),
    .S1(\ConfigBits[239] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net460));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(LG_O),
    .A1(\J2MID_EFb_BEG[0] ),
    .A2(\JS2BEG[0] ),
    .A3(\J_l_EF_BEG[2] ),
    .S0(\ConfigBits[240] ),
    .S1(\ConfigBits[241] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net461));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(LH_O),
    .A1(\J2MID_GHb_BEG[1] ),
    .A2(\JS2BEG[1] ),
    .A3(\J_l_GH_BEG[3] ),
    .S0(\ConfigBits[242] ),
    .S1(\ConfigBits[243] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net462));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(LA_O),
    .A1(\J2MID_ABb_BEG[2] ),
    .A2(\JS2BEG[2] ),
    .A3(\J_l_AB_BEG[0] ),
    .S0(\ConfigBits[244] ),
    .S1(\ConfigBits[245] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net463));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net156),
    .A3(LF_O),
    .S0(\ConfigBits[190] ),
    .S1(\ConfigBits[191] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_inst1  (.A0(LG_O),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[0] ),
    .S0(\ConfigBits[190] ),
    .S1(\ConfigBits[191] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[192] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net290));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net157),
    .A3(LA_O),
    .S0(\ConfigBits[193] ),
    .S1(\ConfigBits[194] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_inst1  (.A0(LH_O),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[0] ),
    .S0(\ConfigBits[193] ),
    .S1(\ConfigBits[194] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[195] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net291));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net154),
    .A3(LB_O),
    .S0(\ConfigBits[196] ),
    .S1(\ConfigBits[197] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[0] ),
    .S0(\ConfigBits[196] ),
    .S1(\ConfigBits[197] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[198] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net292));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net155),
    .A3(LD_O),
    .S0(\ConfigBits[199] ),
    .S1(\ConfigBits[200] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_inst1  (.A0(LE_O),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[0] ),
    .S0(\ConfigBits[199] ),
    .S1(\ConfigBits[200] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_EE4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[201] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net293));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst0  (.A0(\J2MID_GHa_BEG[3] ),
    .A1(\J2MID_ABb_BEG[3] ),
    .A2(\J2MID_CDb_BEG[3] ),
    .A3(\J2MID_EFb_BEG[3] ),
    .S0(\ConfigBits[613] ),
    .S1(\ConfigBits[614] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_inst1  (.A0(\JN2BEG[2] ),
    .A1(\JE2BEG[2] ),
    .A2(\JS2BEG[2] ),
    .A3(\JW2BEG[2] ),
    .S0(\ConfigBits[613] ),
    .S1(\ConfigBits[614] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_4 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_EN_BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[615] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(J_EN_BEG));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst0  (.A0(\J2MID_GHa_BEG[0] ),
    .A1(\J2MID_ABb_BEG[0] ),
    .A2(\J2MID_CDb_BEG[0] ),
    .A3(\J2MID_EFb_BEG[0] ),
    .S0(\ConfigBits[610] ),
    .S1(\ConfigBits[611] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_inst1  (.A0(\JN2BEG[1] ),
    .A1(\JE2BEG[1] ),
    .A2(\JS2BEG[1] ),
    .A3(\JW2BEG[1] ),
    .S0(\ConfigBits[610] ),
    .S1(\ConfigBits[611] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_4 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_J_SR_BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[612] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(J_SR_BEG));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net208),
    .A3(LF_O),
    .S0(\ConfigBits[170] ),
    .S1(\ConfigBits[171] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_inst1  (.A0(LG_O),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[1] ),
    .S0(\ConfigBits[170] ),
    .S1(\ConfigBits[171] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[172] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net394));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net209),
    .A3(LA_O),
    .S0(\ConfigBits[173] ),
    .S1(\ConfigBits[174] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_inst1  (.A0(LH_O),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[1] ),
    .S0(\ConfigBits[173] ),
    .S1(\ConfigBits[174] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[175] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net395));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net206),
    .A3(LB_O),
    .S0(\ConfigBits[176] ),
    .S1(\ConfigBits[177] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[1] ),
    .S0(\ConfigBits[176] ),
    .S1(\ConfigBits[177] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[178] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net396));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net207),
    .A3(LD_O),
    .S0(\ConfigBits[179] ),
    .S1(\ConfigBits[180] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_inst1  (.A0(LE_O),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[1] ),
    .S0(\ConfigBits[179] ),
    .S1(\ConfigBits[180] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_NN4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[181] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net397));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net4),
    .A2(net208),
    .A3(LF_O),
    .S0(\ConfigBits[226] ),
    .S1(\ConfigBits[227] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_inst1  (.A0(LG_O),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[3] ),
    .S0(\ConfigBits[226] ),
    .S1(\ConfigBits[227] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[228] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net446));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net5),
    .A2(net209),
    .A3(LA_O),
    .S0(\ConfigBits[229] ),
    .S1(\ConfigBits[230] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_inst1  (.A0(LH_O),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[3] ),
    .S0(\ConfigBits[229] ),
    .S1(\ConfigBits[230] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[231] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net447));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net2),
    .A2(net206),
    .A3(LB_O),
    .S0(\ConfigBits[232] ),
    .S1(\ConfigBits[233] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[3] ),
    .S0(\ConfigBits[232] ),
    .S1(\ConfigBits[233] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[234] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net448));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net3),
    .A2(net207),
    .A3(LD_O),
    .S0(\ConfigBits[235] ),
    .S1(\ConfigBits[236] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_inst1  (.A0(LE_O),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[3] ),
    .S0(\ConfigBits[235] ),
    .S1(\ConfigBits[236] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_SS4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[237] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net449));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst0  (.A0(net104),
    .A1(net156),
    .A2(net208),
    .A3(LF_O),
    .S0(\ConfigBits[246] ),
    .S1(\ConfigBits[247] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_inst1  (.A0(LG_O),
    .A1(\J2MID_ABb_BEG[1] ),
    .A2(\J2MID_CDb_BEG[1] ),
    .A3(\J2END_GH_BEG[2] ),
    .S0(\ConfigBits[246] ),
    .S1(\ConfigBits[247] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG0/cus_mux41_buf_out1 ),
    .S(\ConfigBits[248] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net495));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst0  (.A0(net105),
    .A1(net157),
    .A2(net209),
    .A3(LA_O),
    .S0(\ConfigBits[249] ),
    .S1(\ConfigBits[250] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_inst1  (.A0(LH_O),
    .A1(\J2MID_ABa_BEG[2] ),
    .A2(\J2MID_CDa_BEG[2] ),
    .A3(\J2END_EF_BEG[2] ),
    .S0(\ConfigBits[249] ),
    .S1(\ConfigBits[250] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG1/cus_mux41_buf_out1 ),
    .S(\ConfigBits[251] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net496));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst0  (.A0(net102),
    .A1(net154),
    .A2(net206),
    .A3(LB_O),
    .S0(\ConfigBits[252] ),
    .S1(\ConfigBits[253] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_inst1  (.A0(LC_O),
    .A1(\J2MID_EFb_BEG[1] ),
    .A2(\J2MID_GHb_BEG[1] ),
    .A3(\J2END_CD_BEG[2] ),
    .S0(\ConfigBits[252] ),
    .S1(\ConfigBits[253] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG2/cus_mux41_buf_out1 ),
    .S(\ConfigBits[254] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net497));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst0  (.A0(net103),
    .A1(net155),
    .A2(net207),
    .A3(LD_O),
    .S0(\ConfigBits[255] ),
    .S1(\ConfigBits[256] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_inst1  (.A0(LE_O),
    .A1(\J2MID_EFa_BEG[2] ),
    .A2(\J2MID_GHa_BEG[2] ),
    .A3(\J2END_AB_BEG[2] ),
    .S0(\ConfigBits[255] ),
    .S1(\ConfigBits[256] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__mux2_1 \Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/my_mux2_inst/_0_  (.A0(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out0 ),
    .A1(\Inst_LUT4AB_switch_matrix/inst_cus_mux81_buf_WW4BEG3/cus_mux41_buf_out1 ),
    .S(\ConfigBits[257] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net498));
 sky130_fd_sc_hd__mux2_8 \Inst_MUX8LUT_frame_config_mux/cus_mux21_AB/_0_  (.A0(A),
    .A1(B),
    .S(S0),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(M_AB));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_AD/_0_  (.A0(M_AB),
    .A1(\Inst_MUX8LUT_frame_config_mux/CD ),
    .S(S1),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/AD ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_AH/_0_  (.A0(\Inst_MUX8LUT_frame_config_mux/AD ),
    .A1(\Inst_MUX8LUT_frame_config_mux/EH ),
    .S(S3),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/AH ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_CD/_0_  (.A0(C),
    .A1(D),
    .S(\Inst_MUX8LUT_frame_config_mux/sCD ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/CD ));
 sky130_fd_sc_hd__mux2_4 \Inst_MUX8LUT_frame_config_mux/cus_mux21_EF/_0_  (.A0(E),
    .A1(F),
    .S(\Inst_MUX8LUT_frame_config_mux/sEF ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(M_EF));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_EH/_0_  (.A0(M_EF),
    .A1(\Inst_MUX8LUT_frame_config_mux/GH ),
    .S(\Inst_MUX8LUT_frame_config_mux/sEH ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/EH ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_EH_GH/_0_  (.A0(\Inst_MUX8LUT_frame_config_mux/GH ),
    .A1(\Inst_MUX8LUT_frame_config_mux/EH ),
    .S(\ConfigBits[152] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/EH_GH ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_GH/_0_  (.A0(G),
    .A1(H),
    .S(\Inst_MUX8LUT_frame_config_mux/sGH ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/GH ));
 sky130_fd_sc_hd__mux2_4 \Inst_MUX8LUT_frame_config_mux/cus_mux21_M_AD/_0_  (.A0(\Inst_MUX8LUT_frame_config_mux/CD ),
    .A1(\Inst_MUX8LUT_frame_config_mux/AD ),
    .S(\ConfigBits[152] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(M_AD));
 sky130_fd_sc_hd__mux2_4 \Inst_MUX8LUT_frame_config_mux/cus_mux21_M_AH/_0_  (.A0(\Inst_MUX8LUT_frame_config_mux/EH_GH ),
    .A1(\Inst_MUX8LUT_frame_config_mux/AH ),
    .S(\ConfigBits[153] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(M_AH));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_sCD/_0_  (.A0(S1),
    .A1(S0),
    .S(\ConfigBits[152] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/sCD ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_sEF/_0_  (.A0(S2),
    .A1(S0),
    .S(\ConfigBits[153] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/sEF ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_sEH/_0_  (.A0(S3),
    .A1(S1),
    .S(\ConfigBits[153] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/sEH ));
 sky130_fd_sc_hd__mux2_1 \Inst_MUX8LUT_frame_config_mux/cus_mux21_sGH/_0_  (.A0(\Inst_MUX8LUT_frame_config_mux/sEH ),
    .A1(\Inst_MUX8LUT_frame_config_mux/sEF ),
    .S(\ConfigBits[152] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\Inst_MUX8LUT_frame_config_mux/sGH ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_0/_0_  (.A(\N4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_1/_0_  (.A(\N4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_10/_0_  (.A(\N4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_11/_0_  (.A(\N4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_2/_0_  (.A(\N4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_3/_0_  (.A(\N4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_4/_0_  (.A(\N4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_5/_0_  (.A(\N4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_6/_0_  (.A(\N4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_7/_0_  (.A(\N4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_8/_0_  (.A(\N4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_9/_0_  (.A(\N4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net390));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_0/_0_  (.A(net132),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_1/_0_  (.A(net133),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_10/_0_  (.A(net127),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_11/_0_  (.A(net128),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_4 \N4END_inbuf_2/_0_  (.A(net134),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_3/_0_  (.A(net135),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_4/_0_  (.A(net136),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_5/_0_  (.A(net137),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[5] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_6/_0_  (.A(net123),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_7/_0_  (.A(net124),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_8/_0_  (.A(net125),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_9/_0_  (.A(net126),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\N4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_0/_0_  (.A(\NN4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_1/_0_  (.A(\NN4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_10/_0_  (.A(\NN4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_11/_0_  (.A(\NN4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_2/_0_  (.A(\NN4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_3/_0_  (.A(\NN4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_4/_0_  (.A(\NN4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_5/_0_  (.A(\NN4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_6/_0_  (.A(\NN4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_7/_0_  (.A(\NN4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_8/_0_  (.A(\NN4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 \NN4BEG_outbuf_9/_0_  (.A(\NN4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_0/_0_  (.A(net148),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_1/_0_  (.A(net149),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_10/_0_  (.A(net143),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_11/_0_  (.A(net144),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_2/_0_  (.A(net150),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_3/_0_  (.A(net151),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_4/_0_  (.A(net152),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_4 \NN4END_inbuf_5/_0_  (.A(net153),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_6/_0_  (.A(net139),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_7/_0_  (.A(net140),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[7] ));
 sky130_fd_sc_hd__buf_2 \NN4END_inbuf_8/_0_  (.A(net141),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \NN4END_inbuf_9/_0_  (.A(net142),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\NN4BEG_i[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_10 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_100 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_101 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_102 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_103 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_104 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_105 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_106 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_107 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_108 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_109 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_11 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_110 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_111 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_112 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_113 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_114 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_115 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_116 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_117 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_118 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_119 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_12 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_120 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_121 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_122 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_123 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_124 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_125 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_126 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_127 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_128 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_129 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_13 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_130 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_131 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_132 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_133 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_134 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_135 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_136 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_137 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_138 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_139 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_14 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_140 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_141 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_142 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_143 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_144 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_145 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_146 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_147 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_148 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_149 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_15 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_150 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_151 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_152 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_153 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_154 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_155 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_16 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_17 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_18 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_19 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_20 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_21 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_22 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_23 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_24 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_25 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_26 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_27 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_28 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_29 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_30 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_31 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_32 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_33 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_34 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_35 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_36 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_37 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_38 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_39 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_40 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_41 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_42 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_43 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_44 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_45 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_46 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_47 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_48 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_49 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_50 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_51 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_52 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_53 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_54 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_55 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_56 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_57 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_58 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_59 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_6 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_60 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_61 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_62 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_63 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_64 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_65 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_66 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_67 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_68 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_69 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_7 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_70 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_71 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_72 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_73 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_74 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_75 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_76 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_77 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_78 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_79 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_8 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_80 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_81 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_82 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_83 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_84 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_85 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_86 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_87 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_88 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_89 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_9 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_90 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_91 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_92 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_93 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_94 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_95 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_96 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_97 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_98 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__decap_3 PHY_99 (.VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_0/_0_  (.A(\S4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_1/_0_  (.A(\S4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_10/_0_  (.A(\S4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_11/_0_  (.A(\S4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_2/_0_  (.A(\S4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_3/_0_  (.A(\S4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_4/_0_  (.A(\S4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_5/_0_  (.A(\S4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_6/_0_  (.A(\S4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_7/_0_  (.A(\S4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_8/_0_  (.A(\S4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_9/_0_  (.A(\S4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net442));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_0/_0_  (.A(net184),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[0] ));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_1/_0_  (.A(net185),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_10/_0_  (.A(net179),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_11/_0_  (.A(net180),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[11] ));
 sky130_fd_sc_hd__buf_2 \S4END_inbuf_2/_0_  (.A(net186),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_3/_0_  (.A(net187),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_4/_0_  (.A(net188),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_5/_0_  (.A(net189),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_6/_0_  (.A(net175),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_7/_0_  (.A(net176),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_8/_0_  (.A(net177),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_9/_0_  (.A(net178),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\S4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_0/_0_  (.A(\SS4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_1/_0_  (.A(\SS4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_10/_0_  (.A(\SS4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_11/_0_  (.A(\SS4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_2/_0_  (.A(\SS4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_3/_0_  (.A(\SS4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_4/_0_  (.A(\SS4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_5/_0_  (.A(\SS4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_6/_0_  (.A(\SS4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_7/_0_  (.A(\SS4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_8/_0_  (.A(\SS4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 \SS4BEG_outbuf_9/_0_  (.A(\SS4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_0/_0_  (.A(net200),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_1/_0_  (.A(net201),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \SS4END_inbuf_10/_0_  (.A(net195),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[10] ));
 sky130_fd_sc_hd__buf_2 \SS4END_inbuf_11/_0_  (.A(net196),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_2/_0_  (.A(net202),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_3/_0_  (.A(net203),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_4/_0_  (.A(net204),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_5/_0_  (.A(net205),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_6/_0_  (.A(net191),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_7/_0_  (.A(net192),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_8/_0_  (.A(net193),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \SS4END_inbuf_9/_0_  (.A(net194),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\SS4BEG_i[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 (.VGND(vssd1),
    .VPWR(vccd1));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_0/_0_  (.A(\W6BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_1/_0_  (.A(\W6BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_2/_0_  (.A(\W6BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_3/_0_  (.A(\W6BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_4/_0_  (.A(\W6BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_5/_0_  (.A(\W6BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_6/_0_  (.A(\W6BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_7/_0_  (.A(\W6BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net489));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_8/_0_  (.A(\W6BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_1 \W6BEG_outbuf_9/_0_  (.A(\W6BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_0/_0_  (.A(net230),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_1/_0_  (.A(net231),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_2/_0_  (.A(net232),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_3/_0_  (.A(net233),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_4/_0_  (.A(net234),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_5/_0_  (.A(net235),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_6/_0_  (.A(net236),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_7/_0_  (.A(net237),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_8/_0_  (.A(net227),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \W6END_inbuf_9/_0_  (.A(net228),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\W6BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_0/_0_  (.A(\WW4BEG_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_1/_0_  (.A(\WW4BEG_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_10/_0_  (.A(\WW4BEG_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_11/_0_  (.A(\WW4BEG_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_2/_0_  (.A(\WW4BEG_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_3/_0_  (.A(\WW4BEG_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_4/_0_  (.A(\WW4BEG_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_5/_0_  (.A(\WW4BEG_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_6/_0_  (.A(\WW4BEG_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_7/_0_  (.A(\WW4BEG_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_8/_0_  (.A(\WW4BEG_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_1 \WW4BEG_outbuf_9/_0_  (.A(\WW4BEG_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net507));
 sky130_fd_sc_hd__buf_2 \WW4END_inbuf_0/_0_  (.A(net248),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_1/_0_  (.A(net249),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_10/_0_  (.A(net243),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_11/_0_  (.A(net244),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_2/_0_  (.A(net250),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_3/_0_  (.A(net251),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_4/_0_  (.A(net252),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_5/_0_  (.A(net253),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_6/_0_  (.A(net239),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_7/_0_  (.A(net240),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_8/_0_  (.A(net241),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \WW4END_inbuf_9/_0_  (.A(net242),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\WW4BEG_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0/_0_  (.A(net50),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1/_0_  (.A(net61),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10/_0_  (.A(net51),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11/_0_  (.A(net52),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12/_0_  (.A(net53),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13/_0_  (.A(net54),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14/_0_  (.A(net55),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15/_0_  (.A(net56),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16/_0_  (.A(net57),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17/_0_  (.A(net58),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18/_0_  (.A(net59),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19/_0_  (.A(net60),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2/_0_  (.A(net72),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20/_0_  (.A(net62),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21/_0_  (.A(net63),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22/_0_  (.A(net64),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23/_0_  (.A(net65),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24/_0_  (.A(net66),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25/_0_  (.A(net67),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26/_0_  (.A(net68),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27/_0_  (.A(net69),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28/_0_  (.A(net70),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29/_0_  (.A(net71),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3/_0_  (.A(net75),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30/_0_  (.A(net73),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31/_0_  (.A(net74),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4/_0_  (.A(net76),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5/_0_  (.A(net77),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6/_0_  (.A(net78),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7/_0_  (.A(net79),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8/_0_  (.A(net80),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9/_0_  (.A(net81),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0/_0_  (.A(\FrameData_O_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1/_0_  (.A(\FrameData_O_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10/_0_  (.A(\FrameData_O_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11/_0_  (.A(\FrameData_O_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12/_0_  (.A(\FrameData_O_i[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13/_0_  (.A(\FrameData_O_i[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14/_0_  (.A(\FrameData_O_i[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15/_0_  (.A(\FrameData_O_i[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16/_0_  (.A(\FrameData_O_i[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17/_0_  (.A(\FrameData_O_i[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18/_0_  (.A(\FrameData_O_i[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19/_0_  (.A(\FrameData_O_i[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2/_0_  (.A(\FrameData_O_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20/_0_  (.A(\FrameData_O_i[20] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21/_0_  (.A(\FrameData_O_i[21] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22/_0_  (.A(\FrameData_O_i[22] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23/_0_  (.A(\FrameData_O_i[23] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24/_0_  (.A(\FrameData_O_i[24] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25/_0_  (.A(\FrameData_O_i[25] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26/_0_  (.A(\FrameData_O_i[26] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27/_0_  (.A(\FrameData_O_i[27] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28/_0_  (.A(\FrameData_O_i[28] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29/_0_  (.A(\FrameData_O_i[29] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3/_0_  (.A(\FrameData_O_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30/_0_  (.A(\FrameData_O_i[30] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31/_0_  (.A(\FrameData_O_i[31] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4/_0_  (.A(\FrameData_O_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5/_0_  (.A(\FrameData_O_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6/_0_  (.A(\FrameData_O_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7/_0_  (.A(\FrameData_O_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8/_0_  (.A(\FrameData_O_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9/_0_  (.A(\FrameData_O_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\Inst_LE_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\Inst_LH_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\Inst_LB_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\Inst_LG_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\Inst_LF_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\Inst_LC_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\Inst_LD_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\Inst_LA_LUT4c_frame_config_dffesr/LUT_flop ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(Ci),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(E2END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net10));
 sky130_fd_sc_hd__buf_12 input100 (.A(FrameStrobe[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_16 input101 (.A(FrameStrobe[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 input102 (.A(N1END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net102));
 sky130_fd_sc_hd__buf_4 input103 (.A(N1END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net103));
 sky130_fd_sc_hd__buf_4 input104 (.A(N1END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net104));
 sky130_fd_sc_hd__buf_4 input105 (.A(N1END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 input106 (.A(N2END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(N2END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(N2END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net108));
 sky130_fd_sc_hd__buf_2 input109 (.A(N2END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net109));
 sky130_fd_sc_hd__buf_2 input11 (.A(E2END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input110 (.A(N2END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net110));
 sky130_fd_sc_hd__buf_2 input111 (.A(N2END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(N2END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 input113 (.A(N2END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 input114 (.A(N2MID[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 input115 (.A(N2MID[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_4 input116 (.A(N2MID[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(N2MID[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net117));
 sky130_fd_sc_hd__buf_2 input118 (.A(N2MID[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 input119 (.A(N2MID[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net119));
 sky130_fd_sc_hd__buf_2 input12 (.A(E2END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input120 (.A(N2MID[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 input121 (.A(N2MID[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net121));
 sky130_fd_sc_hd__buf_2 input122 (.A(N4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(N4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(N4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(N4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(N4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(N4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(N4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(N4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net129));
 sky130_fd_sc_hd__buf_2 input13 (.A(E2END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input130 (.A(N4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(N4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(N4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(N4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(N4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(N4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(N4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(N4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net137));
 sky130_fd_sc_hd__dlymetal6s2s_1 input138 (.A(NN4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(NN4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(E2MID[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(NN4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(NN4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 input142 (.A(NN4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(NN4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(NN4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net144));
 sky130_fd_sc_hd__dlymetal6s2s_1 input145 (.A(NN4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(NN4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 input147 (.A(NN4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(NN4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 input149 (.A(NN4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(E2MID[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(NN4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(NN4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(NN4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 input153 (.A(NN4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(S1END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(S1END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(S1END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(S1END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(S2END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(S2END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net159));
 sky130_fd_sc_hd__buf_2 input16 (.A(E2MID[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input160 (.A(S2END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(S2END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(S2END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net162));
 sky130_fd_sc_hd__buf_2 input163 (.A(S2END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(S2END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(S2END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(S2MID[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(S2MID[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(S2MID[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net168));
 sky130_fd_sc_hd__buf_4 input169 (.A(S2MID[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input170 (.A(S2MID[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(S2MID[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(S2MID[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(S2MID[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net173));
 sky130_fd_sc_hd__buf_2 input174 (.A(S4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(S4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(S4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(S4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(S4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(S4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(E2MID[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(S4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net180));
 sky130_fd_sc_hd__buf_2 input181 (.A(S4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(S4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net182));
 sky130_fd_sc_hd__buf_2 input183 (.A(S4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(S4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(S4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(S4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(S4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(S4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 input189 (.A(S4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input19 (.A(E2MID[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(SS4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 input191 (.A(SS4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(SS4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(SS4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(SS4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(SS4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(SS4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(SS4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 input198 (.A(SS4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net198));
 sky130_fd_sc_hd__dlymetal6s2s_1 input199 (.A(SS4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net199));
 sky130_fd_sc_hd__buf_4 input2 (.A(E1END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(E2MID[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(SS4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(SS4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(SS4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(SS4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(SS4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(SS4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net205));
 sky130_fd_sc_hd__buf_4 input206 (.A(W1END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net206));
 sky130_fd_sc_hd__buf_4 input207 (.A(W1END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net207));
 sky130_fd_sc_hd__buf_4 input208 (.A(W1END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net208));
 sky130_fd_sc_hd__buf_4 input209 (.A(W1END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net209));
 sky130_fd_sc_hd__buf_2 input21 (.A(E2MID[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(W2END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net210));
 sky130_fd_sc_hd__buf_2 input211 (.A(W2END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net211));
 sky130_fd_sc_hd__buf_2 input212 (.A(W2END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net212));
 sky130_fd_sc_hd__buf_2 input213 (.A(W2END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net213));
 sky130_fd_sc_hd__buf_2 input214 (.A(W2END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 input215 (.A(W2END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 input216 (.A(W2END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_2 input217 (.A(W2END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net217));
 sky130_fd_sc_hd__buf_2 input218 (.A(W2MID[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 input219 (.A(W2MID[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net219));
 sky130_fd_sc_hd__buf_4 input22 (.A(E6END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input220 (.A(W2MID[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net220));
 sky130_fd_sc_hd__buf_2 input221 (.A(W2MID[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net221));
 sky130_fd_sc_hd__buf_2 input222 (.A(W2MID[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(W2MID[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 input224 (.A(W2MID[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 input225 (.A(W2MID[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 input226 (.A(W6END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(W6END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(W6END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net228));
 sky130_fd_sc_hd__buf_4 input229 (.A(W6END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(E6END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input230 (.A(W6END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(W6END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(W6END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 input233 (.A(W6END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(W6END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(W6END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(W6END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(W6END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 input238 (.A(WW4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(WW4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(E6END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(WW4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(WW4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(WW4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(WW4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(WW4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 input245 (.A(WW4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(WW4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net246));
 sky130_fd_sc_hd__dlymetal6s2s_1 input247 (.A(WW4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 input248 (.A(WW4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 input249 (.A(WW4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net249));
 sky130_fd_sc_hd__buf_4 input25 (.A(E6END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input250 (.A(WW4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(WW4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 input252 (.A(WW4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 input253 (.A(WW4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(E6END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(E6END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(E6END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(E6END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(E1END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(E6END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(E6END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(E6END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(E6END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(EE4END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(EE4END[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(EE4END[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(EE4END[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(EE4END[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(EE4END[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(E1END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(EE4END[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(EE4END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(EE4END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net42));
 sky130_fd_sc_hd__buf_2 input43 (.A(EE4END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(EE4END[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(EE4END[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(EE4END[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(EE4END[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(EE4END[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(EE4END[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net49));
 sky130_fd_sc_hd__buf_4 input5 (.A(E1END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net5));
 sky130_fd_sc_hd__buf_6 input50 (.A(FrameData[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net50));
 sky130_fd_sc_hd__buf_8 input51 (.A(FrameData[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net51));
 sky130_fd_sc_hd__buf_8 input52 (.A(FrameData[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net52));
 sky130_fd_sc_hd__buf_8 input53 (.A(FrameData[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net53));
 sky130_fd_sc_hd__buf_8 input54 (.A(FrameData[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net54));
 sky130_fd_sc_hd__buf_8 input55 (.A(FrameData[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net55));
 sky130_fd_sc_hd__buf_8 input56 (.A(FrameData[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net56));
 sky130_fd_sc_hd__buf_8 input57 (.A(FrameData[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net57));
 sky130_fd_sc_hd__buf_8 input58 (.A(FrameData[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net58));
 sky130_fd_sc_hd__buf_8 input59 (.A(FrameData[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net6));
 sky130_fd_sc_hd__buf_8 input60 (.A(FrameData[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(FrameData[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net61));
 sky130_fd_sc_hd__buf_8 input62 (.A(FrameData[20]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net62));
 sky130_fd_sc_hd__buf_8 input63 (.A(FrameData[21]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net63));
 sky130_fd_sc_hd__buf_8 input64 (.A(FrameData[22]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net64));
 sky130_fd_sc_hd__buf_8 input65 (.A(FrameData[23]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_16 input66 (.A(FrameData[24]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net66));
 sky130_fd_sc_hd__buf_8 input67 (.A(FrameData[25]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net67));
 sky130_fd_sc_hd__buf_8 input68 (.A(FrameData[26]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net68));
 sky130_fd_sc_hd__buf_8 input69 (.A(FrameData[27]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(E2END[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net7));
 sky130_fd_sc_hd__buf_8 input70 (.A(FrameData[28]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net70));
 sky130_fd_sc_hd__buf_8 input71 (.A(FrameData[29]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net71));
 sky130_fd_sc_hd__buf_8 input72 (.A(FrameData[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net72));
 sky130_fd_sc_hd__buf_8 input73 (.A(FrameData[30]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net73));
 sky130_fd_sc_hd__buf_8 input74 (.A(FrameData[31]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net74));
 sky130_fd_sc_hd__buf_8 input75 (.A(FrameData[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net75));
 sky130_fd_sc_hd__buf_8 input76 (.A(FrameData[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_16 input77 (.A(FrameData[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net77));
 sky130_fd_sc_hd__buf_8 input78 (.A(FrameData[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net78));
 sky130_fd_sc_hd__buf_8 input79 (.A(FrameData[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(E2END[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net8));
 sky130_fd_sc_hd__buf_8 input80 (.A(FrameData[8]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net80));
 sky130_fd_sc_hd__buf_8 input81 (.A(FrameData[9]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net81));
 sky130_fd_sc_hd__buf_8 input82 (.A(FrameStrobe[0]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net82));
 sky130_fd_sc_hd__buf_12 input83 (.A(FrameStrobe[10]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_16 input84 (.A(FrameStrobe[11]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net84));
 sky130_fd_sc_hd__buf_8 input85 (.A(FrameStrobe[12]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_16 input86 (.A(FrameStrobe[13]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net86));
 sky130_fd_sc_hd__buf_8 input87 (.A(FrameStrobe[14]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net87));
 sky130_fd_sc_hd__buf_8 input88 (.A(FrameStrobe[15]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net88));
 sky130_fd_sc_hd__buf_8 input89 (.A(FrameStrobe[16]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net89));
 sky130_fd_sc_hd__buf_2 input9 (.A(E2END[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net9));
 sky130_fd_sc_hd__buf_8 input90 (.A(FrameStrobe[17]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net90));
 sky130_fd_sc_hd__buf_8 input91 (.A(FrameStrobe[18]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net91));
 sky130_fd_sc_hd__buf_8 input92 (.A(FrameStrobe[19]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_16 input93 (.A(FrameStrobe[1]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_16 input94 (.A(FrameStrobe[2]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 input95 (.A(FrameStrobe[3]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_16 input96 (.A(FrameStrobe[4]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 input97 (.A(FrameStrobe[5]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 input98 (.A(FrameStrobe[6]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_16 input99 (.A(FrameStrobe[7]),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(Co));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E1BEG[0]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E1BEG[1]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[2]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net262),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output265 (.A(net265),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[6]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEG[7]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[4]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E2BEGb[7]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[0]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[5]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(E6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output288 (.A(net288),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[10]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[12]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output292 (.A(net292),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[15]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output296 (.A(net296),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output298 (.A(net298),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[6]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net300),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output301 (.A(net301),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output302 (.A(net302),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(EE4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output305 (.A(net305),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output306 (.A(net306),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net312),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output313 (.A(net313),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__clkbuf_4 output316 (.A(net316),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net317),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net319),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output322 (.A(net322),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output324 (.A(net324),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output327 (.A(net327),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__clkbuf_4 output328 (.A(net328),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output339 (.A(net339),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output345 (.A(net345),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net365),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output368 (.A(net368),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output369 (.A(net369),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output392 (.A(net392),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[11]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output395 (.A(net395),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[13]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output397 (.A(net397),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output398 (.A(net398),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output399 (.A(net399),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[2]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output401 (.A(net401),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output402 (.A(net402),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output403 (.A(net403),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output404 (.A(net404),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[7]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output406 (.A(net406),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(NN4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output407 (.A(net407),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output408 (.A(net408),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output409 (.A(net409),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__buf_2 output410 (.A(net410),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output412 (.A(net412),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output413 (.A(net413),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output416 (.A(net416),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output417 (.A(net417),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output418 (.A(net418),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__buf_2 output419 (.A(net419),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output420 (.A(net420),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output421 (.A(net421),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output422 (.A(net422),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output423 (.A(net423),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output424 (.A(net424),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output425 (.A(net425),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output426 (.A(net426),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output427 (.A(net427),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output428 (.A(net428),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output429 (.A(net429),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output430 (.A(net430),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output431 (.A(net431),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output432 (.A(net432),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__buf_2 output433 (.A(net433),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output434 (.A(net434),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output435 (.A(net435),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output436 (.A(net436),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output437 (.A(net437),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output438 (.A(net438),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__buf_2 output439 (.A(net439),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output440 (.A(net440),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output441 (.A(net441),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output442 (.A(net442),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output443 (.A(net443),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output444 (.A(net444),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output445 (.A(net445),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output446 (.A(net446),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output447 (.A(net447),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output448 (.A(net448),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output449 (.A(net449),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output450 (.A(net450),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output451 (.A(net451),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output452 (.A(net452),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output453 (.A(net453),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output454 (.A(net454),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output455 (.A(net455),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output456 (.A(net456),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output457 (.A(net457),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output458 (.A(net458),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(SS4BEG[9]));
 sky130_fd_sc_hd__buf_1 output459 (.A(net459),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(UserCLKo));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output461 (.A(net461),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__buf_2 output463 (.A(net463),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output470 (.A(net470),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__buf_2 output472 (.A(net472),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output473 (.A(net473),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net475),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output476 (.A(net476),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output477 (.A(net477),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net478),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net479),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output480 (.A(net480),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net481),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output482 (.A(net482),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output483 (.A(net483),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net484),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output485 (.A(net485),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net487),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output488 (.A(net488),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output489 (.A(net489),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output490 (.A(net490),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output491 (.A(net491),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output493 (.A(net493),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net494),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output495 (.A(net495),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net497),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output499 (.A(net499),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net503),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__buf_2 output504 (.A(net504),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__buf_2 output505 (.A(net505),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__buf_2 output506 (.A(net506),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0/_0_  (.A(net82),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1/_0_  (.A(net93),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_10/_0_  (.A(net83),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_11/_0_  (.A(net84),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_12/_0_  (.A(net85),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_13/_0_  (.A(net86),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_14/_0_  (.A(net87),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_15/_0_  (.A(net88),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_16/_0_  (.A(net89),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_17/_0_  (.A(net90),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_18/_0_  (.A(net91),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_19/_0_  (.A(net92),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2/_0_  (.A(net94),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3/_0_  (.A(net95),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4/_0_  (.A(net96),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_5/_0_  (.A(net97),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6/_0_  (.A(net98),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_7/_0_  (.A(net99),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_8/_0_  (.A(net100),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_9/_0_  (.A(net101),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(\FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0/_0_  (.A(\FrameStrobe_O_i[0] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1/_0_  (.A(\FrameStrobe_O_i[1] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10/_0_  (.A(\FrameStrobe_O_i[10] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11/_0_  (.A(\FrameStrobe_O_i[11] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12/_0_  (.A(\FrameStrobe_O_i[12] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13/_0_  (.A(\FrameStrobe_O_i[13] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14/_0_  (.A(\FrameStrobe_O_i[14] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15/_0_  (.A(\FrameStrobe_O_i[15] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16/_0_  (.A(\FrameStrobe_O_i[16] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17/_0_  (.A(\FrameStrobe_O_i[17] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_18/_0_  (.A(\FrameStrobe_O_i[18] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19/_0_  (.A(\FrameStrobe_O_i[19] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2/_0_  (.A(\FrameStrobe_O_i[2] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3/_0_  (.A(\FrameStrobe_O_i[3] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4/_0_  (.A(\FrameStrobe_O_i[4] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5/_0_  (.A(\FrameStrobe_O_i[5] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6/_0_  (.A(\FrameStrobe_O_i[6] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7/_0_  (.A(\FrameStrobe_O_i[7] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8/_0_  (.A(\FrameStrobe_O_i[8] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9/_0_  (.A(\FrameStrobe_O_i[9] ),
    .VGND(vssd1),
    .VNB(vssd1),
    .VPB(vccd1),
    .VPWR(vccd1),
    .X(net354));
endmodule
