magic
tech sky130A
magscale 1 2
timestamp 1732489415
<< viali >>
rect 1593 6409 1627 6443
rect 2421 6409 2455 6443
rect 4169 6409 4203 6443
rect 4629 6409 4663 6443
rect 6377 6409 6411 6443
rect 7205 6409 7239 6443
rect 7389 6409 7423 6443
rect 8401 6409 8435 6443
rect 8585 6409 8619 6443
rect 9413 6409 9447 6443
rect 9781 6409 9815 6443
rect 10609 6409 10643 6443
rect 10977 6409 11011 6443
rect 11989 6409 12023 6443
rect 12173 6409 12207 6443
rect 12449 6409 12483 6443
rect 13185 6409 13219 6443
rect 13369 6409 13403 6443
rect 14289 6409 14323 6443
rect 14933 6409 14967 6443
rect 15393 6409 15427 6443
rect 15761 6409 15795 6443
rect 16865 6409 16899 6443
rect 17233 6409 17267 6443
rect 17969 6409 18003 6443
rect 18153 6409 18187 6443
rect 19441 6409 19475 6443
rect 19809 6409 19843 6443
rect 20361 6409 20395 6443
rect 20821 6409 20855 6443
rect 21557 6409 21591 6443
rect 21833 6409 21867 6443
rect 22569 6409 22603 6443
rect 22937 6409 22971 6443
rect 23489 6409 23523 6443
rect 23949 6409 23983 6443
rect 5733 6341 5767 6375
rect 6101 6341 6135 6375
rect 6929 6341 6963 6375
rect 8125 6341 8159 6375
rect 9321 6341 9355 6375
rect 10517 6341 10551 6375
rect 14197 6341 14231 6375
rect 15301 6341 15335 6375
rect 16773 6341 16807 6375
rect 17693 6341 17727 6375
rect 19349 6341 19383 6375
rect 22477 6341 22511 6375
rect 23857 6341 23891 6375
rect 1501 6273 1535 6307
rect 2237 6273 2271 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 6561 6273 6595 6307
rect 7573 6273 7607 6307
rect 8769 6273 8803 6307
rect 9965 6273 9999 6307
rect 11161 6273 11195 6307
rect 11805 6273 11839 6307
rect 12357 6273 12391 6307
rect 12633 6273 12667 6307
rect 13001 6273 13035 6307
rect 13553 6273 13587 6307
rect 14657 6273 14691 6307
rect 15117 6273 15151 6307
rect 15945 6273 15979 6307
rect 17417 6273 17451 6307
rect 18337 6273 18371 6307
rect 19993 6273 20027 6307
rect 20177 6273 20211 6307
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 21373 6273 21407 6307
rect 22017 6273 22051 6307
rect 23121 6273 23155 6307
rect 23673 6273 23707 6307
rect 20729 6137 20763 6171
rect 14841 6069 14875 6103
rect 6101 5865 6135 5899
rect 7389 5865 7423 5899
rect 8585 5865 8619 5899
rect 9689 5865 9723 5899
rect 10885 5865 10919 5899
rect 12265 5865 12299 5899
rect 13277 5865 13311 5899
rect 14381 5865 14415 5899
rect 15761 5865 15795 5899
rect 16957 5865 16991 5899
rect 18245 5865 18279 5899
rect 19809 5865 19843 5899
rect 24133 5865 24167 5899
rect 11805 5797 11839 5831
rect 6285 5661 6319 5695
rect 7573 5661 7607 5695
rect 8769 5661 8803 5695
rect 9873 5661 9907 5695
rect 11069 5661 11103 5695
rect 11989 5661 12023 5695
rect 12449 5661 12483 5695
rect 13461 5661 13495 5695
rect 14565 5661 14599 5695
rect 14841 5661 14875 5695
rect 15945 5661 15979 5695
rect 17141 5661 17175 5695
rect 18429 5661 18463 5695
rect 19993 5661 20027 5695
rect 23857 5593 23891 5627
rect 14657 5525 14691 5559
rect 6377 5321 6411 5355
rect 7573 5321 7607 5355
rect 8769 5321 8803 5355
rect 9873 5321 9907 5355
rect 11069 5321 11103 5355
rect 11989 5321 12023 5355
rect 12449 5321 12483 5355
rect 13461 5321 13495 5355
rect 14565 5321 14599 5355
rect 14841 5321 14875 5355
rect 15945 5321 15979 5355
rect 17141 5321 17175 5355
rect 18429 5321 18463 5355
rect 19993 5321 20027 5355
rect 24133 5321 24167 5355
rect 6561 5185 6595 5219
rect 7297 5185 7331 5219
rect 7757 5185 7791 5219
rect 8953 5185 8987 5219
rect 10057 5185 10091 5219
rect 11253 5185 11287 5219
rect 12173 5185 12207 5219
rect 12633 5185 12667 5219
rect 13645 5185 13679 5219
rect 14749 5185 14783 5219
rect 15025 5185 15059 5219
rect 16129 5185 16163 5219
rect 17325 5185 17359 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 24317 5185 24351 5219
rect 6929 4981 6963 5015
rect 24041 4777 24075 4811
rect 23949 4573 23983 4607
rect 24225 4573 24259 4607
rect 23765 4437 23799 4471
rect 23949 3689 23983 3723
rect 24133 3485 24167 3519
rect 24133 3145 24167 3179
rect 23489 3009 23523 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 24317 3009 24351 3043
rect 23305 2805 23339 2839
rect 23581 2805 23615 2839
rect 23857 2805 23891 2839
rect 1685 2601 1719 2635
rect 16313 2601 16347 2635
rect 22569 2601 22603 2635
rect 22937 2601 22971 2635
rect 23213 2601 23247 2635
rect 23765 2601 23799 2635
rect 1593 2533 1627 2567
rect 1961 2533 1995 2567
rect 15117 2533 15151 2567
rect 16589 2533 16623 2567
rect 23489 2533 23523 2567
rect 1409 2397 1443 2431
rect 1869 2397 1903 2431
rect 2145 2397 2179 2431
rect 2237 2397 2271 2431
rect 4905 2397 4939 2431
rect 6101 2397 6135 2431
rect 7389 2397 7423 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 10425 2397 10459 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 12817 2397 12851 2431
rect 13277 2397 13311 2431
rect 15301 2393 15335 2427
rect 15577 2397 15611 2431
rect 15945 2397 15979 2431
rect 16497 2397 16531 2431
rect 16773 2397 16807 2431
rect 17049 2397 17083 2431
rect 17325 2397 17359 2431
rect 17601 2397 17635 2431
rect 17877 2397 17911 2431
rect 18153 2397 18187 2431
rect 18429 2397 18463 2431
rect 18705 2397 18739 2431
rect 18981 2397 19015 2431
rect 19441 2397 19475 2431
rect 19717 2397 19751 2431
rect 19993 2397 20027 2431
rect 20269 2397 20303 2431
rect 20545 2397 20579 2431
rect 20821 2397 20855 2431
rect 22385 2397 22419 2431
rect 22845 2397 22879 2431
rect 23121 2397 23155 2431
rect 23397 2397 23431 2431
rect 23673 2397 23707 2431
rect 23949 2397 23983 2431
rect 24225 2397 24259 2431
rect 2421 2261 2455 2295
rect 4721 2261 4755 2295
rect 6285 2261 6319 2295
rect 7205 2261 7239 2295
rect 9413 2261 9447 2295
rect 9689 2261 9723 2295
rect 10241 2261 10275 2295
rect 10977 2261 11011 2295
rect 11529 2261 11563 2295
rect 11805 2261 11839 2295
rect 12081 2261 12115 2295
rect 12357 2261 12391 2295
rect 12633 2261 12667 2295
rect 13093 2261 13127 2295
rect 15393 2261 15427 2295
rect 16129 2261 16163 2295
rect 16865 2261 16899 2295
rect 17141 2261 17175 2295
rect 17417 2261 17451 2295
rect 17693 2261 17727 2295
rect 17969 2261 18003 2295
rect 18245 2261 18279 2295
rect 18521 2261 18555 2295
rect 18797 2261 18831 2295
rect 19257 2261 19291 2295
rect 19533 2261 19567 2295
rect 19809 2261 19843 2295
rect 20085 2261 20119 2295
rect 20361 2261 20395 2295
rect 20637 2261 20671 2295
rect 22661 2261 22695 2295
rect 24041 2261 24075 2295
rect 2421 2057 2455 2091
rect 2697 2057 2731 2091
rect 7573 2057 7607 2091
rect 7849 2057 7883 2091
rect 8125 2057 8159 2091
rect 13553 2057 13587 2091
rect 14197 2057 14231 2091
rect 17417 2057 17451 2091
rect 17693 2057 17727 2091
rect 21465 2057 21499 2091
rect 21833 2057 21867 2091
rect 22293 2057 22327 2091
rect 22753 2057 22787 2091
rect 24409 2057 24443 2091
rect 10425 1989 10459 2023
rect 10977 1989 11011 2023
rect 11989 1989 12023 2023
rect 12817 1989 12851 2023
rect 15853 1989 15887 2023
rect 18061 1989 18095 2023
rect 18613 1989 18647 2023
rect 19717 1989 19751 2023
rect 20821 1989 20855 2023
rect 1685 1921 1719 1955
rect 1777 1921 1811 1955
rect 2145 1921 2179 1955
rect 2605 1921 2639 1955
rect 2881 1921 2915 1955
rect 3157 1921 3191 1955
rect 3433 1921 3467 1955
rect 3709 1921 3743 1955
rect 3985 1921 4019 1955
rect 4261 1921 4295 1955
rect 4537 1921 4571 1955
rect 4813 1921 4847 1955
rect 5089 1921 5123 1955
rect 5365 1921 5399 1955
rect 5641 1921 5675 1955
rect 5733 1921 5767 1955
rect 6193 1921 6227 1955
rect 6653 1921 6687 1955
rect 6929 1921 6963 1955
rect 7021 1921 7055 1955
rect 7481 1921 7515 1955
rect 7757 1921 7791 1955
rect 8033 1921 8067 1955
rect 8309 1921 8343 1955
rect 8585 1921 8619 1955
rect 8861 1921 8895 1955
rect 9137 1921 9171 1955
rect 9405 1921 9439 1955
rect 9689 1921 9723 1955
rect 9965 1921 9999 1955
rect 10241 1921 10275 1955
rect 11529 1921 11563 1955
rect 12633 1921 12667 1955
rect 13461 1921 13495 1955
rect 13737 1921 13771 1955
rect 14105 1921 14139 1955
rect 14381 1921 14415 1955
rect 14473 1921 14507 1955
rect 14841 1921 14875 1955
rect 15393 1921 15427 1955
rect 15669 1921 15703 1955
rect 16497 1921 16531 1955
rect 16957 1921 16991 1955
rect 17601 1921 17635 1955
rect 17877 1921 17911 1955
rect 19165 1921 19199 1955
rect 20269 1921 20303 1955
rect 21097 1921 21131 1955
rect 21649 1921 21683 1955
rect 22017 1921 22051 1955
rect 22109 1921 22143 1955
rect 22661 1921 22695 1955
rect 22937 1921 22971 1955
rect 23029 1921 23063 1955
rect 23581 1921 23615 1955
rect 23857 1921 23891 1955
rect 24133 1921 24167 1955
rect 24225 1921 24259 1955
rect 3525 1785 3559 1819
rect 3801 1785 3835 1819
rect 4629 1785 4663 1819
rect 4905 1785 4939 1819
rect 5917 1785 5951 1819
rect 7205 1785 7239 1819
rect 8953 1785 8987 1819
rect 9505 1785 9539 1819
rect 10057 1785 10091 1819
rect 15209 1785 15243 1819
rect 22477 1785 22511 1819
rect 23397 1785 23431 1819
rect 23949 1785 23983 1819
rect 1501 1717 1535 1751
rect 1961 1717 1995 1751
rect 2329 1717 2363 1751
rect 2973 1717 3007 1751
rect 3249 1717 3283 1751
rect 4077 1717 4111 1751
rect 4353 1717 4387 1751
rect 5181 1717 5215 1751
rect 5457 1717 5491 1751
rect 6009 1717 6043 1751
rect 6469 1717 6503 1751
rect 6745 1717 6779 1751
rect 7297 1717 7331 1751
rect 8401 1717 8435 1751
rect 8677 1717 8711 1751
rect 9229 1717 9263 1751
rect 9781 1717 9815 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11713 1717 11747 1751
rect 12081 1717 12115 1751
rect 12449 1717 12483 1751
rect 12909 1717 12943 1751
rect 13277 1717 13311 1751
rect 13921 1717 13955 1751
rect 14657 1717 14691 1751
rect 15025 1717 15059 1751
rect 15485 1717 15519 1751
rect 15945 1717 15979 1751
rect 16313 1717 16347 1751
rect 17049 1717 17083 1751
rect 18153 1717 18187 1751
rect 18705 1717 18739 1751
rect 19257 1717 19291 1751
rect 19809 1717 19843 1751
rect 20361 1717 20395 1751
rect 20913 1717 20947 1751
rect 21281 1717 21315 1751
rect 23213 1717 23247 1751
rect 23673 1717 23707 1751
rect 2605 1513 2639 1547
rect 2881 1513 2915 1547
rect 5089 1513 5123 1547
rect 6193 1513 6227 1547
rect 14289 1513 14323 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 18521 1513 18555 1547
rect 19441 1513 19475 1547
rect 21097 1513 21131 1547
rect 21465 1513 21499 1547
rect 23213 1513 23247 1547
rect 3433 1445 3467 1479
rect 6653 1445 6687 1479
rect 7205 1445 7239 1479
rect 7481 1445 7515 1479
rect 8585 1445 8619 1479
rect 20085 1445 20119 1479
rect 20637 1445 20671 1479
rect 21833 1445 21867 1479
rect 11069 1377 11103 1411
rect 1685 1309 1719 1343
rect 1777 1309 1811 1343
rect 2237 1309 2271 1343
rect 2513 1309 2547 1343
rect 2789 1309 2823 1343
rect 3065 1309 3099 1343
rect 3341 1309 3375 1343
rect 3617 1309 3651 1343
rect 3985 1309 4019 1343
rect 4261 1309 4295 1343
rect 4537 1309 4571 1343
rect 4629 1309 4663 1343
rect 4905 1309 4939 1343
rect 5365 1309 5399 1343
rect 5641 1309 5675 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6561 1309 6595 1343
rect 6837 1309 6871 1343
rect 7113 1309 7147 1343
rect 7389 1309 7423 1343
rect 7665 1309 7699 1343
rect 7941 1309 7975 1343
rect 8217 1309 8251 1343
rect 8493 1309 8527 1343
rect 8769 1285 8803 1319
rect 9045 1309 9079 1343
rect 9505 1309 9539 1343
rect 9597 1309 9631 1343
rect 9965 1309 9999 1343
rect 10333 1309 10367 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12909 1309 12943 1343
rect 13277 1309 13311 1343
rect 14197 1309 14231 1343
rect 14657 1309 14691 1343
rect 15301 1309 15335 1343
rect 15853 1309 15887 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 17877 1309 17911 1343
rect 19073 1309 19107 1343
rect 19901 1309 19935 1343
rect 21005 1309 21039 1343
rect 21649 1309 21683 1343
rect 22017 1309 22051 1343
rect 22109 1309 22143 1343
rect 22385 1309 22419 1343
rect 22661 1309 22695 1343
rect 22937 1309 22971 1343
rect 23397 1309 23431 1343
rect 23489 1309 23523 1343
rect 23765 1309 23799 1343
rect 24041 1309 24075 1343
rect 10793 1241 10827 1275
rect 12265 1241 12299 1275
rect 17325 1241 17359 1275
rect 18429 1241 18463 1275
rect 19349 1241 19383 1275
rect 20453 1241 20487 1275
rect 1501 1173 1535 1207
rect 1961 1173 1995 1207
rect 2053 1173 2087 1207
rect 2329 1173 2363 1207
rect 3157 1173 3191 1207
rect 3801 1173 3835 1207
rect 4077 1173 4111 1207
rect 4353 1173 4387 1207
rect 4813 1173 4847 1207
rect 5181 1173 5215 1207
rect 5457 1173 5491 1207
rect 5917 1173 5951 1207
rect 6377 1173 6411 1207
rect 6929 1173 6963 1207
rect 7757 1173 7791 1207
rect 8033 1173 8067 1207
rect 8309 1173 8343 1207
rect 9229 1173 9263 1207
rect 9321 1173 9355 1207
rect 9781 1173 9815 1207
rect 10149 1173 10183 1207
rect 10517 1173 10551 1207
rect 11529 1173 11563 1207
rect 11989 1173 12023 1207
rect 12357 1173 12391 1207
rect 13093 1173 13127 1207
rect 13461 1173 13495 1207
rect 14841 1173 14875 1207
rect 17969 1173 18003 1207
rect 18889 1173 18923 1207
rect 22293 1173 22327 1207
rect 22569 1173 22603 1207
rect 22845 1173 22879 1207
rect 23121 1173 23155 1207
rect 23673 1173 23707 1207
rect 23949 1173 23983 1207
rect 24225 1173 24259 1207
<< metal1 >>
rect 1104 6554 25000 6576
rect 1104 6502 6884 6554
rect 6936 6502 6948 6554
rect 7000 6502 7012 6554
rect 7064 6502 7076 6554
rect 7128 6502 7140 6554
rect 7192 6502 12818 6554
rect 12870 6502 12882 6554
rect 12934 6502 12946 6554
rect 12998 6502 13010 6554
rect 13062 6502 13074 6554
rect 13126 6502 18752 6554
rect 18804 6502 18816 6554
rect 18868 6502 18880 6554
rect 18932 6502 18944 6554
rect 18996 6502 19008 6554
rect 19060 6502 24686 6554
rect 24738 6502 24750 6554
rect 24802 6502 24814 6554
rect 24866 6502 24878 6554
rect 24930 6502 24942 6554
rect 24994 6502 25000 6554
rect 1104 6480 25000 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1360 6412 1593 6440
rect 1360 6400 1366 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 2188 6412 2421 6440
rect 2188 6400 2194 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 2409 6403 2467 6409
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 3844 6412 4169 6440
rect 3844 6400 3850 6412
rect 4157 6409 4169 6412
rect 4203 6409 4215 6443
rect 4157 6403 4215 6409
rect 4614 6400 4620 6452
rect 4672 6400 4678 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 5736 6412 6377 6440
rect 5626 6372 5632 6384
rect 2240 6344 5632 6372
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 2240 6313 2268 6344
rect 5626 6332 5632 6344
rect 5684 6332 5690 6384
rect 5736 6381 5764 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7282 6440 7288 6452
rect 7239 6412 7288 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6409 7435 6443
rect 7377 6403 7435 6409
rect 5721 6375 5779 6381
rect 5721 6341 5733 6375
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 6086 6332 6092 6384
rect 6144 6332 6150 6384
rect 6917 6375 6975 6381
rect 6917 6341 6929 6375
rect 6963 6372 6975 6375
rect 7392 6372 7420 6403
rect 8386 6400 8392 6452
rect 8444 6400 8450 6452
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6409 8631 6443
rect 8573 6403 8631 6409
rect 6963 6344 7420 6372
rect 8113 6375 8171 6381
rect 6963 6341 6975 6344
rect 6917 6335 6975 6341
rect 8113 6341 8125 6375
rect 8159 6372 8171 6375
rect 8588 6372 8616 6403
rect 9398 6400 9404 6452
rect 9456 6400 9462 6452
rect 9769 6443 9827 6449
rect 9769 6409 9781 6443
rect 9815 6409 9827 6443
rect 9769 6403 9827 6409
rect 8159 6344 8616 6372
rect 9309 6375 9367 6381
rect 8159 6341 8171 6344
rect 8113 6335 8171 6341
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9784 6372 9812 6403
rect 10594 6400 10600 6452
rect 10652 6400 10658 6452
rect 10965 6443 11023 6449
rect 10965 6409 10977 6443
rect 11011 6409 11023 6443
rect 10965 6403 11023 6409
rect 9355 6344 9812 6372
rect 10505 6375 10563 6381
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 10505 6341 10517 6375
rect 10551 6372 10563 6375
rect 10980 6372 11008 6403
rect 11974 6400 11980 6452
rect 12032 6400 12038 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6409 12219 6443
rect 12161 6403 12219 6409
rect 12437 6443 12495 6449
rect 12437 6409 12449 6443
rect 12483 6409 12495 6443
rect 12437 6403 12495 6409
rect 10551 6344 11008 6372
rect 10551 6341 10563 6344
rect 10505 6335 10563 6341
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 3896 6100 3924 6267
rect 4540 6236 4568 6267
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 8754 6264 8760 6316
rect 8812 6264 8818 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 9953 6307 10011 6313
rect 9953 6304 9965 6307
rect 9732 6276 9965 6304
rect 9732 6264 9738 6276
rect 9953 6273 9965 6276
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6304 11851 6307
rect 12176 6304 12204 6403
rect 11839 6276 12204 6304
rect 11839 6273 11851 6276
rect 11793 6267 11851 6273
rect 12342 6264 12348 6316
rect 12400 6264 12406 6316
rect 12452 6236 12480 6403
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6409 13415 6443
rect 13357 6403 13415 6409
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 12989 6307 13047 6313
rect 12989 6273 13001 6307
rect 13035 6304 13047 6307
rect 13372 6304 13400 6403
rect 14274 6400 14280 6452
rect 14332 6400 14338 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6409 14979 6443
rect 14921 6403 14979 6409
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6372 14243 6375
rect 14936 6372 14964 6403
rect 15378 6400 15384 6452
rect 15436 6400 15442 6452
rect 15749 6443 15807 6449
rect 15749 6409 15761 6443
rect 15795 6409 15807 6443
rect 15749 6403 15807 6409
rect 14231 6344 14964 6372
rect 15289 6375 15347 6381
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 15289 6341 15301 6375
rect 15335 6372 15347 6375
rect 15764 6372 15792 6403
rect 16850 6400 16856 6452
rect 16908 6400 16914 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 15335 6344 15792 6372
rect 16761 6375 16819 6381
rect 15335 6341 15347 6344
rect 15289 6335 15347 6341
rect 16761 6341 16773 6375
rect 16807 6372 16819 6375
rect 17236 6372 17264 6403
rect 17954 6400 17960 6452
rect 18012 6400 18018 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6409 18199 6443
rect 18141 6403 18199 6409
rect 16807 6344 17264 6372
rect 17681 6375 17739 6381
rect 16807 6341 16819 6344
rect 16761 6335 16819 6341
rect 17681 6341 17693 6375
rect 17727 6372 17739 6375
rect 18156 6372 18184 6403
rect 19426 6400 19432 6452
rect 19484 6400 19490 6452
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6409 19855 6443
rect 19797 6403 19855 6409
rect 17727 6344 18184 6372
rect 19337 6375 19395 6381
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 19337 6341 19349 6375
rect 19383 6372 19395 6375
rect 19812 6372 19840 6403
rect 20346 6400 20352 6452
rect 20404 6400 20410 6452
rect 20809 6443 20867 6449
rect 20809 6409 20821 6443
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 20824 6372 20852 6403
rect 21542 6400 21548 6452
rect 21600 6400 21606 6452
rect 21821 6443 21879 6449
rect 21821 6409 21833 6443
rect 21867 6409 21879 6443
rect 21821 6403 21879 6409
rect 19383 6344 19840 6372
rect 20180 6344 20852 6372
rect 19383 6341 19395 6344
rect 19337 6335 19395 6341
rect 13035 6276 13400 6304
rect 13035 6273 13047 6276
rect 12989 6267 13047 6273
rect 13538 6264 13544 6316
rect 13596 6264 13602 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 15102 6264 15108 6316
rect 15160 6264 15166 6316
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15712 6276 15945 6304
rect 15712 6264 15718 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 18322 6264 18328 6316
rect 18380 6264 18386 6316
rect 19978 6264 19984 6316
rect 20036 6264 20042 6316
rect 20180 6313 20208 6344
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20993 6307 21051 6313
rect 20993 6273 21005 6307
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6304 21419 6307
rect 21836 6304 21864 6403
rect 22554 6400 22560 6452
rect 22612 6400 22618 6452
rect 22925 6443 22983 6449
rect 22925 6409 22937 6443
rect 22971 6409 22983 6443
rect 22925 6403 22983 6409
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 23523 6412 23888 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 22465 6375 22523 6381
rect 22465 6341 22477 6375
rect 22511 6372 22523 6375
rect 22940 6372 22968 6403
rect 23860 6381 23888 6412
rect 23934 6400 23940 6452
rect 23992 6400 23998 6452
rect 22511 6344 22968 6372
rect 23845 6375 23903 6381
rect 22511 6341 22523 6344
rect 22465 6335 22523 6341
rect 23845 6341 23857 6375
rect 23891 6341 23903 6375
rect 23845 6335 23903 6341
rect 21407 6276 21864 6304
rect 22005 6307 22063 6313
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 22005 6273 22017 6307
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 4540 6208 12480 6236
rect 5626 6128 5632 6180
rect 5684 6168 5690 6180
rect 20717 6171 20775 6177
rect 20717 6168 20729 6171
rect 5684 6140 20729 6168
rect 5684 6128 5690 6140
rect 20717 6137 20729 6140
rect 20763 6137 20775 6171
rect 21008 6168 21036 6267
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 22020 6236 22048 6267
rect 23106 6264 23112 6316
rect 23164 6264 23170 6316
rect 23658 6264 23664 6316
rect 23716 6264 23722 6316
rect 21692 6208 22048 6236
rect 21692 6196 21698 6208
rect 24210 6168 24216 6180
rect 21008 6140 24216 6168
rect 20717 6131 20775 6137
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 3896 6072 14841 6100
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 1104 6010 24840 6032
rect 1104 5958 3917 6010
rect 3969 5958 3981 6010
rect 4033 5958 4045 6010
rect 4097 5958 4109 6010
rect 4161 5958 4173 6010
rect 4225 5958 9851 6010
rect 9903 5958 9915 6010
rect 9967 5958 9979 6010
rect 10031 5958 10043 6010
rect 10095 5958 10107 6010
rect 10159 5958 15785 6010
rect 15837 5958 15849 6010
rect 15901 5958 15913 6010
rect 15965 5958 15977 6010
rect 16029 5958 16041 6010
rect 16093 5958 21719 6010
rect 21771 5958 21783 6010
rect 21835 5958 21847 6010
rect 21899 5958 21911 6010
rect 21963 5958 21975 6010
rect 22027 5958 24840 6010
rect 1104 5936 24840 5958
rect 6089 5899 6147 5905
rect 6089 5865 6101 5899
rect 6135 5896 6147 5899
rect 6546 5896 6552 5908
rect 6135 5868 6552 5896
rect 6135 5865 6147 5868
rect 6089 5859 6147 5865
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7558 5896 7564 5908
rect 7423 5868 7564 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 8573 5899 8631 5905
rect 8573 5865 8585 5899
rect 8619 5896 8631 5899
rect 8754 5896 8760 5908
rect 8619 5868 8760 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9674 5856 9680 5908
rect 9732 5856 9738 5908
rect 10873 5899 10931 5905
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11146 5896 11152 5908
rect 10919 5868 11152 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11146 5856 11152 5868
rect 11204 5856 11210 5908
rect 12253 5899 12311 5905
rect 12253 5865 12265 5899
rect 12299 5896 12311 5899
rect 12342 5896 12348 5908
rect 12299 5868 12348 5896
rect 12299 5865 12311 5868
rect 12253 5859 12311 5865
rect 12342 5856 12348 5868
rect 12400 5856 12406 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13538 5896 13544 5908
rect 13311 5868 13544 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14642 5896 14648 5908
rect 14415 5868 14648 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14642 5856 14648 5868
rect 14700 5856 14706 5908
rect 15102 5856 15108 5908
rect 15160 5856 15166 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15712 5868 15761 5896
rect 15712 5856 15718 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 16945 5899 17003 5905
rect 16945 5865 16957 5899
rect 16991 5896 17003 5899
rect 17402 5896 17408 5908
rect 16991 5868 17408 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 18233 5899 18291 5905
rect 18233 5865 18245 5899
rect 18279 5896 18291 5899
rect 18322 5896 18328 5908
rect 18279 5868 18328 5896
rect 18279 5865 18291 5868
rect 18233 5859 18291 5865
rect 18322 5856 18328 5868
rect 18380 5856 18386 5908
rect 19797 5899 19855 5905
rect 19797 5865 19809 5899
rect 19843 5896 19855 5899
rect 20530 5896 20536 5908
rect 19843 5868 20536 5896
rect 19843 5865 19855 5868
rect 19797 5859 19855 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 24486 5896 24492 5908
rect 24167 5868 24492 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 11793 5831 11851 5837
rect 11793 5797 11805 5831
rect 11839 5828 11851 5831
rect 12636 5828 12664 5856
rect 11839 5800 12664 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 9858 5652 9864 5704
rect 9916 5652 9922 5704
rect 11054 5652 11060 5704
rect 11112 5652 11118 5704
rect 11974 5652 11980 5704
rect 12032 5652 12038 5704
rect 12434 5652 12440 5704
rect 12492 5652 12498 5704
rect 13446 5652 13452 5704
rect 13504 5652 13510 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14826 5652 14832 5704
rect 14884 5652 14890 5704
rect 14645 5559 14703 5565
rect 14645 5525 14657 5559
rect 14691 5556 14703 5559
rect 15120 5556 15148 5856
rect 19978 5788 19984 5840
rect 20036 5828 20042 5840
rect 24026 5828 24032 5840
rect 20036 5800 24032 5828
rect 20036 5788 20042 5800
rect 24026 5788 24032 5800
rect 24084 5788 24090 5840
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 18414 5652 18420 5704
rect 18472 5652 18478 5704
rect 19978 5652 19984 5704
rect 20036 5652 20042 5704
rect 23842 5584 23848 5636
rect 23900 5584 23906 5636
rect 14691 5528 15148 5556
rect 14691 5525 14703 5528
rect 14645 5519 14703 5525
rect 1104 5466 25000 5488
rect 1104 5414 6884 5466
rect 6936 5414 6948 5466
rect 7000 5414 7012 5466
rect 7064 5414 7076 5466
rect 7128 5414 7140 5466
rect 7192 5414 12818 5466
rect 12870 5414 12882 5466
rect 12934 5414 12946 5466
rect 12998 5414 13010 5466
rect 13062 5414 13074 5466
rect 13126 5414 18752 5466
rect 18804 5414 18816 5466
rect 18868 5414 18880 5466
rect 18932 5414 18944 5466
rect 18996 5414 19008 5466
rect 19060 5414 24686 5466
rect 24738 5414 24750 5466
rect 24802 5414 24814 5466
rect 24866 5414 24878 5466
rect 24930 5414 24942 5466
rect 24994 5414 25000 5466
rect 1104 5392 25000 5414
rect 6270 5312 6276 5364
rect 6328 5352 6334 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 6328 5324 6377 5352
rect 6328 5312 6334 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 7558 5312 7564 5364
rect 7616 5312 7622 5364
rect 8754 5312 8760 5364
rect 8812 5312 8818 5364
rect 9858 5312 9864 5364
rect 9916 5312 9922 5364
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 11974 5312 11980 5364
rect 12032 5312 12038 5364
rect 12434 5312 12440 5364
rect 12492 5312 12498 5364
rect 13446 5312 13452 5364
rect 13504 5312 13510 5364
rect 14550 5312 14556 5364
rect 14608 5312 14614 5364
rect 14826 5312 14832 5364
rect 14884 5312 14890 5364
rect 15930 5312 15936 5364
rect 15988 5312 15994 5364
rect 17126 5312 17132 5364
rect 17184 5312 17190 5364
rect 18414 5312 18420 5364
rect 18472 5312 18478 5364
rect 19978 5312 19984 5364
rect 20036 5312 20042 5364
rect 23842 5312 23848 5364
rect 23900 5352 23906 5364
rect 24121 5355 24179 5361
rect 24121 5352 24133 5355
rect 23900 5324 24133 5352
rect 23900 5312 23906 5324
rect 24121 5321 24133 5324
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 13170 5284 13176 5296
rect 7760 5256 13176 5284
rect 7760 5225 7788 5256
rect 13170 5244 13176 5256
rect 13228 5244 13234 5296
rect 24394 5284 24400 5296
rect 16132 5256 24400 5284
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 7285 5219 7343 5225
rect 6595 5188 6960 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6932 5021 6960 5188
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7331 5188 7757 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5185 8999 5219
rect 8941 5179 8999 5185
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10962 5216 10968 5228
rect 10091 5188 10968 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 6917 5015 6975 5021
rect 6917 4981 6929 5015
rect 6963 5012 6975 5015
rect 8202 5012 8208 5024
rect 6963 4984 8208 5012
rect 6963 4981 6975 4984
rect 6917 4975 6975 4981
rect 8202 4972 8208 4984
rect 8260 4972 8266 5024
rect 8956 5012 8984 5179
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11238 5176 11244 5228
rect 11296 5176 11302 5228
rect 12161 5219 12219 5225
rect 12161 5185 12173 5219
rect 12207 5216 12219 5219
rect 12621 5219 12679 5225
rect 12207 5188 12434 5216
rect 12207 5185 12219 5188
rect 12161 5179 12219 5185
rect 12406 5080 12434 5188
rect 12621 5185 12633 5219
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12636 5148 12664 5179
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 16132 5225 16160 5256
rect 24394 5244 24400 5256
rect 24452 5244 24458 5296
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14516 5188 14749 5216
rect 14516 5176 14522 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 14182 5148 14188 5160
rect 12636 5120 14188 5148
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 15028 5148 15056 5179
rect 17126 5148 17132 5160
rect 15028 5120 17132 5148
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 17328 5148 17356 5179
rect 18598 5176 18604 5228
rect 18656 5176 18662 5228
rect 20165 5219 20223 5225
rect 20165 5185 20177 5219
rect 20211 5216 20223 5219
rect 21174 5216 21180 5228
rect 20211 5188 21180 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 23750 5148 23756 5160
rect 17328 5120 23756 5148
rect 23750 5108 23756 5120
rect 23808 5108 23814 5160
rect 22554 5080 22560 5092
rect 12406 5052 22560 5080
rect 22554 5040 22560 5052
rect 22612 5040 22618 5092
rect 17218 5012 17224 5024
rect 8956 4984 17224 5012
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 1104 4922 24840 4944
rect 1104 4870 3917 4922
rect 3969 4870 3981 4922
rect 4033 4870 4045 4922
rect 4097 4870 4109 4922
rect 4161 4870 4173 4922
rect 4225 4870 9851 4922
rect 9903 4870 9915 4922
rect 9967 4870 9979 4922
rect 10031 4870 10043 4922
rect 10095 4870 10107 4922
rect 10159 4870 15785 4922
rect 15837 4870 15849 4922
rect 15901 4870 15913 4922
rect 15965 4870 15977 4922
rect 16029 4870 16041 4922
rect 16093 4870 21719 4922
rect 21771 4870 21783 4922
rect 21835 4870 21847 4922
rect 21899 4870 21911 4922
rect 21963 4870 21975 4922
rect 22027 4870 24840 4922
rect 1104 4848 24840 4870
rect 24029 4811 24087 4817
rect 24029 4777 24041 4811
rect 24075 4808 24087 4811
rect 24302 4808 24308 4820
rect 24075 4780 24308 4808
rect 24075 4777 24087 4780
rect 24029 4771 24087 4777
rect 24302 4768 24308 4780
rect 24360 4768 24366 4820
rect 22922 4564 22928 4616
rect 22980 4604 22986 4616
rect 23937 4607 23995 4613
rect 23937 4604 23949 4607
rect 22980 4576 23949 4604
rect 22980 4564 22986 4576
rect 23937 4573 23949 4576
rect 23983 4573 23995 4607
rect 23937 4567 23995 4573
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 24228 4536 24256 4567
rect 23768 4508 24256 4536
rect 23768 4477 23796 4508
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4437 23811 4471
rect 23753 4431 23811 4437
rect 1104 4378 25000 4400
rect 1104 4326 6884 4378
rect 6936 4326 6948 4378
rect 7000 4326 7012 4378
rect 7064 4326 7076 4378
rect 7128 4326 7140 4378
rect 7192 4326 12818 4378
rect 12870 4326 12882 4378
rect 12934 4326 12946 4378
rect 12998 4326 13010 4378
rect 13062 4326 13074 4378
rect 13126 4326 18752 4378
rect 18804 4326 18816 4378
rect 18868 4326 18880 4378
rect 18932 4326 18944 4378
rect 18996 4326 19008 4378
rect 19060 4326 24686 4378
rect 24738 4326 24750 4378
rect 24802 4326 24814 4378
rect 24866 4326 24878 4378
rect 24930 4326 24942 4378
rect 24994 4326 25000 4378
rect 1104 4304 25000 4326
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 7708 4236 18000 4264
rect 7708 4224 7714 4236
rect 17972 4208 18000 4236
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 17862 4196 17868 4208
rect 17184 4168 17868 4196
rect 17184 4156 17190 4168
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 17954 4156 17960 4208
rect 18012 4156 18018 4208
rect 1104 3834 24840 3856
rect 1104 3782 3917 3834
rect 3969 3782 3981 3834
rect 4033 3782 4045 3834
rect 4097 3782 4109 3834
rect 4161 3782 4173 3834
rect 4225 3782 9851 3834
rect 9903 3782 9915 3834
rect 9967 3782 9979 3834
rect 10031 3782 10043 3834
rect 10095 3782 10107 3834
rect 10159 3782 15785 3834
rect 15837 3782 15849 3834
rect 15901 3782 15913 3834
rect 15965 3782 15977 3834
rect 16029 3782 16041 3834
rect 16093 3782 21719 3834
rect 21771 3782 21783 3834
rect 21835 3782 21847 3834
rect 21899 3782 21911 3834
rect 21963 3782 21975 3834
rect 22027 3782 24840 3834
rect 1104 3760 24840 3782
rect 23658 3680 23664 3732
rect 23716 3720 23722 3732
rect 23937 3723 23995 3729
rect 23937 3720 23949 3723
rect 23716 3692 23949 3720
rect 23716 3680 23722 3692
rect 23937 3689 23949 3692
rect 23983 3689 23995 3723
rect 23937 3683 23995 3689
rect 24118 3476 24124 3528
rect 24176 3476 24182 3528
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 22186 3448 22192 3460
rect 13688 3420 22192 3448
rect 13688 3408 13694 3420
rect 22186 3408 22192 3420
rect 22244 3408 22250 3460
rect 1104 3290 25000 3312
rect 1104 3238 6884 3290
rect 6936 3238 6948 3290
rect 7000 3238 7012 3290
rect 7064 3238 7076 3290
rect 7128 3238 7140 3290
rect 7192 3238 12818 3290
rect 12870 3238 12882 3290
rect 12934 3238 12946 3290
rect 12998 3238 13010 3290
rect 13062 3238 13074 3290
rect 13126 3238 18752 3290
rect 18804 3238 18816 3290
rect 18868 3238 18880 3290
rect 18932 3238 18944 3290
rect 18996 3238 19008 3290
rect 19060 3238 24686 3290
rect 24738 3238 24750 3290
rect 24802 3238 24814 3290
rect 24866 3238 24878 3290
rect 24930 3238 24942 3290
rect 24994 3238 25000 3290
rect 1104 3216 25000 3238
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 16666 3108 16672 3120
rect 11020 3080 16672 3108
rect 11020 3068 11026 3080
rect 16666 3068 16672 3080
rect 16724 3068 16730 3120
rect 25038 3108 25044 3120
rect 23492 3080 25044 3108
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 10410 3040 10416 3052
rect 1452 3012 10416 3040
rect 1452 3000 1458 3012
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 15194 3040 15200 3052
rect 11296 3012 15200 3040
rect 11296 3000 11302 3012
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 23492 3049 23520 3080
rect 25038 3068 25044 3080
rect 25096 3068 25102 3120
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23753 3043 23811 3049
rect 23753 3009 23765 3043
rect 23799 3009 23811 3043
rect 23753 3003 23811 3009
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 5902 2932 5908 2984
rect 5960 2972 5966 2984
rect 9582 2972 9588 2984
rect 5960 2944 9588 2972
rect 5960 2932 5966 2944
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 10778 2932 10784 2984
rect 10836 2972 10842 2984
rect 10836 2944 16804 2972
rect 10836 2932 10842 2944
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 7466 2904 7472 2916
rect 2740 2876 7472 2904
rect 2740 2864 2746 2876
rect 7466 2864 7472 2876
rect 7524 2864 7530 2916
rect 8018 2864 8024 2916
rect 8076 2904 8082 2916
rect 15010 2904 15016 2916
rect 8076 2876 15016 2904
rect 8076 2864 8082 2876
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 16776 2848 16804 2944
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 22278 2972 22284 2984
rect 17276 2944 22284 2972
rect 17276 2932 17282 2944
rect 22278 2932 22284 2944
rect 22336 2932 22342 2984
rect 23768 2904 23796 3003
rect 24044 2972 24072 3003
rect 24302 3000 24308 3052
rect 24360 3000 24366 3052
rect 24486 2972 24492 2984
rect 24044 2944 24492 2972
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 24578 2904 24584 2916
rect 23768 2876 24584 2904
rect 24578 2864 24584 2876
rect 24636 2864 24642 2916
rect 1946 2796 1952 2848
rect 2004 2836 2010 2848
rect 6730 2836 6736 2848
rect 2004 2808 6736 2836
rect 2004 2796 2010 2808
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 9490 2796 9496 2848
rect 9548 2836 9554 2848
rect 12434 2836 12440 2848
rect 9548 2808 12440 2836
rect 9548 2796 9554 2808
rect 12434 2796 12440 2808
rect 12492 2796 12498 2848
rect 16758 2796 16764 2848
rect 16816 2796 16822 2848
rect 22830 2796 22836 2848
rect 22888 2836 22894 2848
rect 23293 2839 23351 2845
rect 23293 2836 23305 2839
rect 22888 2808 23305 2836
rect 22888 2796 22894 2808
rect 23293 2805 23305 2808
rect 23339 2805 23351 2839
rect 23293 2799 23351 2805
rect 23569 2839 23627 2845
rect 23569 2805 23581 2839
rect 23615 2836 23627 2839
rect 23658 2836 23664 2848
rect 23615 2808 23664 2836
rect 23615 2805 23627 2808
rect 23569 2799 23627 2805
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24026 2836 24032 2848
rect 23891 2808 24032 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 1104 2746 24840 2768
rect 1104 2694 3917 2746
rect 3969 2694 3981 2746
rect 4033 2694 4045 2746
rect 4097 2694 4109 2746
rect 4161 2694 4173 2746
rect 4225 2694 9851 2746
rect 9903 2694 9915 2746
rect 9967 2694 9979 2746
rect 10031 2694 10043 2746
rect 10095 2694 10107 2746
rect 10159 2694 15785 2746
rect 15837 2694 15849 2746
rect 15901 2694 15913 2746
rect 15965 2694 15977 2746
rect 16029 2694 16041 2746
rect 16093 2694 21719 2746
rect 21771 2694 21783 2746
rect 21835 2694 21847 2746
rect 21899 2694 21911 2746
rect 21963 2694 21975 2746
rect 22027 2694 24840 2746
rect 1104 2672 24840 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 3418 2632 3424 2644
rect 1719 2604 3424 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 3418 2592 3424 2604
rect 3476 2592 3482 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 10686 2632 10692 2644
rect 7248 2604 10692 2632
rect 7248 2592 7254 2604
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 16301 2635 16359 2641
rect 11112 2604 16068 2632
rect 11112 2592 11118 2604
rect 1578 2524 1584 2576
rect 1636 2524 1642 2576
rect 1946 2524 1952 2576
rect 2004 2524 2010 2576
rect 7834 2524 7840 2576
rect 7892 2564 7898 2576
rect 10778 2564 10784 2576
rect 7892 2536 10784 2564
rect 7892 2524 7898 2536
rect 10778 2524 10784 2536
rect 10836 2524 10842 2576
rect 11974 2524 11980 2576
rect 12032 2564 12038 2576
rect 15105 2567 15163 2573
rect 12032 2536 13308 2564
rect 12032 2524 12038 2536
rect 474 2456 480 2508
rect 532 2496 538 2508
rect 532 2468 2176 2496
rect 532 2456 538 2468
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 2148 2437 2176 2468
rect 2590 2456 2596 2508
rect 2648 2496 2654 2508
rect 10870 2496 10876 2508
rect 2648 2468 7328 2496
rect 2648 2456 2654 2468
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 1360 2400 1409 2428
rect 1360 2388 1366 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2397 2191 2431
rect 2133 2391 2191 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1872 2360 1900 2391
rect 256 2332 1900 2360
rect 256 2320 262 2332
rect 1946 2320 1952 2372
rect 2004 2360 2010 2372
rect 2240 2360 2268 2391
rect 4614 2388 4620 2440
rect 4672 2428 4678 2440
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 4672 2400 4905 2428
rect 4672 2388 4678 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 6086 2388 6092 2440
rect 6144 2388 6150 2440
rect 7190 2388 7196 2440
rect 7248 2388 7254 2440
rect 7208 2360 7236 2388
rect 2004 2332 2268 2360
rect 2424 2332 7236 2360
rect 7300 2360 7328 2468
rect 9232 2468 10876 2496
rect 7374 2388 7380 2440
rect 7432 2388 7438 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 9232 2428 9260 2468
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 11020 2468 12848 2496
rect 11020 2456 11026 2468
rect 7800 2400 9260 2428
rect 7800 2388 7806 2400
rect 9306 2388 9312 2440
rect 9364 2428 9370 2440
rect 9585 2431 9643 2437
rect 9585 2428 9597 2431
rect 9364 2400 9597 2428
rect 9364 2388 9370 2400
rect 9585 2397 9597 2400
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9732 2400 9873 2428
rect 9732 2388 9738 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 7300 2332 9168 2360
rect 2004 2320 2010 2332
rect 2424 2301 2452 2332
rect 9140 2304 9168 2332
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 10428 2360 10456 2391
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 10652 2400 11161 2428
rect 10652 2388 10658 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11701 2431 11759 2437
rect 11701 2397 11713 2431
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11716 2360 11744 2391
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11848 2400 11989 2428
rect 11848 2388 11854 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12253 2431 12311 2437
rect 12253 2397 12265 2431
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 12268 2360 12296 2391
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12820 2437 12848 2468
rect 13280 2437 13308 2536
rect 15105 2533 15117 2567
rect 15151 2564 15163 2567
rect 15151 2536 15700 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 13446 2456 13452 2508
rect 13504 2496 13510 2508
rect 13504 2468 15608 2496
rect 13504 2456 13510 2468
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 15286 2388 15292 2440
rect 15344 2388 15350 2440
rect 15580 2437 15608 2468
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2397 15623 2431
rect 15672 2428 15700 2536
rect 16040 2508 16068 2604
rect 16301 2601 16313 2635
rect 16347 2632 16359 2635
rect 17402 2632 17408 2644
rect 16347 2604 17408 2632
rect 16347 2601 16359 2604
rect 16301 2595 16359 2601
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 17862 2592 17868 2644
rect 17920 2632 17926 2644
rect 22557 2635 22615 2641
rect 22557 2632 22569 2635
rect 17920 2604 22569 2632
rect 17920 2592 17926 2604
rect 22557 2601 22569 2604
rect 22603 2601 22615 2635
rect 22557 2595 22615 2601
rect 22922 2592 22928 2644
rect 22980 2592 22986 2644
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2632 23259 2635
rect 23247 2604 23612 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 16577 2567 16635 2573
rect 16577 2533 16589 2567
rect 16623 2533 16635 2567
rect 16577 2527 16635 2533
rect 16022 2456 16028 2508
rect 16080 2456 16086 2508
rect 16592 2496 16620 2527
rect 18598 2524 18604 2576
rect 18656 2564 18662 2576
rect 23477 2567 23535 2573
rect 23477 2564 23489 2567
rect 18656 2536 20668 2564
rect 18656 2524 18662 2536
rect 16592 2468 17356 2496
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15672 2400 15945 2428
rect 15565 2391 15623 2397
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16482 2388 16488 2440
rect 16540 2388 16546 2440
rect 16758 2388 16764 2440
rect 16816 2388 16822 2440
rect 17328 2437 17356 2468
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 20640 2496 20668 2536
rect 23308 2536 23489 2564
rect 23308 2496 23336 2536
rect 23477 2533 23489 2536
rect 23523 2533 23535 2567
rect 23584 2564 23612 2604
rect 23750 2592 23756 2644
rect 23808 2592 23814 2644
rect 24302 2592 24308 2644
rect 24360 2592 24366 2644
rect 24320 2564 24348 2592
rect 23584 2536 24348 2564
rect 23477 2527 23535 2533
rect 18012 2468 19012 2496
rect 18012 2456 18018 2468
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 15289 2387 15347 2388
rect 17052 2360 17080 2391
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 17862 2388 17868 2440
rect 17920 2388 17926 2440
rect 18138 2388 18144 2440
rect 18196 2388 18202 2440
rect 18414 2388 18420 2440
rect 18472 2388 18478 2440
rect 18690 2388 18696 2440
rect 18748 2388 18754 2440
rect 18984 2437 19012 2468
rect 19352 2468 20576 2496
rect 20640 2468 23336 2496
rect 18969 2431 19027 2437
rect 18969 2397 18981 2431
rect 19015 2397 19027 2431
rect 18969 2391 19027 2397
rect 18322 2360 18328 2372
rect 9272 2332 10456 2360
rect 10980 2332 11744 2360
rect 11808 2332 12296 2360
rect 16776 2332 17080 2360
rect 17420 2332 18328 2360
rect 9272 2320 9278 2332
rect 2409 2295 2467 2301
rect 2409 2261 2421 2295
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 4246 2292 4252 2304
rect 2924 2264 4252 2292
rect 2924 2252 2930 2264
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4338 2252 4344 2304
rect 4396 2292 4402 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4396 2264 4721 2292
rect 4396 2252 4402 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 6270 2252 6276 2304
rect 6328 2252 6334 2304
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2292 7251 2295
rect 8110 2292 8116 2304
rect 7239 2264 8116 2292
rect 7239 2261 7251 2264
rect 7193 2255 7251 2261
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 9122 2252 9128 2304
rect 9180 2252 9186 2304
rect 9398 2252 9404 2304
rect 9456 2252 9462 2304
rect 9677 2295 9735 2301
rect 9677 2261 9689 2295
rect 9723 2292 9735 2295
rect 9766 2292 9772 2304
rect 9723 2264 9772 2292
rect 9723 2261 9735 2264
rect 9677 2255 9735 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10229 2295 10287 2301
rect 10229 2261 10241 2295
rect 10275 2292 10287 2295
rect 10870 2292 10876 2304
rect 10275 2264 10876 2292
rect 10275 2261 10287 2264
rect 10229 2255 10287 2261
rect 10870 2252 10876 2264
rect 10928 2252 10934 2304
rect 10980 2301 11008 2332
rect 10965 2295 11023 2301
rect 10965 2261 10977 2295
rect 11011 2261 11023 2295
rect 10965 2255 11023 2261
rect 11514 2252 11520 2304
rect 11572 2252 11578 2304
rect 11808 2301 11836 2332
rect 11793 2295 11851 2301
rect 11793 2261 11805 2295
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12066 2252 12072 2304
rect 12124 2252 12130 2304
rect 12342 2252 12348 2304
rect 12400 2252 12406 2304
rect 12618 2252 12624 2304
rect 12676 2252 12682 2304
rect 13081 2295 13139 2301
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 13998 2292 14004 2304
rect 13127 2264 14004 2292
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 13998 2252 14004 2264
rect 14056 2252 14062 2304
rect 14090 2252 14096 2304
rect 14148 2292 14154 2304
rect 15102 2292 15108 2304
rect 14148 2264 15108 2292
rect 14148 2252 14154 2264
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 15378 2252 15384 2304
rect 15436 2252 15442 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15620 2264 16129 2292
rect 15620 2252 15626 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16298 2252 16304 2304
rect 16356 2292 16362 2304
rect 16776 2292 16804 2332
rect 16356 2264 16804 2292
rect 16356 2252 16362 2264
rect 16850 2252 16856 2304
rect 16908 2252 16914 2304
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17420 2301 17448 2332
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 17000 2264 17141 2292
rect 17000 2252 17006 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17405 2295 17463 2301
rect 17405 2261 17417 2295
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17681 2295 17739 2301
rect 17681 2261 17693 2295
rect 17727 2292 17739 2295
rect 17770 2292 17776 2304
rect 17727 2264 17776 2292
rect 17727 2261 17739 2264
rect 17681 2255 17739 2261
rect 17770 2252 17776 2264
rect 17828 2252 17834 2304
rect 17957 2295 18015 2301
rect 17957 2261 17969 2295
rect 18003 2292 18015 2295
rect 18138 2292 18144 2304
rect 18003 2264 18144 2292
rect 18003 2261 18015 2264
rect 17957 2255 18015 2261
rect 18138 2252 18144 2264
rect 18196 2252 18202 2304
rect 18230 2252 18236 2304
rect 18288 2252 18294 2304
rect 18509 2295 18567 2301
rect 18509 2261 18521 2295
rect 18555 2292 18567 2295
rect 18598 2292 18604 2304
rect 18555 2264 18604 2292
rect 18555 2261 18567 2264
rect 18509 2255 18567 2261
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 18785 2295 18843 2301
rect 18785 2261 18797 2295
rect 18831 2292 18843 2295
rect 19150 2292 19156 2304
rect 18831 2264 19156 2292
rect 18831 2261 18843 2264
rect 18785 2255 18843 2261
rect 19150 2252 19156 2264
rect 19208 2252 19214 2304
rect 19242 2252 19248 2304
rect 19300 2252 19306 2304
rect 19352 2292 19380 2468
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2397 19487 2431
rect 19429 2391 19487 2397
rect 19444 2360 19472 2391
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2428 20039 2431
rect 20162 2428 20168 2440
rect 20027 2400 20168 2428
rect 20027 2397 20039 2400
rect 19981 2391 20039 2397
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 20254 2388 20260 2440
rect 20312 2388 20318 2440
rect 20548 2437 20576 2468
rect 20533 2431 20591 2437
rect 20533 2397 20545 2431
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2397 20867 2431
rect 20809 2391 20867 2397
rect 19444 2332 20116 2360
rect 19521 2295 19579 2301
rect 19521 2292 19533 2295
rect 19352 2264 19533 2292
rect 19521 2261 19533 2264
rect 19567 2261 19579 2295
rect 19521 2255 19579 2261
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2292 19855 2295
rect 19978 2292 19984 2304
rect 19843 2264 19984 2292
rect 19843 2261 19855 2264
rect 19797 2255 19855 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20088 2301 20116 2332
rect 20438 2320 20444 2372
rect 20496 2360 20502 2372
rect 20824 2360 20852 2391
rect 22370 2388 22376 2440
rect 22428 2388 22434 2440
rect 22830 2388 22836 2440
rect 22888 2388 22894 2440
rect 23109 2431 23167 2437
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23290 2428 23296 2440
rect 23155 2400 23296 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23382 2388 23388 2440
rect 23440 2388 23446 2440
rect 23661 2431 23719 2437
rect 23661 2397 23673 2431
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 20496 2332 20852 2360
rect 23676 2360 23704 2391
rect 23934 2388 23940 2440
rect 23992 2388 23998 2440
rect 24026 2388 24032 2440
rect 24084 2428 24090 2440
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 24084 2400 24225 2428
rect 24084 2388 24090 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 23676 2332 24256 2360
rect 20496 2320 20502 2332
rect 24228 2304 24256 2332
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20346 2252 20352 2304
rect 20404 2252 20410 2304
rect 20622 2252 20628 2304
rect 20680 2252 20686 2304
rect 22649 2295 22707 2301
rect 22649 2261 22661 2295
rect 22695 2292 22707 2295
rect 22738 2292 22744 2304
rect 22695 2264 22744 2292
rect 22695 2261 22707 2264
rect 22649 2255 22707 2261
rect 22738 2252 22744 2264
rect 22796 2252 22802 2304
rect 24026 2252 24032 2304
rect 24084 2252 24090 2304
rect 24210 2252 24216 2304
rect 24268 2252 24274 2304
rect 1104 2202 25000 2224
rect 1104 2150 6884 2202
rect 6936 2150 6948 2202
rect 7000 2150 7012 2202
rect 7064 2150 7076 2202
rect 7128 2150 7140 2202
rect 7192 2150 12818 2202
rect 12870 2150 12882 2202
rect 12934 2150 12946 2202
rect 12998 2150 13010 2202
rect 13062 2150 13074 2202
rect 13126 2150 18752 2202
rect 18804 2150 18816 2202
rect 18868 2150 18880 2202
rect 18932 2150 18944 2202
rect 18996 2150 19008 2202
rect 19060 2150 24686 2202
rect 24738 2150 24750 2202
rect 24802 2150 24814 2202
rect 24866 2150 24878 2202
rect 24930 2150 24942 2202
rect 24994 2150 25000 2202
rect 1104 2128 25000 2150
rect 2409 2091 2467 2097
rect 2409 2088 2421 2091
rect 1688 2060 2421 2088
rect 1688 1961 1716 2060
rect 2409 2057 2421 2060
rect 2455 2057 2467 2091
rect 2409 2051 2467 2057
rect 2682 2048 2688 2100
rect 2740 2048 2746 2100
rect 3896 2060 6868 2088
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 1762 1912 1768 1964
rect 1820 1912 1826 1964
rect 2130 1912 2136 1964
rect 2188 1912 2194 1964
rect 2593 1955 2651 1961
rect 2593 1921 2605 1955
rect 2639 1921 2651 1955
rect 2869 1955 2927 1961
rect 2869 1952 2881 1955
rect 2593 1915 2651 1921
rect 2746 1924 2881 1952
rect 750 1844 756 1896
rect 808 1884 814 1896
rect 2608 1884 2636 1915
rect 808 1856 2636 1884
rect 808 1844 814 1856
rect 1026 1776 1032 1828
rect 1084 1816 1090 1828
rect 2746 1816 2774 1924
rect 2869 1921 2881 1924
rect 2915 1921 2927 1955
rect 2869 1915 2927 1921
rect 3142 1912 3148 1964
rect 3200 1912 3206 1964
rect 3421 1956 3479 1961
rect 3421 1955 3556 1956
rect 3421 1921 3433 1955
rect 3467 1952 3556 1955
rect 3602 1952 3608 1964
rect 3467 1928 3608 1952
rect 3467 1921 3479 1928
rect 3528 1924 3608 1928
rect 3421 1915 3479 1921
rect 3602 1912 3608 1924
rect 3660 1912 3666 1964
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1952 3755 1955
rect 3786 1952 3792 1964
rect 3743 1924 3792 1952
rect 3743 1921 3755 1924
rect 3697 1915 3755 1921
rect 3786 1912 3792 1924
rect 3844 1912 3850 1964
rect 1084 1788 2774 1816
rect 1084 1776 1090 1788
rect 3326 1776 3332 1828
rect 3384 1816 3390 1828
rect 3513 1819 3571 1825
rect 3513 1816 3525 1819
rect 3384 1788 3525 1816
rect 3384 1776 3390 1788
rect 3513 1785 3525 1788
rect 3559 1785 3571 1819
rect 3513 1779 3571 1785
rect 3602 1776 3608 1828
rect 3660 1816 3666 1828
rect 3789 1819 3847 1825
rect 3789 1816 3801 1819
rect 3660 1788 3801 1816
rect 3660 1776 3666 1788
rect 3789 1785 3801 1788
rect 3835 1785 3847 1819
rect 3789 1779 3847 1785
rect 1486 1708 1492 1760
rect 1544 1708 1550 1760
rect 1949 1751 2007 1757
rect 1949 1717 1961 1751
rect 1995 1748 2007 1751
rect 2222 1748 2228 1760
rect 1995 1720 2228 1748
rect 1995 1717 2007 1720
rect 1949 1711 2007 1717
rect 2222 1708 2228 1720
rect 2280 1708 2286 1760
rect 2314 1708 2320 1760
rect 2372 1708 2378 1760
rect 2958 1708 2964 1760
rect 3016 1708 3022 1760
rect 3237 1751 3295 1757
rect 3237 1717 3249 1751
rect 3283 1748 3295 1751
rect 3896 1748 3924 2060
rect 3973 1955 4031 1961
rect 3973 1921 3985 1955
rect 4019 1921 4031 1955
rect 3973 1915 4031 1921
rect 3988 1884 4016 1915
rect 4246 1912 4252 1964
rect 4304 1912 4310 1964
rect 4525 1955 4583 1961
rect 4525 1921 4537 1955
rect 4571 1952 4583 1955
rect 4706 1952 4712 1964
rect 4571 1924 4712 1952
rect 4571 1921 4583 1924
rect 4525 1915 4583 1921
rect 4706 1912 4712 1924
rect 4764 1912 4770 1964
rect 4801 1955 4859 1961
rect 4801 1921 4813 1955
rect 4847 1952 4859 1955
rect 4982 1952 4988 1964
rect 4847 1924 4988 1952
rect 4847 1921 4859 1924
rect 4801 1915 4859 1921
rect 4982 1912 4988 1924
rect 5040 1912 5046 1964
rect 5077 1955 5135 1961
rect 5077 1921 5089 1955
rect 5123 1952 5135 1955
rect 5258 1952 5264 1964
rect 5123 1924 5264 1952
rect 5123 1921 5135 1924
rect 5077 1915 5135 1921
rect 5258 1912 5264 1924
rect 5316 1912 5322 1964
rect 5353 1955 5411 1961
rect 5353 1921 5365 1955
rect 5399 1921 5411 1955
rect 5353 1915 5411 1921
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 5629 1915 5687 1921
rect 5721 1955 5779 1961
rect 5721 1921 5733 1955
rect 5767 1921 5779 1955
rect 5721 1915 5779 1921
rect 6181 1955 6239 1961
rect 6181 1921 6193 1955
rect 6227 1952 6239 1955
rect 6546 1952 6552 1964
rect 6227 1924 6552 1952
rect 6227 1921 6239 1924
rect 6181 1915 6239 1921
rect 4430 1884 4436 1896
rect 3988 1856 4436 1884
rect 4430 1844 4436 1856
rect 4488 1844 4494 1896
rect 5368 1884 5396 1915
rect 4632 1856 5396 1884
rect 4632 1825 4660 1856
rect 4617 1819 4675 1825
rect 4617 1785 4629 1819
rect 4663 1785 4675 1819
rect 4617 1779 4675 1785
rect 4893 1819 4951 1825
rect 4893 1785 4905 1819
rect 4939 1816 4951 1819
rect 5644 1816 5672 1915
rect 5736 1884 5764 1915
rect 6546 1912 6552 1924
rect 6604 1912 6610 1964
rect 6638 1912 6644 1964
rect 6696 1912 6702 1964
rect 6840 1952 6868 2060
rect 7466 2048 7472 2100
rect 7524 2048 7530 2100
rect 7561 2091 7619 2097
rect 7561 2057 7573 2091
rect 7607 2088 7619 2091
rect 7742 2088 7748 2100
rect 7607 2060 7748 2088
rect 7607 2057 7619 2060
rect 7561 2051 7619 2057
rect 7742 2048 7748 2060
rect 7800 2048 7806 2100
rect 7834 2048 7840 2100
rect 7892 2048 7898 2100
rect 8018 2048 8024 2100
rect 8076 2088 8082 2100
rect 8113 2091 8171 2097
rect 8113 2088 8125 2091
rect 8076 2060 8125 2088
rect 8076 2048 8082 2060
rect 8113 2057 8125 2060
rect 8159 2057 8171 2091
rect 8113 2051 8171 2057
rect 8680 2060 11008 2088
rect 7484 2020 7512 2048
rect 7484 1992 8616 2020
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 6840 1924 6929 1952
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7009 1955 7067 1961
rect 7009 1921 7021 1955
rect 7055 1952 7067 1955
rect 7374 1952 7380 1964
rect 7055 1924 7380 1952
rect 7055 1921 7067 1924
rect 7009 1915 7067 1921
rect 7374 1912 7380 1924
rect 7432 1912 7438 1964
rect 7466 1912 7472 1964
rect 7524 1912 7530 1964
rect 7742 1912 7748 1964
rect 7800 1912 7806 1964
rect 8018 1912 8024 1964
rect 8076 1912 8082 1964
rect 8294 1912 8300 1964
rect 8352 1912 8358 1964
rect 8588 1961 8616 1992
rect 8573 1955 8631 1961
rect 8573 1921 8585 1955
rect 8619 1921 8631 1955
rect 8573 1915 8631 1921
rect 6270 1884 6276 1896
rect 5736 1856 6276 1884
rect 6270 1844 6276 1856
rect 6328 1844 6334 1896
rect 7558 1884 7564 1896
rect 6840 1856 7564 1884
rect 4939 1788 5672 1816
rect 5905 1819 5963 1825
rect 4939 1785 4951 1788
rect 4893 1779 4951 1785
rect 5905 1785 5917 1819
rect 5951 1816 5963 1819
rect 6840 1816 6868 1856
rect 7558 1844 7564 1856
rect 7616 1844 7622 1896
rect 7834 1844 7840 1896
rect 7892 1884 7898 1896
rect 8680 1884 8708 2060
rect 8754 1980 8760 2032
rect 8812 2020 8818 2032
rect 8812 1992 9996 2020
rect 8812 1980 8818 1992
rect 8846 1912 8852 1964
rect 8904 1912 8910 1964
rect 9122 1912 9128 1964
rect 9180 1912 9186 1964
rect 9398 1961 9404 1964
rect 9393 1952 9404 1961
rect 9359 1924 9404 1952
rect 9393 1915 9404 1924
rect 9398 1912 9404 1915
rect 9456 1912 9462 1964
rect 9968 1961 9996 1992
rect 10410 1980 10416 2032
rect 10468 1980 10474 2032
rect 10980 2029 11008 2060
rect 12618 2048 12624 2100
rect 12676 2088 12682 2100
rect 13541 2091 13599 2097
rect 12676 2060 13492 2088
rect 12676 2048 12682 2060
rect 10965 2023 11023 2029
rect 10965 1989 10977 2023
rect 11011 1989 11023 2023
rect 10965 1983 11023 1989
rect 11238 1980 11244 2032
rect 11296 2020 11302 2032
rect 11977 2023 12035 2029
rect 11977 2020 11989 2023
rect 11296 1992 11989 2020
rect 11296 1980 11302 1992
rect 11977 1989 11989 1992
rect 12023 1989 12035 2023
rect 12805 2023 12863 2029
rect 12805 2020 12817 2023
rect 11977 1983 12035 1989
rect 12084 1992 12817 2020
rect 9677 1955 9735 1961
rect 9677 1952 9689 1955
rect 9600 1936 9689 1952
rect 9508 1924 9689 1936
rect 9508 1908 9628 1924
rect 9677 1921 9689 1924
rect 9723 1921 9735 1955
rect 9677 1915 9735 1921
rect 9953 1955 10011 1961
rect 9953 1921 9965 1955
rect 9999 1921 10011 1955
rect 9953 1915 10011 1921
rect 10042 1912 10048 1964
rect 10100 1912 10106 1964
rect 10229 1955 10287 1961
rect 10229 1921 10241 1955
rect 10275 1952 10287 1955
rect 10318 1952 10324 1964
rect 10275 1924 10324 1952
rect 10275 1921 10287 1924
rect 10229 1915 10287 1921
rect 10318 1912 10324 1924
rect 10376 1912 10382 1964
rect 11330 1912 11336 1964
rect 11388 1952 11394 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 11388 1924 11529 1952
rect 11388 1912 11394 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 12084 1952 12112 1992
rect 12805 1989 12817 1992
rect 12851 1989 12863 2023
rect 12805 1983 12863 1989
rect 11517 1915 11575 1921
rect 11624 1924 12112 1952
rect 9508 1884 9536 1908
rect 7892 1856 8708 1884
rect 8956 1856 9536 1884
rect 10060 1884 10088 1912
rect 11624 1884 11652 1924
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 13464 1961 13492 2060
rect 13541 2057 13553 2091
rect 13587 2088 13599 2091
rect 13587 2060 13952 2088
rect 13587 2057 13599 2060
rect 13541 2051 13599 2057
rect 12621 1956 12679 1961
rect 12452 1955 12679 1956
rect 12452 1952 12633 1955
rect 12400 1928 12633 1952
rect 12400 1924 12480 1928
rect 12400 1912 12406 1924
rect 12621 1921 12633 1928
rect 12667 1921 12679 1955
rect 12621 1915 12679 1921
rect 13449 1955 13507 1961
rect 13449 1921 13461 1955
rect 13495 1921 13507 1955
rect 13449 1915 13507 1921
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 13725 1955 13783 1961
rect 13725 1952 13737 1955
rect 13596 1924 13737 1952
rect 13596 1912 13602 1924
rect 13725 1921 13737 1924
rect 13771 1921 13783 1955
rect 13924 1952 13952 2060
rect 13998 2048 14004 2100
rect 14056 2048 14062 2100
rect 14185 2091 14243 2097
rect 14185 2057 14197 2091
rect 14231 2088 14243 2091
rect 15286 2088 15292 2100
rect 14231 2060 15292 2088
rect 14231 2057 14243 2060
rect 14185 2051 14243 2057
rect 15286 2048 15292 2060
rect 15344 2048 15350 2100
rect 15378 2048 15384 2100
rect 15436 2088 15442 2100
rect 17405 2091 17463 2097
rect 15436 2060 15884 2088
rect 15436 2048 15442 2060
rect 14016 2020 14044 2048
rect 15856 2029 15884 2060
rect 17405 2057 17417 2091
rect 17451 2088 17463 2091
rect 17586 2088 17592 2100
rect 17451 2060 17592 2088
rect 17451 2057 17463 2060
rect 17405 2051 17463 2057
rect 17586 2048 17592 2060
rect 17644 2048 17650 2100
rect 17681 2091 17739 2097
rect 17681 2057 17693 2091
rect 17727 2088 17739 2091
rect 17862 2088 17868 2100
rect 17727 2060 17868 2088
rect 17727 2057 17739 2060
rect 17681 2051 17739 2057
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 18230 2048 18236 2100
rect 18288 2048 18294 2100
rect 18322 2048 18328 2100
rect 18380 2088 18386 2100
rect 18380 2060 18736 2088
rect 18380 2048 18386 2060
rect 15841 2023 15899 2029
rect 14016 1992 14872 2020
rect 13998 1952 14004 1964
rect 13924 1924 14004 1952
rect 13725 1915 13783 1921
rect 13998 1912 14004 1924
rect 14056 1912 14062 1964
rect 14093 1955 14151 1961
rect 14093 1921 14105 1955
rect 14139 1952 14151 1955
rect 14274 1952 14280 1964
rect 14139 1924 14280 1952
rect 14139 1921 14151 1924
rect 14093 1915 14151 1921
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14366 1912 14372 1964
rect 14424 1912 14430 1964
rect 14844 1961 14872 1992
rect 15028 1992 15700 2020
rect 14461 1955 14519 1961
rect 14461 1921 14473 1955
rect 14507 1921 14519 1955
rect 14461 1915 14519 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1921 14887 1955
rect 14829 1915 14887 1921
rect 10060 1856 11652 1884
rect 7892 1844 7898 1856
rect 5951 1788 6868 1816
rect 7193 1819 7251 1825
rect 5951 1785 5963 1788
rect 5905 1779 5963 1785
rect 7193 1785 7205 1819
rect 7239 1816 7251 1819
rect 8110 1816 8116 1828
rect 7239 1788 8116 1816
rect 7239 1785 7251 1788
rect 7193 1779 7251 1785
rect 8110 1776 8116 1788
rect 8168 1776 8174 1828
rect 8956 1825 8984 1856
rect 12066 1844 12072 1896
rect 12124 1884 12130 1896
rect 14476 1884 14504 1915
rect 12124 1856 14504 1884
rect 12124 1844 12130 1856
rect 8941 1819 8999 1825
rect 8941 1785 8953 1819
rect 8987 1785 8999 1819
rect 8941 1779 8999 1785
rect 9030 1776 9036 1828
rect 9088 1816 9094 1828
rect 9088 1788 9168 1816
rect 9088 1776 9094 1788
rect 3283 1720 3924 1748
rect 3283 1717 3295 1720
rect 3237 1711 3295 1717
rect 4062 1708 4068 1760
rect 4120 1708 4126 1760
rect 4246 1708 4252 1760
rect 4304 1748 4310 1760
rect 4341 1751 4399 1757
rect 4341 1748 4353 1751
rect 4304 1720 4353 1748
rect 4304 1708 4310 1720
rect 4341 1717 4353 1720
rect 4387 1717 4399 1751
rect 4341 1711 4399 1717
rect 5166 1708 5172 1760
rect 5224 1708 5230 1760
rect 5445 1751 5503 1757
rect 5445 1717 5457 1751
rect 5491 1748 5503 1751
rect 5534 1748 5540 1760
rect 5491 1720 5540 1748
rect 5491 1717 5503 1720
rect 5445 1711 5503 1717
rect 5534 1708 5540 1720
rect 5592 1708 5598 1760
rect 5994 1708 6000 1760
rect 6052 1708 6058 1760
rect 6454 1708 6460 1760
rect 6512 1708 6518 1760
rect 6730 1708 6736 1760
rect 6788 1708 6794 1760
rect 7098 1708 7104 1760
rect 7156 1748 7162 1760
rect 7285 1751 7343 1757
rect 7285 1748 7297 1751
rect 7156 1720 7297 1748
rect 7156 1708 7162 1720
rect 7285 1717 7297 1720
rect 7331 1717 7343 1751
rect 7285 1711 7343 1717
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 8389 1751 8447 1757
rect 8389 1748 8401 1751
rect 8260 1720 8401 1748
rect 8260 1708 8266 1720
rect 8389 1717 8401 1720
rect 8435 1717 8447 1751
rect 8389 1711 8447 1717
rect 8662 1708 8668 1760
rect 8720 1708 8726 1760
rect 9140 1748 9168 1788
rect 9490 1776 9496 1828
rect 9548 1776 9554 1828
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 10045 1819 10103 1825
rect 10045 1816 10057 1819
rect 9732 1788 10057 1816
rect 9732 1776 9738 1788
rect 10045 1785 10057 1788
rect 10091 1785 10103 1819
rect 13446 1816 13452 1828
rect 10045 1779 10103 1785
rect 10428 1788 13452 1816
rect 9217 1751 9275 1757
rect 9217 1748 9229 1751
rect 9140 1720 9229 1748
rect 9217 1717 9229 1720
rect 9263 1717 9275 1751
rect 9217 1711 9275 1717
rect 9769 1751 9827 1757
rect 9769 1717 9781 1751
rect 9815 1748 9827 1751
rect 10428 1748 10456 1788
rect 13446 1776 13452 1788
rect 13504 1776 13510 1828
rect 15028 1816 15056 1992
rect 15102 1912 15108 1964
rect 15160 1952 15166 1964
rect 15672 1961 15700 1992
rect 15841 1989 15853 2023
rect 15887 1989 15899 2023
rect 15841 1983 15899 1989
rect 16022 1980 16028 2032
rect 16080 2020 16086 2032
rect 16080 1992 17632 2020
rect 16080 1980 16086 1992
rect 15381 1955 15439 1961
rect 15381 1952 15393 1955
rect 15160 1924 15393 1952
rect 15160 1912 15166 1924
rect 15381 1921 15393 1924
rect 15427 1921 15439 1955
rect 15381 1915 15439 1921
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1921 15715 1955
rect 15657 1915 15715 1921
rect 16114 1912 16120 1964
rect 16172 1952 16178 1964
rect 17604 1961 17632 1992
rect 17770 1980 17776 2032
rect 17828 2020 17834 2032
rect 18049 2023 18107 2029
rect 18049 2020 18061 2023
rect 17828 1992 18061 2020
rect 17828 1980 17834 1992
rect 18049 1989 18061 1992
rect 18095 1989 18107 2023
rect 18248 2020 18276 2048
rect 18601 2023 18659 2029
rect 18601 2020 18613 2023
rect 18248 1992 18613 2020
rect 18049 1983 18107 1989
rect 18601 1989 18613 1992
rect 18647 1989 18659 2023
rect 18601 1983 18659 1989
rect 16485 1955 16543 1961
rect 16485 1952 16497 1955
rect 16172 1924 16497 1952
rect 16172 1912 16178 1924
rect 16485 1921 16497 1924
rect 16531 1921 16543 1955
rect 16485 1915 16543 1921
rect 16945 1955 17003 1961
rect 16945 1921 16957 1955
rect 16991 1921 17003 1955
rect 16945 1915 17003 1921
rect 17589 1955 17647 1961
rect 17589 1921 17601 1955
rect 17635 1921 17647 1955
rect 17589 1915 17647 1921
rect 17865 1955 17923 1961
rect 17865 1921 17877 1955
rect 17911 1921 17923 1955
rect 17865 1915 17923 1921
rect 16960 1884 16988 1915
rect 17880 1884 17908 1915
rect 18414 1912 18420 1964
rect 18472 1912 18478 1964
rect 18708 1952 18736 2060
rect 19150 2048 19156 2100
rect 19208 2048 19214 2100
rect 19242 2048 19248 2100
rect 19300 2088 19306 2100
rect 19300 2060 19840 2088
rect 19300 2048 19306 2060
rect 19168 2020 19196 2048
rect 19705 2023 19763 2029
rect 19705 2020 19717 2023
rect 19168 1992 19717 2020
rect 19705 1989 19717 1992
rect 19751 1989 19763 2023
rect 19705 1983 19763 1989
rect 19153 1955 19211 1961
rect 19153 1952 19165 1955
rect 18708 1924 19165 1952
rect 19153 1921 19165 1924
rect 19199 1921 19211 1955
rect 19812 1952 19840 2060
rect 20346 2048 20352 2100
rect 20404 2088 20410 2100
rect 21082 2088 21088 2100
rect 20404 2060 21088 2088
rect 20404 2048 20410 2060
rect 21082 2048 21088 2060
rect 21140 2048 21146 2100
rect 21174 2048 21180 2100
rect 21232 2088 21238 2100
rect 21453 2091 21511 2097
rect 21453 2088 21465 2091
rect 21232 2060 21465 2088
rect 21232 2048 21238 2060
rect 21453 2057 21465 2060
rect 21499 2057 21511 2091
rect 21453 2051 21511 2057
rect 21634 2048 21640 2100
rect 21692 2088 21698 2100
rect 21821 2091 21879 2097
rect 21821 2088 21833 2091
rect 21692 2060 21833 2088
rect 21692 2048 21698 2060
rect 21821 2057 21833 2060
rect 21867 2057 21879 2091
rect 21821 2051 21879 2057
rect 22278 2048 22284 2100
rect 22336 2048 22342 2100
rect 22741 2091 22799 2097
rect 22741 2057 22753 2091
rect 22787 2088 22799 2091
rect 23106 2088 23112 2100
rect 22787 2060 23112 2088
rect 22787 2057 22799 2060
rect 22741 2051 22799 2057
rect 23106 2048 23112 2060
rect 23164 2048 23170 2100
rect 24026 2048 24032 2100
rect 24084 2048 24090 2100
rect 24394 2048 24400 2100
rect 24452 2048 24458 2100
rect 19886 1980 19892 2032
rect 19944 2020 19950 2032
rect 19944 1992 20484 2020
rect 19944 1980 19950 1992
rect 20257 1955 20315 1961
rect 20257 1952 20269 1955
rect 19812 1924 20269 1952
rect 19153 1915 19211 1921
rect 20257 1921 20269 1924
rect 20303 1921 20315 1955
rect 20257 1915 20315 1921
rect 15212 1856 16988 1884
rect 17052 1856 17908 1884
rect 18432 1884 18460 1912
rect 20456 1884 20484 1992
rect 20622 1980 20628 2032
rect 20680 2020 20686 2032
rect 20809 2023 20867 2029
rect 20809 2020 20821 2023
rect 20680 1992 20821 2020
rect 20680 1980 20686 1992
rect 20809 1989 20821 1992
rect 20855 1989 20867 2023
rect 20809 1983 20867 1989
rect 23382 1980 23388 2032
rect 23440 2020 23446 2032
rect 23440 1992 23980 2020
rect 23440 1980 23446 1992
rect 21082 1912 21088 1964
rect 21140 1912 21146 1964
rect 21266 1912 21272 1964
rect 21324 1952 21330 1964
rect 21637 1955 21695 1961
rect 21637 1952 21649 1955
rect 21324 1924 21649 1952
rect 21324 1912 21330 1924
rect 21637 1921 21649 1924
rect 21683 1921 21695 1955
rect 21637 1915 21695 1921
rect 22002 1912 22008 1964
rect 22060 1912 22066 1964
rect 22097 1955 22155 1961
rect 22097 1921 22109 1955
rect 22143 1921 22155 1955
rect 22097 1915 22155 1921
rect 18432 1856 20208 1884
rect 20456 1856 21312 1884
rect 15212 1825 15240 1856
rect 14200 1788 15056 1816
rect 15197 1819 15255 1825
rect 9815 1720 10456 1748
rect 9815 1717 9827 1720
rect 9769 1711 9827 1717
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 10962 1708 10968 1760
rect 11020 1748 11026 1760
rect 11057 1751 11115 1757
rect 11057 1748 11069 1751
rect 11020 1720 11069 1748
rect 11020 1708 11026 1720
rect 11057 1717 11069 1720
rect 11103 1717 11115 1751
rect 11057 1711 11115 1717
rect 11698 1708 11704 1760
rect 11756 1708 11762 1760
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 12069 1751 12127 1757
rect 12069 1748 12081 1751
rect 11848 1720 12081 1748
rect 11848 1708 11854 1720
rect 12069 1717 12081 1720
rect 12115 1717 12127 1751
rect 12069 1711 12127 1717
rect 12437 1751 12495 1757
rect 12437 1717 12449 1751
rect 12483 1748 12495 1751
rect 12802 1748 12808 1760
rect 12483 1720 12808 1748
rect 12483 1717 12495 1720
rect 12437 1711 12495 1717
rect 12802 1708 12808 1720
rect 12860 1708 12866 1760
rect 12894 1708 12900 1760
rect 12952 1708 12958 1760
rect 13265 1751 13323 1757
rect 13265 1717 13277 1751
rect 13311 1748 13323 1751
rect 13814 1748 13820 1760
rect 13311 1720 13820 1748
rect 13311 1717 13323 1720
rect 13265 1711 13323 1717
rect 13814 1708 13820 1720
rect 13872 1708 13878 1760
rect 13909 1751 13967 1757
rect 13909 1717 13921 1751
rect 13955 1748 13967 1751
rect 14200 1748 14228 1788
rect 15197 1785 15209 1819
rect 15243 1785 15255 1819
rect 15197 1779 15255 1785
rect 15378 1776 15384 1828
rect 15436 1816 15442 1828
rect 17052 1816 17080 1856
rect 15436 1788 17080 1816
rect 15436 1776 15442 1788
rect 17770 1776 17776 1828
rect 17828 1816 17834 1828
rect 17828 1788 19288 1816
rect 17828 1776 17834 1788
rect 13955 1720 14228 1748
rect 13955 1717 13967 1720
rect 13909 1711 13967 1717
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14645 1751 14703 1757
rect 14645 1748 14657 1751
rect 14332 1720 14657 1748
rect 14332 1708 14338 1720
rect 14645 1717 14657 1720
rect 14691 1717 14703 1751
rect 14645 1711 14703 1717
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14792 1720 15025 1748
rect 14792 1708 14798 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15470 1708 15476 1760
rect 15528 1708 15534 1760
rect 15654 1708 15660 1760
rect 15712 1748 15718 1760
rect 15933 1751 15991 1757
rect 15933 1748 15945 1751
rect 15712 1720 15945 1748
rect 15712 1708 15718 1720
rect 15933 1717 15945 1720
rect 15979 1717 15991 1751
rect 15933 1711 15991 1717
rect 16301 1751 16359 1757
rect 16301 1717 16313 1751
rect 16347 1748 16359 1751
rect 16574 1748 16580 1760
rect 16347 1720 16580 1748
rect 16347 1717 16359 1720
rect 16301 1711 16359 1717
rect 16574 1708 16580 1720
rect 16632 1708 16638 1760
rect 16758 1708 16764 1760
rect 16816 1748 16822 1760
rect 17037 1751 17095 1757
rect 17037 1748 17049 1751
rect 16816 1720 17049 1748
rect 16816 1708 16822 1720
rect 17037 1717 17049 1720
rect 17083 1717 17095 1751
rect 17037 1711 17095 1717
rect 17954 1708 17960 1760
rect 18012 1748 18018 1760
rect 18141 1751 18199 1757
rect 18141 1748 18153 1751
rect 18012 1720 18153 1748
rect 18012 1708 18018 1720
rect 18141 1717 18153 1720
rect 18187 1717 18199 1751
rect 18141 1711 18199 1717
rect 18230 1708 18236 1760
rect 18288 1748 18294 1760
rect 19260 1757 19288 1788
rect 19426 1776 19432 1828
rect 19484 1816 19490 1828
rect 20180 1816 20208 1856
rect 21174 1816 21180 1828
rect 19484 1788 19932 1816
rect 20180 1788 21180 1816
rect 19484 1776 19490 1788
rect 18693 1751 18751 1757
rect 18693 1748 18705 1751
rect 18288 1720 18705 1748
rect 18288 1708 18294 1720
rect 18693 1717 18705 1720
rect 18739 1717 18751 1751
rect 18693 1711 18751 1717
rect 19245 1751 19303 1757
rect 19245 1717 19257 1751
rect 19291 1717 19303 1751
rect 19245 1711 19303 1717
rect 19334 1708 19340 1760
rect 19392 1748 19398 1760
rect 19797 1751 19855 1757
rect 19797 1748 19809 1751
rect 19392 1720 19809 1748
rect 19392 1708 19398 1720
rect 19797 1717 19809 1720
rect 19843 1717 19855 1751
rect 19904 1748 19932 1788
rect 21174 1776 21180 1788
rect 21232 1776 21238 1828
rect 20349 1751 20407 1757
rect 20349 1748 20361 1751
rect 19904 1720 20361 1748
rect 19797 1711 19855 1717
rect 20349 1717 20361 1720
rect 20395 1717 20407 1751
rect 20349 1711 20407 1717
rect 20898 1708 20904 1760
rect 20956 1708 20962 1760
rect 21284 1757 21312 1856
rect 21726 1844 21732 1896
rect 21784 1884 21790 1896
rect 22112 1884 22140 1915
rect 22462 1912 22468 1964
rect 22520 1952 22526 1964
rect 22649 1955 22707 1961
rect 22649 1952 22661 1955
rect 22520 1924 22661 1952
rect 22520 1912 22526 1924
rect 22649 1921 22661 1924
rect 22695 1921 22707 1955
rect 22649 1915 22707 1921
rect 22738 1912 22744 1964
rect 22796 1952 22802 1964
rect 22925 1955 22983 1961
rect 22925 1952 22937 1955
rect 22796 1924 22937 1952
rect 22796 1912 22802 1924
rect 22925 1921 22937 1924
rect 22971 1921 22983 1955
rect 22925 1915 22983 1921
rect 23014 1912 23020 1964
rect 23072 1912 23078 1964
rect 23569 1955 23627 1961
rect 23569 1952 23581 1955
rect 23308 1924 23581 1952
rect 21784 1856 22140 1884
rect 21784 1844 21790 1856
rect 22186 1844 22192 1896
rect 22244 1844 22250 1896
rect 22370 1844 22376 1896
rect 22428 1884 22434 1896
rect 23106 1884 23112 1896
rect 22428 1856 23112 1884
rect 22428 1844 22434 1856
rect 23106 1844 23112 1856
rect 23164 1844 23170 1896
rect 21269 1751 21327 1757
rect 21269 1717 21281 1751
rect 21315 1717 21327 1751
rect 22204 1748 22232 1844
rect 22465 1819 22523 1825
rect 22465 1785 22477 1819
rect 22511 1816 22523 1819
rect 23308 1816 23336 1924
rect 23569 1921 23581 1924
rect 23615 1921 23627 1955
rect 23569 1915 23627 1921
rect 23845 1955 23903 1961
rect 23845 1921 23857 1955
rect 23891 1921 23903 1955
rect 23845 1915 23903 1921
rect 23860 1884 23888 1915
rect 23400 1856 23888 1884
rect 23952 1884 23980 1992
rect 24044 1952 24072 2048
rect 24121 1955 24179 1961
rect 24121 1952 24133 1955
rect 24044 1924 24133 1952
rect 24121 1921 24133 1924
rect 24167 1921 24179 1955
rect 24121 1915 24179 1921
rect 24213 1955 24271 1961
rect 24213 1921 24225 1955
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 24228 1884 24256 1915
rect 23952 1856 24256 1884
rect 23400 1825 23428 1856
rect 24302 1844 24308 1896
rect 24360 1844 24366 1896
rect 22511 1788 23336 1816
rect 23385 1819 23443 1825
rect 22511 1785 22523 1788
rect 22465 1779 22523 1785
rect 23385 1785 23397 1819
rect 23431 1785 23443 1819
rect 23385 1779 23443 1785
rect 23474 1776 23480 1828
rect 23532 1816 23538 1828
rect 23750 1816 23756 1828
rect 23532 1788 23756 1816
rect 23532 1776 23538 1788
rect 23750 1776 23756 1788
rect 23808 1776 23814 1828
rect 23937 1819 23995 1825
rect 23937 1785 23949 1819
rect 23983 1816 23995 1819
rect 24320 1816 24348 1844
rect 23983 1788 24348 1816
rect 23983 1785 23995 1788
rect 23937 1779 23995 1785
rect 23201 1751 23259 1757
rect 23201 1748 23213 1751
rect 22204 1720 23213 1748
rect 21269 1711 21327 1717
rect 23201 1717 23213 1720
rect 23247 1717 23259 1751
rect 23201 1711 23259 1717
rect 23661 1751 23719 1757
rect 23661 1717 23673 1751
rect 23707 1748 23719 1751
rect 24118 1748 24124 1760
rect 23707 1720 24124 1748
rect 23707 1717 23719 1720
rect 23661 1711 23719 1717
rect 24118 1708 24124 1720
rect 24176 1708 24182 1760
rect 1104 1658 24840 1680
rect 1104 1606 3917 1658
rect 3969 1606 3981 1658
rect 4033 1606 4045 1658
rect 4097 1606 4109 1658
rect 4161 1606 4173 1658
rect 4225 1606 9851 1658
rect 9903 1606 9915 1658
rect 9967 1606 9979 1658
rect 10031 1606 10043 1658
rect 10095 1606 10107 1658
rect 10159 1606 15785 1658
rect 15837 1606 15849 1658
rect 15901 1606 15913 1658
rect 15965 1606 15977 1658
rect 16029 1606 16041 1658
rect 16093 1606 21719 1658
rect 21771 1606 21783 1658
rect 21835 1606 21847 1658
rect 21899 1606 21911 1658
rect 21963 1606 21975 1658
rect 22027 1606 24840 1658
rect 1104 1584 24840 1606
rect 2590 1504 2596 1556
rect 2648 1504 2654 1556
rect 2866 1504 2872 1556
rect 2924 1504 2930 1556
rect 4338 1544 4344 1556
rect 3344 1516 4344 1544
rect 3234 1408 3240 1420
rect 2700 1380 3240 1408
rect 1394 1300 1400 1352
rect 1452 1300 1458 1352
rect 1486 1300 1492 1352
rect 1544 1340 1550 1352
rect 1673 1343 1731 1349
rect 1673 1340 1685 1343
rect 1544 1312 1685 1340
rect 1544 1300 1550 1312
rect 1673 1309 1685 1312
rect 1719 1309 1731 1343
rect 1673 1303 1731 1309
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 2501 1343 2559 1349
rect 2501 1309 2513 1343
rect 2547 1340 2559 1343
rect 2700 1340 2728 1380
rect 3234 1368 3240 1380
rect 3292 1368 3298 1420
rect 2547 1312 2728 1340
rect 2547 1309 2559 1312
rect 2501 1303 2559 1309
rect 1412 1204 1440 1300
rect 1780 1272 1808 1303
rect 2240 1272 2268 1303
rect 2774 1300 2780 1352
rect 2832 1300 2838 1352
rect 3050 1300 3056 1352
rect 3108 1300 3114 1352
rect 3344 1349 3372 1516
rect 4338 1504 4344 1516
rect 4396 1504 4402 1556
rect 5077 1547 5135 1553
rect 5077 1513 5089 1547
rect 5123 1544 5135 1547
rect 5902 1544 5908 1556
rect 5123 1516 5908 1544
rect 5123 1513 5135 1516
rect 5077 1507 5135 1513
rect 5902 1504 5908 1516
rect 5960 1504 5966 1556
rect 5994 1504 6000 1556
rect 6052 1504 6058 1556
rect 6181 1547 6239 1553
rect 6181 1513 6193 1547
rect 6227 1544 6239 1547
rect 6914 1544 6920 1556
rect 6227 1516 6920 1544
rect 6227 1513 6239 1516
rect 6181 1507 6239 1513
rect 6914 1504 6920 1516
rect 6972 1504 6978 1556
rect 7098 1504 7104 1556
rect 7156 1544 7162 1556
rect 7156 1516 13768 1544
rect 7156 1504 7162 1516
rect 3421 1479 3479 1485
rect 3421 1445 3433 1479
rect 3467 1476 3479 1479
rect 3467 1448 4292 1476
rect 3467 1445 3479 1448
rect 3421 1439 3479 1445
rect 4264 1408 4292 1448
rect 6012 1408 6040 1504
rect 6641 1479 6699 1485
rect 6641 1445 6653 1479
rect 6687 1445 6699 1479
rect 6641 1439 6699 1445
rect 7193 1479 7251 1485
rect 7193 1445 7205 1479
rect 7239 1476 7251 1479
rect 7469 1479 7527 1485
rect 7239 1448 7420 1476
rect 7239 1445 7251 1448
rect 7193 1439 7251 1445
rect 3528 1380 4108 1408
rect 4264 1380 4384 1408
rect 3528 1352 3556 1380
rect 3329 1343 3387 1349
rect 3329 1309 3341 1343
rect 3375 1309 3387 1343
rect 3329 1303 3387 1309
rect 3510 1300 3516 1352
rect 3568 1300 3574 1352
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1340 3663 1343
rect 3878 1340 3884 1352
rect 3651 1312 3884 1340
rect 3651 1309 3663 1312
rect 3605 1303 3663 1309
rect 3878 1300 3884 1312
rect 3936 1300 3942 1352
rect 3973 1343 4031 1349
rect 3973 1309 3985 1343
rect 4019 1309 4031 1343
rect 4080 1340 4108 1380
rect 4249 1343 4307 1349
rect 4249 1340 4261 1343
rect 4080 1312 4261 1340
rect 3973 1303 4031 1309
rect 4249 1309 4261 1312
rect 4295 1309 4307 1343
rect 4356 1340 4384 1380
rect 4816 1380 5028 1408
rect 4525 1343 4583 1349
rect 4525 1340 4537 1343
rect 4356 1312 4537 1340
rect 4249 1303 4307 1309
rect 4525 1309 4537 1312
rect 4571 1309 4583 1343
rect 4525 1303 4583 1309
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1340 4675 1343
rect 4816 1340 4844 1380
rect 4663 1312 4844 1340
rect 4893 1343 4951 1349
rect 4663 1309 4675 1312
rect 4617 1303 4675 1309
rect 4893 1309 4905 1343
rect 4939 1309 4951 1343
rect 4893 1303 4951 1309
rect 2682 1272 2688 1284
rect 1780 1244 2176 1272
rect 2240 1244 2688 1272
rect 1489 1207 1547 1213
rect 1489 1204 1501 1207
rect 1412 1176 1501 1204
rect 1489 1173 1501 1176
rect 1535 1173 1547 1207
rect 1489 1167 1547 1173
rect 1670 1164 1676 1216
rect 1728 1204 1734 1216
rect 1949 1207 2007 1213
rect 1949 1204 1961 1207
rect 1728 1176 1961 1204
rect 1728 1164 1734 1176
rect 1949 1173 1961 1176
rect 1995 1173 2007 1207
rect 1949 1167 2007 1173
rect 2038 1164 2044 1216
rect 2096 1164 2102 1216
rect 2148 1204 2176 1244
rect 2682 1232 2688 1244
rect 2740 1232 2746 1284
rect 3988 1272 4016 1303
rect 4908 1272 4936 1303
rect 3160 1244 4016 1272
rect 4080 1244 4936 1272
rect 5000 1272 5028 1380
rect 5736 1380 6040 1408
rect 6656 1408 6684 1439
rect 7392 1408 7420 1448
rect 7469 1445 7481 1479
rect 7515 1476 7527 1479
rect 8478 1476 8484 1488
rect 7515 1448 8484 1476
rect 7515 1445 7527 1448
rect 7469 1439 7527 1445
rect 8478 1436 8484 1448
rect 8536 1436 8542 1488
rect 8570 1436 8576 1488
rect 8628 1436 8634 1488
rect 8938 1436 8944 1488
rect 8996 1476 9002 1488
rect 11974 1476 11980 1488
rect 8996 1448 9996 1476
rect 8996 1436 9002 1448
rect 7834 1408 7840 1420
rect 6656 1380 7236 1408
rect 7392 1380 7840 1408
rect 5166 1300 5172 1352
rect 5224 1340 5230 1352
rect 5353 1343 5411 1349
rect 5353 1340 5365 1343
rect 5224 1312 5365 1340
rect 5224 1300 5230 1312
rect 5353 1309 5365 1312
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 5534 1300 5540 1352
rect 5592 1340 5598 1352
rect 5736 1349 5764 1380
rect 5629 1343 5687 1349
rect 5629 1340 5641 1343
rect 5592 1312 5641 1340
rect 5592 1300 5598 1312
rect 5629 1309 5641 1312
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5997 1343 6055 1349
rect 5997 1309 6009 1343
rect 6043 1340 6055 1343
rect 6454 1340 6460 1352
rect 6043 1312 6460 1340
rect 6043 1309 6055 1312
rect 5997 1303 6055 1309
rect 6454 1300 6460 1312
rect 6512 1300 6518 1352
rect 6549 1343 6607 1349
rect 6549 1309 6561 1343
rect 6595 1340 6607 1343
rect 6730 1340 6736 1352
rect 6595 1312 6736 1340
rect 6595 1309 6607 1312
rect 6549 1303 6607 1309
rect 6730 1300 6736 1312
rect 6788 1300 6794 1352
rect 6822 1300 6828 1352
rect 6880 1300 6886 1352
rect 6914 1300 6920 1352
rect 6972 1300 6978 1352
rect 7006 1300 7012 1352
rect 7064 1340 7070 1352
rect 7101 1343 7159 1349
rect 7101 1340 7113 1343
rect 7064 1312 7113 1340
rect 7064 1300 7070 1312
rect 7101 1309 7113 1312
rect 7147 1309 7159 1343
rect 7208 1340 7236 1380
rect 7834 1368 7840 1380
rect 7892 1368 7898 1420
rect 8386 1408 8392 1420
rect 8128 1380 8392 1408
rect 7377 1343 7435 1349
rect 7377 1340 7389 1343
rect 7208 1312 7389 1340
rect 7101 1303 7159 1309
rect 7377 1309 7389 1312
rect 7423 1309 7435 1343
rect 7377 1303 7435 1309
rect 7653 1343 7711 1349
rect 7653 1309 7665 1343
rect 7699 1309 7711 1343
rect 7653 1303 7711 1309
rect 7929 1343 7987 1349
rect 7929 1309 7941 1343
rect 7975 1340 7987 1343
rect 8128 1340 8156 1380
rect 8386 1368 8392 1380
rect 8444 1368 8450 1420
rect 9048 1380 9720 1408
rect 7975 1312 8156 1340
rect 7975 1309 7987 1312
rect 7929 1303 7987 1309
rect 6932 1272 6960 1300
rect 7668 1272 7696 1303
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8478 1300 8484 1352
rect 8536 1300 8542 1352
rect 9048 1349 9076 1380
rect 9033 1343 9091 1349
rect 8757 1319 8815 1325
rect 8757 1285 8769 1319
rect 8803 1316 8815 1319
rect 8803 1288 8892 1316
rect 9033 1309 9045 1343
rect 9079 1309 9091 1343
rect 9033 1303 9091 1309
rect 9214 1300 9220 1352
rect 9272 1300 9278 1352
rect 9490 1300 9496 1352
rect 9548 1300 9554 1352
rect 9585 1343 9643 1349
rect 9585 1309 9597 1343
rect 9631 1309 9643 1343
rect 9692 1340 9720 1380
rect 9766 1340 9772 1352
rect 9692 1312 9772 1340
rect 9585 1303 9643 1309
rect 8803 1285 8815 1288
rect 5000 1244 5580 1272
rect 2222 1204 2228 1216
rect 2148 1176 2228 1204
rect 2222 1164 2228 1176
rect 2280 1164 2286 1216
rect 2314 1164 2320 1216
rect 2372 1164 2378 1216
rect 3160 1213 3188 1244
rect 3145 1207 3203 1213
rect 3145 1173 3157 1207
rect 3191 1173 3203 1207
rect 3145 1167 3203 1173
rect 3326 1164 3332 1216
rect 3384 1204 3390 1216
rect 3510 1204 3516 1216
rect 3384 1176 3516 1204
rect 3384 1164 3390 1176
rect 3510 1164 3516 1176
rect 3568 1164 3574 1216
rect 3789 1207 3847 1213
rect 3789 1173 3801 1207
rect 3835 1204 3847 1207
rect 3970 1204 3976 1216
rect 3835 1176 3976 1204
rect 3835 1173 3847 1176
rect 3789 1167 3847 1173
rect 3970 1164 3976 1176
rect 4028 1164 4034 1216
rect 4080 1213 4108 1244
rect 5552 1216 5580 1244
rect 5920 1244 6960 1272
rect 7116 1244 7696 1272
rect 4065 1207 4123 1213
rect 4065 1173 4077 1207
rect 4111 1173 4123 1207
rect 4065 1167 4123 1173
rect 4338 1164 4344 1216
rect 4396 1164 4402 1216
rect 4798 1164 4804 1216
rect 4856 1164 4862 1216
rect 5166 1164 5172 1216
rect 5224 1164 5230 1216
rect 5442 1164 5448 1216
rect 5500 1164 5506 1216
rect 5534 1164 5540 1216
rect 5592 1164 5598 1216
rect 5920 1213 5948 1244
rect 5905 1207 5963 1213
rect 5905 1173 5917 1207
rect 5951 1173 5963 1207
rect 5905 1167 5963 1173
rect 6362 1164 6368 1216
rect 6420 1164 6426 1216
rect 6917 1207 6975 1213
rect 6917 1173 6929 1207
rect 6963 1204 6975 1207
rect 7116 1204 7144 1244
rect 7834 1232 7840 1284
rect 7892 1272 7898 1284
rect 8757 1279 8815 1285
rect 8864 1272 8892 1288
rect 9122 1272 9128 1284
rect 7892 1244 8064 1272
rect 8864 1244 9128 1272
rect 7892 1232 7898 1244
rect 6963 1176 7144 1204
rect 6963 1173 6975 1176
rect 6917 1167 6975 1173
rect 7190 1164 7196 1216
rect 7248 1204 7254 1216
rect 7650 1204 7656 1216
rect 7248 1176 7656 1204
rect 7248 1164 7254 1176
rect 7650 1164 7656 1176
rect 7708 1164 7714 1216
rect 7745 1207 7803 1213
rect 7745 1173 7757 1207
rect 7791 1204 7803 1207
rect 7926 1204 7932 1216
rect 7791 1176 7932 1204
rect 7791 1173 7803 1176
rect 7745 1167 7803 1173
rect 7926 1164 7932 1176
rect 7984 1164 7990 1216
rect 8036 1213 8064 1244
rect 9122 1232 9128 1244
rect 9180 1232 9186 1284
rect 9232 1272 9260 1300
rect 9600 1272 9628 1303
rect 9766 1300 9772 1312
rect 9824 1300 9830 1352
rect 9968 1349 9996 1448
rect 11440 1448 11980 1476
rect 11054 1368 11060 1420
rect 11112 1368 11118 1420
rect 9953 1343 10011 1349
rect 9953 1309 9965 1343
rect 9999 1309 10011 1343
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 9953 1303 10011 1309
rect 10060 1312 10333 1340
rect 9232 1244 9628 1272
rect 9858 1232 9864 1284
rect 9916 1272 9922 1284
rect 10060 1272 10088 1312
rect 10321 1309 10333 1312
rect 10367 1309 10379 1343
rect 10321 1303 10379 1309
rect 10686 1272 10692 1284
rect 9916 1244 10088 1272
rect 10152 1244 10692 1272
rect 9916 1232 9922 1244
rect 8021 1207 8079 1213
rect 8021 1173 8033 1207
rect 8067 1173 8079 1207
rect 8021 1167 8079 1173
rect 8202 1164 8208 1216
rect 8260 1204 8266 1216
rect 8297 1207 8355 1213
rect 8297 1204 8309 1207
rect 8260 1176 8309 1204
rect 8260 1164 8266 1176
rect 8297 1173 8309 1176
rect 8343 1173 8355 1207
rect 8297 1167 8355 1173
rect 9214 1164 9220 1216
rect 9272 1164 9278 1216
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1204 9367 1207
rect 9674 1204 9680 1216
rect 9355 1176 9680 1204
rect 9355 1173 9367 1176
rect 9309 1167 9367 1173
rect 9674 1164 9680 1176
rect 9732 1164 9738 1216
rect 9769 1207 9827 1213
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10042 1204 10048 1216
rect 9815 1176 10048 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10042 1164 10048 1176
rect 10100 1164 10106 1216
rect 10152 1213 10180 1244
rect 10686 1232 10692 1244
rect 10744 1232 10750 1284
rect 10778 1232 10784 1284
rect 10836 1232 10842 1284
rect 10137 1207 10195 1213
rect 10137 1173 10149 1207
rect 10183 1173 10195 1207
rect 10137 1167 10195 1173
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 11146 1204 11152 1216
rect 10551 1176 11152 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 11146 1164 11152 1176
rect 11204 1164 11210 1216
rect 11440 1204 11468 1448
rect 11974 1436 11980 1448
rect 12032 1436 12038 1488
rect 12526 1436 12532 1488
rect 12584 1476 12590 1488
rect 13740 1476 13768 1516
rect 13814 1504 13820 1556
rect 13872 1544 13878 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13872 1516 14289 1544
rect 13872 1504 13878 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14918 1504 14924 1556
rect 14976 1544 14982 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 14976 1516 15393 1544
rect 14976 1504 14982 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 16301 1547 16359 1553
rect 16301 1513 16313 1547
rect 16347 1544 16359 1547
rect 16482 1544 16488 1556
rect 16347 1516 16488 1544
rect 16347 1513 16359 1516
rect 16301 1507 16359 1513
rect 12584 1448 12664 1476
rect 13740 1448 14320 1476
rect 12584 1436 12590 1448
rect 11514 1368 11520 1420
rect 11572 1408 11578 1420
rect 11572 1380 12572 1408
rect 11572 1368 11578 1380
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11793 1343 11851 1349
rect 11793 1309 11805 1343
rect 11839 1309 11851 1343
rect 12434 1340 12440 1352
rect 11793 1303 11851 1309
rect 11992 1312 12440 1340
rect 11808 1272 11836 1303
rect 11624 1244 11836 1272
rect 11624 1216 11652 1244
rect 11517 1207 11575 1213
rect 11517 1204 11529 1207
rect 11440 1176 11529 1204
rect 11517 1173 11529 1176
rect 11563 1173 11575 1207
rect 11517 1167 11575 1173
rect 11606 1164 11612 1216
rect 11664 1164 11670 1216
rect 11992 1213 12020 1312
rect 12434 1300 12440 1312
rect 12492 1300 12498 1352
rect 12253 1275 12311 1281
rect 12253 1272 12265 1275
rect 12084 1244 12265 1272
rect 12084 1216 12112 1244
rect 12253 1241 12265 1244
rect 12299 1241 12311 1275
rect 12544 1272 12572 1380
rect 12636 1340 12664 1448
rect 12802 1368 12808 1420
rect 12860 1408 12866 1420
rect 14292 1408 14320 1448
rect 15286 1436 15292 1488
rect 15344 1476 15350 1488
rect 15948 1476 15976 1507
rect 16482 1504 16488 1516
rect 16540 1504 16546 1556
rect 16853 1547 16911 1553
rect 16853 1513 16865 1547
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1513 17463 1547
rect 17405 1507 17463 1513
rect 15344 1448 15976 1476
rect 15344 1436 15350 1448
rect 16022 1436 16028 1488
rect 16080 1476 16086 1488
rect 16868 1476 16896 1507
rect 16080 1448 16896 1476
rect 16080 1436 16086 1448
rect 15378 1408 15384 1420
rect 12860 1380 14228 1408
rect 14292 1380 15384 1408
rect 12860 1368 12866 1380
rect 12897 1343 12955 1349
rect 12897 1340 12909 1343
rect 12636 1312 12909 1340
rect 12897 1309 12909 1312
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 13265 1343 13323 1349
rect 13265 1309 13277 1343
rect 13311 1309 13323 1343
rect 13265 1303 13323 1309
rect 13280 1272 13308 1303
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 14200 1349 14228 1380
rect 15378 1368 15384 1380
rect 15436 1368 15442 1420
rect 16206 1368 16212 1420
rect 16264 1408 16270 1420
rect 17420 1408 17448 1507
rect 17586 1504 17592 1556
rect 17644 1544 17650 1556
rect 18509 1547 18567 1553
rect 18509 1544 18521 1547
rect 17644 1516 18521 1544
rect 17644 1504 17650 1516
rect 18509 1513 18521 1516
rect 18555 1513 18567 1547
rect 19429 1547 19487 1553
rect 19429 1544 19441 1547
rect 18509 1507 18567 1513
rect 18616 1516 19441 1544
rect 18616 1476 18644 1516
rect 19429 1513 19441 1516
rect 19475 1513 19487 1547
rect 19429 1507 19487 1513
rect 19794 1504 19800 1556
rect 19852 1544 19858 1556
rect 21085 1547 21143 1553
rect 21085 1544 21097 1547
rect 19852 1516 21097 1544
rect 19852 1504 19858 1516
rect 21085 1513 21097 1516
rect 21131 1513 21143 1547
rect 21085 1507 21143 1513
rect 21174 1504 21180 1556
rect 21232 1544 21238 1556
rect 21453 1547 21511 1553
rect 21453 1544 21465 1547
rect 21232 1516 21465 1544
rect 21232 1504 21238 1516
rect 21453 1513 21465 1516
rect 21499 1513 21511 1547
rect 21453 1507 21511 1513
rect 22094 1504 22100 1556
rect 22152 1544 22158 1556
rect 23201 1547 23259 1553
rect 23201 1544 23213 1547
rect 22152 1516 23213 1544
rect 22152 1504 22158 1516
rect 23201 1513 23213 1516
rect 23247 1513 23259 1547
rect 23201 1507 23259 1513
rect 23308 1516 23612 1544
rect 17604 1448 18644 1476
rect 17604 1420 17632 1448
rect 18690 1436 18696 1488
rect 18748 1476 18754 1488
rect 20073 1479 20131 1485
rect 20073 1476 20085 1479
rect 18748 1448 20085 1476
rect 18748 1436 18754 1448
rect 20073 1445 20085 1448
rect 20119 1445 20131 1479
rect 20073 1439 20131 1445
rect 20625 1479 20683 1485
rect 20625 1445 20637 1479
rect 20671 1445 20683 1479
rect 20625 1439 20683 1445
rect 16264 1380 17448 1408
rect 16264 1368 16270 1380
rect 17586 1368 17592 1420
rect 17644 1368 17650 1420
rect 18138 1368 18144 1420
rect 18196 1368 18202 1420
rect 18598 1368 18604 1420
rect 18656 1408 18662 1420
rect 20640 1408 20668 1439
rect 21542 1436 21548 1488
rect 21600 1476 21606 1488
rect 21600 1448 21680 1476
rect 21600 1436 21606 1448
rect 18656 1380 20668 1408
rect 18656 1368 18662 1380
rect 21450 1368 21456 1420
rect 21508 1408 21514 1420
rect 21652 1408 21680 1448
rect 21818 1436 21824 1488
rect 21876 1436 21882 1488
rect 22002 1436 22008 1488
rect 22060 1476 22066 1488
rect 23308 1476 23336 1516
rect 23474 1476 23480 1488
rect 22060 1448 23336 1476
rect 23400 1448 23480 1476
rect 22060 1436 22066 1448
rect 21508 1380 21588 1408
rect 21652 1380 22692 1408
rect 21508 1368 21514 1380
rect 14185 1343 14243 1349
rect 14185 1309 14197 1343
rect 14231 1309 14243 1343
rect 14185 1303 14243 1309
rect 14642 1300 14648 1352
rect 14700 1300 14706 1352
rect 15289 1343 15347 1349
rect 15289 1309 15301 1343
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 12544 1244 13308 1272
rect 13924 1272 13952 1300
rect 15304 1272 15332 1303
rect 15470 1300 15476 1352
rect 15528 1340 15534 1352
rect 15841 1343 15899 1349
rect 15841 1340 15853 1343
rect 15528 1312 15853 1340
rect 15528 1300 15534 1312
rect 15841 1309 15853 1312
rect 15887 1309 15899 1343
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 15841 1303 15899 1309
rect 15948 1312 16497 1340
rect 13924 1244 15332 1272
rect 12253 1235 12311 1241
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1173 12035 1207
rect 11977 1167 12035 1173
rect 12066 1164 12072 1216
rect 12124 1164 12130 1216
rect 12342 1164 12348 1216
rect 12400 1164 12406 1216
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13446 1164 13452 1216
rect 13504 1164 13510 1216
rect 13998 1164 14004 1216
rect 14056 1204 14062 1216
rect 14829 1207 14887 1213
rect 14829 1204 14841 1207
rect 14056 1176 14841 1204
rect 14056 1164 14062 1176
rect 14829 1173 14841 1176
rect 14875 1173 14887 1207
rect 14829 1167 14887 1173
rect 15010 1164 15016 1216
rect 15068 1204 15074 1216
rect 15948 1204 15976 1312
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16485 1303 16543 1309
rect 16574 1300 16580 1352
rect 16632 1340 16638 1352
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16632 1312 16773 1340
rect 16632 1300 16638 1312
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16761 1303 16819 1309
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 17865 1343 17923 1349
rect 17865 1340 17877 1343
rect 16908 1312 17877 1340
rect 16908 1300 16914 1312
rect 17865 1309 17877 1312
rect 17911 1309 17923 1343
rect 18156 1340 18184 1368
rect 19061 1343 19119 1349
rect 19061 1340 19073 1343
rect 18156 1312 19073 1340
rect 17865 1303 17923 1309
rect 19061 1309 19073 1312
rect 19107 1309 19119 1343
rect 19889 1343 19947 1349
rect 19889 1340 19901 1343
rect 19061 1303 19119 1309
rect 19168 1312 19901 1340
rect 16390 1232 16396 1284
rect 16448 1272 16454 1284
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 16448 1244 17325 1272
rect 16448 1232 16454 1244
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17313 1235 17371 1241
rect 17402 1232 17408 1284
rect 17460 1272 17466 1284
rect 18417 1275 18475 1281
rect 18417 1272 18429 1275
rect 17460 1244 18429 1272
rect 17460 1232 17466 1244
rect 18417 1241 18429 1244
rect 18463 1241 18475 1275
rect 18417 1235 18475 1241
rect 18506 1232 18512 1284
rect 18564 1272 18570 1284
rect 18690 1272 18696 1284
rect 18564 1244 18696 1272
rect 18564 1232 18570 1244
rect 18690 1232 18696 1244
rect 18748 1232 18754 1284
rect 19168 1272 19196 1312
rect 19889 1309 19901 1312
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20993 1343 21051 1349
rect 20993 1340 21005 1343
rect 20036 1312 21005 1340
rect 20036 1300 20042 1312
rect 20993 1309 21005 1312
rect 21039 1309 21051 1343
rect 21560 1340 21588 1380
rect 21637 1343 21695 1349
rect 21637 1340 21649 1343
rect 21560 1312 21649 1340
rect 20993 1303 21051 1309
rect 21637 1309 21649 1312
rect 21683 1309 21695 1343
rect 21637 1303 21695 1309
rect 21726 1300 21732 1352
rect 21784 1340 21790 1352
rect 22005 1343 22063 1349
rect 22005 1340 22017 1343
rect 21784 1312 22017 1340
rect 21784 1300 21790 1312
rect 22005 1309 22017 1312
rect 22051 1309 22063 1343
rect 22005 1303 22063 1309
rect 22097 1343 22155 1349
rect 22097 1309 22109 1343
rect 22143 1309 22155 1343
rect 22373 1343 22431 1349
rect 22373 1340 22385 1343
rect 22097 1303 22155 1309
rect 22204 1312 22385 1340
rect 18892 1244 19196 1272
rect 19337 1275 19395 1281
rect 15068 1176 15976 1204
rect 15068 1164 15074 1176
rect 16482 1164 16488 1216
rect 16540 1204 16546 1216
rect 18892 1213 18920 1244
rect 19337 1241 19349 1275
rect 19383 1272 19395 1275
rect 19610 1272 19616 1284
rect 19383 1244 19616 1272
rect 19383 1241 19395 1244
rect 19337 1235 19395 1241
rect 19610 1232 19616 1244
rect 19668 1232 19674 1284
rect 20441 1275 20499 1281
rect 20441 1241 20453 1275
rect 20487 1241 20499 1275
rect 22112 1272 22140 1303
rect 20441 1235 20499 1241
rect 21744 1244 22140 1272
rect 17957 1207 18015 1213
rect 17957 1204 17969 1207
rect 16540 1176 17969 1204
rect 16540 1164 16546 1176
rect 17957 1173 17969 1176
rect 18003 1173 18015 1207
rect 17957 1167 18015 1173
rect 18877 1207 18935 1213
rect 18877 1173 18889 1207
rect 18923 1173 18935 1207
rect 18877 1167 18935 1173
rect 19058 1164 19064 1216
rect 19116 1204 19122 1216
rect 20456 1204 20484 1235
rect 19116 1176 20484 1204
rect 19116 1164 19122 1176
rect 20530 1164 20536 1216
rect 20588 1204 20594 1216
rect 21744 1204 21772 1244
rect 20588 1176 21772 1204
rect 20588 1164 20594 1176
rect 21910 1164 21916 1216
rect 21968 1204 21974 1216
rect 22204 1204 22232 1312
rect 22373 1309 22385 1312
rect 22419 1309 22431 1343
rect 22373 1303 22431 1309
rect 22554 1300 22560 1352
rect 22612 1300 22618 1352
rect 22664 1349 22692 1380
rect 22649 1343 22707 1349
rect 22649 1309 22661 1343
rect 22695 1309 22707 1343
rect 22649 1303 22707 1309
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 22922 1300 22928 1352
rect 22980 1300 22986 1352
rect 23400 1349 23428 1448
rect 23474 1436 23480 1448
rect 23532 1436 23538 1488
rect 23584 1408 23612 1516
rect 23750 1436 23756 1488
rect 23808 1476 23814 1488
rect 25314 1476 25320 1488
rect 23808 1448 25320 1476
rect 23808 1436 23814 1448
rect 25314 1436 25320 1448
rect 25372 1436 25378 1488
rect 23492 1380 23612 1408
rect 23492 1349 23520 1380
rect 23385 1343 23443 1349
rect 23385 1309 23397 1343
rect 23431 1309 23443 1343
rect 23385 1303 23443 1309
rect 23477 1343 23535 1349
rect 23477 1309 23489 1343
rect 23523 1309 23535 1343
rect 23477 1303 23535 1309
rect 23753 1343 23811 1349
rect 23753 1309 23765 1343
rect 23799 1340 23811 1343
rect 23842 1340 23848 1352
rect 23799 1312 23848 1340
rect 23799 1309 23811 1312
rect 23753 1303 23811 1309
rect 23842 1300 23848 1312
rect 23900 1300 23906 1352
rect 24026 1300 24032 1352
rect 24084 1300 24090 1352
rect 21968 1176 22232 1204
rect 21968 1164 21974 1176
rect 22278 1164 22284 1216
rect 22336 1164 22342 1216
rect 22572 1213 22600 1300
rect 22557 1207 22615 1213
rect 22557 1173 22569 1207
rect 22603 1173 22615 1207
rect 22756 1204 22784 1300
rect 22833 1207 22891 1213
rect 22833 1204 22845 1207
rect 22756 1176 22845 1204
rect 22557 1167 22615 1173
rect 22833 1173 22845 1176
rect 22879 1173 22891 1207
rect 22833 1167 22891 1173
rect 23106 1164 23112 1216
rect 23164 1164 23170 1216
rect 23658 1164 23664 1216
rect 23716 1164 23722 1216
rect 23750 1164 23756 1216
rect 23808 1204 23814 1216
rect 23937 1207 23995 1213
rect 23937 1204 23949 1207
rect 23808 1176 23949 1204
rect 23808 1164 23814 1176
rect 23937 1173 23949 1176
rect 23983 1173 23995 1207
rect 23937 1167 23995 1173
rect 24213 1207 24271 1213
rect 24213 1173 24225 1207
rect 24259 1204 24271 1207
rect 24302 1204 24308 1216
rect 24259 1176 24308 1204
rect 24259 1173 24271 1176
rect 24213 1167 24271 1173
rect 24302 1164 24308 1176
rect 24360 1164 24366 1216
rect 1104 1114 25000 1136
rect 1104 1062 6884 1114
rect 6936 1062 6948 1114
rect 7000 1062 7012 1114
rect 7064 1062 7076 1114
rect 7128 1062 7140 1114
rect 7192 1062 12818 1114
rect 12870 1062 12882 1114
rect 12934 1062 12946 1114
rect 12998 1062 13010 1114
rect 13062 1062 13074 1114
rect 13126 1062 18752 1114
rect 18804 1062 18816 1114
rect 18868 1062 18880 1114
rect 18932 1062 18944 1114
rect 18996 1062 19008 1114
rect 19060 1062 24686 1114
rect 24738 1062 24750 1114
rect 24802 1062 24814 1114
rect 24866 1062 24878 1114
rect 24930 1062 24942 1114
rect 24994 1062 25000 1114
rect 1104 1040 25000 1062
rect 2038 960 2044 1012
rect 2096 1000 2102 1012
rect 2096 972 2774 1000
rect 2096 960 2102 972
rect 2314 892 2320 944
rect 2372 892 2378 944
rect 2746 932 2774 972
rect 5442 960 5448 1012
rect 5500 1000 5506 1012
rect 10778 1000 10784 1012
rect 5500 972 10784 1000
rect 5500 960 5506 972
rect 10778 960 10784 972
rect 10836 960 10842 1012
rect 10870 960 10876 1012
rect 10928 1000 10934 1012
rect 16390 1000 16396 1012
rect 10928 972 16396 1000
rect 10928 960 10934 972
rect 16390 960 16396 972
rect 16448 960 16454 1012
rect 16942 960 16948 1012
rect 17000 1000 17006 1012
rect 19610 1000 19616 1012
rect 17000 972 19616 1000
rect 17000 960 17006 972
rect 19610 960 19616 972
rect 19668 960 19674 1012
rect 21910 960 21916 1012
rect 21968 1000 21974 1012
rect 23106 1000 23112 1012
rect 21968 972 23112 1000
rect 21968 960 21974 972
rect 23106 960 23112 972
rect 23164 960 23170 1012
rect 23658 960 23664 1012
rect 23716 960 23722 1012
rect 24302 960 24308 1012
rect 24360 960 24366 1012
rect 8570 932 8576 944
rect 2746 904 8576 932
rect 8570 892 8576 904
rect 8628 892 8634 944
rect 9674 892 9680 944
rect 9732 932 9738 944
rect 14642 932 14648 944
rect 9732 904 12434 932
rect 9732 892 9738 904
rect 2332 796 2360 892
rect 6362 824 6368 876
rect 6420 864 6426 876
rect 11606 864 11612 876
rect 6420 836 11612 864
rect 6420 824 6426 836
rect 11606 824 11612 836
rect 11664 824 11670 876
rect 2332 768 2774 796
rect 2746 592 2774 768
rect 3418 756 3424 808
rect 3476 796 3482 808
rect 6730 796 6736 808
rect 3476 768 6736 796
rect 3476 756 3482 768
rect 6730 756 6736 768
rect 6788 756 6794 808
rect 7558 756 7564 808
rect 7616 756 7622 808
rect 8018 756 8024 808
rect 8076 796 8082 808
rect 12406 796 12434 904
rect 13556 904 14648 932
rect 13556 796 13584 904
rect 14642 892 14648 904
rect 14700 892 14706 944
rect 16666 892 16672 944
rect 16724 932 16730 944
rect 23676 932 23704 960
rect 16724 904 23704 932
rect 16724 892 16730 904
rect 14182 824 14188 876
rect 14240 864 14246 876
rect 24320 864 24348 960
rect 14240 836 24348 864
rect 14240 824 14246 836
rect 8076 768 10088 796
rect 12406 768 13584 796
rect 8076 756 8082 768
rect 3970 688 3976 740
rect 4028 728 4034 740
rect 7576 728 7604 756
rect 4028 700 7604 728
rect 4028 688 4034 700
rect 9214 620 9220 672
rect 9272 620 9278 672
rect 10060 660 10088 768
rect 20898 756 20904 808
rect 20956 796 20962 808
rect 21726 796 21732 808
rect 20956 768 21732 796
rect 20956 756 20962 768
rect 21726 756 21732 768
rect 21784 756 21790 808
rect 22278 796 22284 808
rect 22066 768 22284 796
rect 12434 688 12440 740
rect 12492 728 12498 740
rect 12894 728 12900 740
rect 12492 700 12900 728
rect 12492 688 12498 700
rect 12894 688 12900 700
rect 12952 688 12958 740
rect 14458 688 14464 740
rect 14516 728 14522 740
rect 22066 728 22094 768
rect 22278 756 22284 768
rect 22336 756 22342 808
rect 22922 756 22928 808
rect 22980 756 22986 808
rect 23290 756 23296 808
rect 23348 796 23354 808
rect 25590 796 25596 808
rect 23348 768 25596 796
rect 23348 756 23354 768
rect 25590 756 25596 768
rect 25648 756 25654 808
rect 14516 700 22094 728
rect 14516 688 14522 700
rect 13538 660 13544 672
rect 10060 632 13544 660
rect 13538 620 13544 632
rect 13596 620 13602 672
rect 15194 620 15200 672
rect 15252 660 15258 672
rect 15252 632 16436 660
rect 15252 620 15258 632
rect 6914 592 6920 604
rect 2746 564 6920 592
rect 6914 552 6920 564
rect 6972 552 6978 604
rect 9232 592 9260 620
rect 16114 592 16120 604
rect 9232 564 16120 592
rect 16114 552 16120 564
rect 16172 552 16178 604
rect 16408 592 16436 632
rect 20346 620 20352 672
rect 20404 660 20410 672
rect 21266 660 21272 672
rect 20404 632 21272 660
rect 20404 620 20410 632
rect 21266 620 21272 632
rect 21324 620 21330 672
rect 21450 620 21456 672
rect 21508 660 21514 672
rect 22940 660 22968 756
rect 23566 688 23572 740
rect 23624 688 23630 740
rect 21508 632 22968 660
rect 21508 620 21514 632
rect 23584 592 23612 688
rect 16408 564 23612 592
rect 2774 484 2780 536
rect 2832 524 2838 536
rect 3510 524 3516 536
rect 2832 496 3516 524
rect 2832 484 2838 496
rect 3510 484 3516 496
rect 3568 484 3574 536
rect 3602 484 3608 536
rect 3660 484 3666 536
rect 5166 484 5172 536
rect 5224 524 5230 536
rect 9858 524 9864 536
rect 5224 496 9864 524
rect 5224 484 5230 496
rect 9858 484 9864 496
rect 9916 484 9922 536
rect 11238 484 11244 536
rect 11296 484 11302 536
rect 13354 484 13360 536
rect 13412 524 13418 536
rect 21910 524 21916 536
rect 13412 496 21916 524
rect 13412 484 13418 496
rect 21910 484 21916 496
rect 21968 484 21974 536
rect 3620 388 3648 484
rect 4338 416 4344 468
rect 4396 456 4402 468
rect 11256 456 11284 484
rect 4396 428 11284 456
rect 4396 416 4402 428
rect 12066 388 12072 400
rect 3620 360 12072 388
rect 12066 348 12072 360
rect 12124 348 12130 400
rect 22646 348 22652 400
rect 22704 388 22710 400
rect 24210 388 24216 400
rect 22704 360 24216 388
rect 22704 348 22710 360
rect 24210 348 24216 360
rect 24268 348 24274 400
rect 8938 280 8944 332
rect 8996 320 9002 332
rect 8996 292 12434 320
rect 8996 280 9002 292
rect 9122 212 9128 264
rect 9180 252 9186 264
rect 9674 252 9680 264
rect 9180 224 9680 252
rect 9180 212 9186 224
rect 9674 212 9680 224
rect 9732 212 9738 264
rect 12406 252 12434 292
rect 16298 252 16304 264
rect 12406 224 16304 252
rect 16298 212 16304 224
rect 16356 212 16362 264
<< via1 >>
rect 6884 6502 6936 6554
rect 6948 6502 7000 6554
rect 7012 6502 7064 6554
rect 7076 6502 7128 6554
rect 7140 6502 7192 6554
rect 12818 6502 12870 6554
rect 12882 6502 12934 6554
rect 12946 6502 12998 6554
rect 13010 6502 13062 6554
rect 13074 6502 13126 6554
rect 18752 6502 18804 6554
rect 18816 6502 18868 6554
rect 18880 6502 18932 6554
rect 18944 6502 18996 6554
rect 19008 6502 19060 6554
rect 24686 6502 24738 6554
rect 24750 6502 24802 6554
rect 24814 6502 24866 6554
rect 24878 6502 24930 6554
rect 24942 6502 24994 6554
rect 1308 6400 1360 6452
rect 2136 6400 2188 6452
rect 3792 6400 3844 6452
rect 4620 6443 4672 6452
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 5632 6332 5684 6384
rect 7288 6400 7340 6452
rect 6092 6375 6144 6384
rect 6092 6341 6101 6375
rect 6101 6341 6135 6375
rect 6135 6341 6144 6375
rect 6092 6332 6144 6341
rect 8392 6443 8444 6452
rect 8392 6409 8401 6443
rect 8401 6409 8435 6443
rect 8435 6409 8444 6443
rect 8392 6400 8444 6409
rect 9404 6443 9456 6452
rect 9404 6409 9413 6443
rect 9413 6409 9447 6443
rect 9447 6409 9456 6443
rect 9404 6400 9456 6409
rect 10600 6443 10652 6452
rect 10600 6409 10609 6443
rect 10609 6409 10643 6443
rect 10643 6409 10652 6443
rect 10600 6400 10652 6409
rect 11980 6443 12032 6452
rect 11980 6409 11989 6443
rect 11989 6409 12023 6443
rect 12023 6409 12032 6443
rect 11980 6400 12032 6409
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 9680 6264 9732 6316
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 14280 6443 14332 6452
rect 14280 6409 14289 6443
rect 14289 6409 14323 6443
rect 14323 6409 14332 6443
rect 14280 6400 14332 6409
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 17960 6443 18012 6452
rect 17960 6409 17969 6443
rect 17969 6409 18003 6443
rect 18003 6409 18012 6443
rect 17960 6400 18012 6409
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 21548 6443 21600 6452
rect 21548 6409 21557 6443
rect 21557 6409 21591 6443
rect 21591 6409 21600 6443
rect 21548 6400 21600 6409
rect 13544 6307 13596 6316
rect 13544 6273 13553 6307
rect 13553 6273 13587 6307
rect 13587 6273 13596 6307
rect 13544 6264 13596 6273
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 15660 6264 15712 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 18328 6307 18380 6316
rect 18328 6273 18337 6307
rect 18337 6273 18371 6307
rect 18371 6273 18380 6307
rect 18328 6264 18380 6273
rect 19984 6307 20036 6316
rect 19984 6273 19993 6307
rect 19993 6273 20027 6307
rect 20027 6273 20036 6307
rect 19984 6264 20036 6273
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 22560 6443 22612 6452
rect 22560 6409 22569 6443
rect 22569 6409 22603 6443
rect 22603 6409 22612 6443
rect 22560 6400 22612 6409
rect 23940 6443 23992 6452
rect 23940 6409 23949 6443
rect 23949 6409 23983 6443
rect 23983 6409 23992 6443
rect 23940 6400 23992 6409
rect 5632 6128 5684 6180
rect 21640 6196 21692 6248
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 23664 6307 23716 6316
rect 23664 6273 23673 6307
rect 23673 6273 23707 6307
rect 23707 6273 23716 6307
rect 23664 6264 23716 6273
rect 24216 6128 24268 6180
rect 3917 5958 3969 6010
rect 3981 5958 4033 6010
rect 4045 5958 4097 6010
rect 4109 5958 4161 6010
rect 4173 5958 4225 6010
rect 9851 5958 9903 6010
rect 9915 5958 9967 6010
rect 9979 5958 10031 6010
rect 10043 5958 10095 6010
rect 10107 5958 10159 6010
rect 15785 5958 15837 6010
rect 15849 5958 15901 6010
rect 15913 5958 15965 6010
rect 15977 5958 16029 6010
rect 16041 5958 16093 6010
rect 21719 5958 21771 6010
rect 21783 5958 21835 6010
rect 21847 5958 21899 6010
rect 21911 5958 21963 6010
rect 21975 5958 22027 6010
rect 6552 5856 6604 5908
rect 7564 5856 7616 5908
rect 8760 5856 8812 5908
rect 9680 5899 9732 5908
rect 9680 5865 9689 5899
rect 9689 5865 9723 5899
rect 9723 5865 9732 5899
rect 9680 5856 9732 5865
rect 11152 5856 11204 5908
rect 12348 5856 12400 5908
rect 12624 5856 12676 5908
rect 13544 5856 13596 5908
rect 14648 5856 14700 5908
rect 15108 5856 15160 5908
rect 15660 5856 15712 5908
rect 17408 5856 17460 5908
rect 18328 5856 18380 5908
rect 20536 5856 20588 5908
rect 24492 5856 24544 5908
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 8760 5695 8812 5704
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9864 5695 9916 5704
rect 9864 5661 9873 5695
rect 9873 5661 9907 5695
rect 9907 5661 9916 5695
rect 9864 5652 9916 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11980 5695 12032 5704
rect 11980 5661 11989 5695
rect 11989 5661 12023 5695
rect 12023 5661 12032 5695
rect 11980 5652 12032 5661
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 13452 5695 13504 5704
rect 13452 5661 13461 5695
rect 13461 5661 13495 5695
rect 13495 5661 13504 5695
rect 13452 5652 13504 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 19984 5788 20036 5840
rect 24032 5788 24084 5840
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 18420 5695 18472 5704
rect 18420 5661 18429 5695
rect 18429 5661 18463 5695
rect 18463 5661 18472 5695
rect 18420 5652 18472 5661
rect 19984 5695 20036 5704
rect 19984 5661 19993 5695
rect 19993 5661 20027 5695
rect 20027 5661 20036 5695
rect 19984 5652 20036 5661
rect 23848 5627 23900 5636
rect 23848 5593 23857 5627
rect 23857 5593 23891 5627
rect 23891 5593 23900 5627
rect 23848 5584 23900 5593
rect 6884 5414 6936 5466
rect 6948 5414 7000 5466
rect 7012 5414 7064 5466
rect 7076 5414 7128 5466
rect 7140 5414 7192 5466
rect 12818 5414 12870 5466
rect 12882 5414 12934 5466
rect 12946 5414 12998 5466
rect 13010 5414 13062 5466
rect 13074 5414 13126 5466
rect 18752 5414 18804 5466
rect 18816 5414 18868 5466
rect 18880 5414 18932 5466
rect 18944 5414 18996 5466
rect 19008 5414 19060 5466
rect 24686 5414 24738 5466
rect 24750 5414 24802 5466
rect 24814 5414 24866 5466
rect 24878 5414 24930 5466
rect 24942 5414 24994 5466
rect 6276 5312 6328 5364
rect 7564 5355 7616 5364
rect 7564 5321 7573 5355
rect 7573 5321 7607 5355
rect 7607 5321 7616 5355
rect 7564 5312 7616 5321
rect 8760 5355 8812 5364
rect 8760 5321 8769 5355
rect 8769 5321 8803 5355
rect 8803 5321 8812 5355
rect 8760 5312 8812 5321
rect 9864 5355 9916 5364
rect 9864 5321 9873 5355
rect 9873 5321 9907 5355
rect 9907 5321 9916 5355
rect 9864 5312 9916 5321
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 12440 5355 12492 5364
rect 12440 5321 12449 5355
rect 12449 5321 12483 5355
rect 12483 5321 12492 5355
rect 12440 5312 12492 5321
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 15936 5355 15988 5364
rect 15936 5321 15945 5355
rect 15945 5321 15979 5355
rect 15979 5321 15988 5355
rect 15936 5312 15988 5321
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 18420 5355 18472 5364
rect 18420 5321 18429 5355
rect 18429 5321 18463 5355
rect 18463 5321 18472 5355
rect 18420 5312 18472 5321
rect 19984 5355 20036 5364
rect 19984 5321 19993 5355
rect 19993 5321 20027 5355
rect 20027 5321 20036 5355
rect 19984 5312 20036 5321
rect 23848 5312 23900 5364
rect 13176 5244 13228 5296
rect 8208 4972 8260 5024
rect 10968 5176 11020 5228
rect 11244 5219 11296 5228
rect 11244 5185 11253 5219
rect 11253 5185 11287 5219
rect 11287 5185 11296 5219
rect 11244 5176 11296 5185
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 14464 5176 14516 5228
rect 24400 5244 24452 5296
rect 14188 5108 14240 5160
rect 17132 5108 17184 5160
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 21180 5176 21232 5228
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 23756 5108 23808 5160
rect 22560 5040 22612 5092
rect 17224 4972 17276 5024
rect 3917 4870 3969 4922
rect 3981 4870 4033 4922
rect 4045 4870 4097 4922
rect 4109 4870 4161 4922
rect 4173 4870 4225 4922
rect 9851 4870 9903 4922
rect 9915 4870 9967 4922
rect 9979 4870 10031 4922
rect 10043 4870 10095 4922
rect 10107 4870 10159 4922
rect 15785 4870 15837 4922
rect 15849 4870 15901 4922
rect 15913 4870 15965 4922
rect 15977 4870 16029 4922
rect 16041 4870 16093 4922
rect 21719 4870 21771 4922
rect 21783 4870 21835 4922
rect 21847 4870 21899 4922
rect 21911 4870 21963 4922
rect 21975 4870 22027 4922
rect 24308 4768 24360 4820
rect 22928 4564 22980 4616
rect 6884 4326 6936 4378
rect 6948 4326 7000 4378
rect 7012 4326 7064 4378
rect 7076 4326 7128 4378
rect 7140 4326 7192 4378
rect 12818 4326 12870 4378
rect 12882 4326 12934 4378
rect 12946 4326 12998 4378
rect 13010 4326 13062 4378
rect 13074 4326 13126 4378
rect 18752 4326 18804 4378
rect 18816 4326 18868 4378
rect 18880 4326 18932 4378
rect 18944 4326 18996 4378
rect 19008 4326 19060 4378
rect 24686 4326 24738 4378
rect 24750 4326 24802 4378
rect 24814 4326 24866 4378
rect 24878 4326 24930 4378
rect 24942 4326 24994 4378
rect 7656 4224 7708 4276
rect 17132 4156 17184 4208
rect 17868 4156 17920 4208
rect 17960 4156 18012 4208
rect 3917 3782 3969 3834
rect 3981 3782 4033 3834
rect 4045 3782 4097 3834
rect 4109 3782 4161 3834
rect 4173 3782 4225 3834
rect 9851 3782 9903 3834
rect 9915 3782 9967 3834
rect 9979 3782 10031 3834
rect 10043 3782 10095 3834
rect 10107 3782 10159 3834
rect 15785 3782 15837 3834
rect 15849 3782 15901 3834
rect 15913 3782 15965 3834
rect 15977 3782 16029 3834
rect 16041 3782 16093 3834
rect 21719 3782 21771 3834
rect 21783 3782 21835 3834
rect 21847 3782 21899 3834
rect 21911 3782 21963 3834
rect 21975 3782 22027 3834
rect 23664 3680 23716 3732
rect 24124 3519 24176 3528
rect 24124 3485 24133 3519
rect 24133 3485 24167 3519
rect 24167 3485 24176 3519
rect 24124 3476 24176 3485
rect 13636 3408 13688 3460
rect 22192 3408 22244 3460
rect 6884 3238 6936 3290
rect 6948 3238 7000 3290
rect 7012 3238 7064 3290
rect 7076 3238 7128 3290
rect 7140 3238 7192 3290
rect 12818 3238 12870 3290
rect 12882 3238 12934 3290
rect 12946 3238 12998 3290
rect 13010 3238 13062 3290
rect 13074 3238 13126 3290
rect 18752 3238 18804 3290
rect 18816 3238 18868 3290
rect 18880 3238 18932 3290
rect 18944 3238 18996 3290
rect 19008 3238 19060 3290
rect 24686 3238 24738 3290
rect 24750 3238 24802 3290
rect 24814 3238 24866 3290
rect 24878 3238 24930 3290
rect 24942 3238 24994 3290
rect 24124 3179 24176 3188
rect 24124 3145 24133 3179
rect 24133 3145 24167 3179
rect 24167 3145 24176 3179
rect 24124 3136 24176 3145
rect 10968 3068 11020 3120
rect 16672 3068 16724 3120
rect 1400 3000 1452 3052
rect 10416 3000 10468 3052
rect 11244 3000 11296 3052
rect 15200 3000 15252 3052
rect 25044 3068 25096 3120
rect 5908 2932 5960 2984
rect 9588 2932 9640 2984
rect 10784 2932 10836 2984
rect 2688 2864 2740 2916
rect 7472 2864 7524 2916
rect 8024 2864 8076 2916
rect 15016 2864 15068 2916
rect 17224 2932 17276 2984
rect 22284 2932 22336 2984
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 24492 2932 24544 2984
rect 24584 2864 24636 2916
rect 1952 2796 2004 2848
rect 6736 2796 6788 2848
rect 9496 2796 9548 2848
rect 12440 2796 12492 2848
rect 16764 2796 16816 2848
rect 22836 2796 22888 2848
rect 23664 2796 23716 2848
rect 24032 2796 24084 2848
rect 3917 2694 3969 2746
rect 3981 2694 4033 2746
rect 4045 2694 4097 2746
rect 4109 2694 4161 2746
rect 4173 2694 4225 2746
rect 9851 2694 9903 2746
rect 9915 2694 9967 2746
rect 9979 2694 10031 2746
rect 10043 2694 10095 2746
rect 10107 2694 10159 2746
rect 15785 2694 15837 2746
rect 15849 2694 15901 2746
rect 15913 2694 15965 2746
rect 15977 2694 16029 2746
rect 16041 2694 16093 2746
rect 21719 2694 21771 2746
rect 21783 2694 21835 2746
rect 21847 2694 21899 2746
rect 21911 2694 21963 2746
rect 21975 2694 22027 2746
rect 3424 2592 3476 2644
rect 7196 2592 7248 2644
rect 10692 2592 10744 2644
rect 11060 2592 11112 2644
rect 1584 2567 1636 2576
rect 1584 2533 1593 2567
rect 1593 2533 1627 2567
rect 1627 2533 1636 2567
rect 1584 2524 1636 2533
rect 1952 2567 2004 2576
rect 1952 2533 1961 2567
rect 1961 2533 1995 2567
rect 1995 2533 2004 2567
rect 1952 2524 2004 2533
rect 7840 2524 7892 2576
rect 10784 2524 10836 2576
rect 11980 2524 12032 2576
rect 480 2456 532 2508
rect 1308 2388 1360 2440
rect 2596 2456 2648 2508
rect 204 2320 256 2372
rect 1952 2320 2004 2372
rect 4620 2388 4672 2440
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 7196 2388 7248 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7748 2388 7800 2440
rect 10876 2456 10928 2508
rect 10968 2456 11020 2508
rect 9312 2388 9364 2440
rect 9680 2388 9732 2440
rect 9220 2320 9272 2372
rect 10600 2388 10652 2440
rect 11796 2388 11848 2440
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 13452 2456 13504 2508
rect 15292 2427 15344 2440
rect 15292 2393 15301 2427
rect 15301 2393 15335 2427
rect 15335 2393 15344 2427
rect 15292 2388 15344 2393
rect 17408 2592 17460 2644
rect 17868 2592 17920 2644
rect 22928 2635 22980 2644
rect 22928 2601 22937 2635
rect 22937 2601 22971 2635
rect 22971 2601 22980 2635
rect 22928 2592 22980 2601
rect 16028 2456 16080 2508
rect 18604 2524 18656 2576
rect 16488 2431 16540 2440
rect 16488 2397 16497 2431
rect 16497 2397 16531 2431
rect 16531 2397 16540 2431
rect 16488 2388 16540 2397
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 17960 2456 18012 2508
rect 23756 2635 23808 2644
rect 23756 2601 23765 2635
rect 23765 2601 23799 2635
rect 23799 2601 23808 2635
rect 23756 2592 23808 2601
rect 24308 2592 24360 2644
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 18696 2431 18748 2440
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 2872 2252 2924 2304
rect 4252 2252 4304 2304
rect 4344 2252 4396 2304
rect 6276 2295 6328 2304
rect 6276 2261 6285 2295
rect 6285 2261 6319 2295
rect 6319 2261 6328 2295
rect 6276 2252 6328 2261
rect 8116 2252 8168 2304
rect 9128 2252 9180 2304
rect 9404 2295 9456 2304
rect 9404 2261 9413 2295
rect 9413 2261 9447 2295
rect 9447 2261 9456 2295
rect 9404 2252 9456 2261
rect 9772 2252 9824 2304
rect 10876 2252 10928 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 12348 2295 12400 2304
rect 12348 2261 12357 2295
rect 12357 2261 12391 2295
rect 12391 2261 12400 2295
rect 12348 2252 12400 2261
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 14004 2252 14056 2304
rect 14096 2252 14148 2304
rect 15108 2252 15160 2304
rect 15384 2295 15436 2304
rect 15384 2261 15393 2295
rect 15393 2261 15427 2295
rect 15427 2261 15436 2295
rect 15384 2252 15436 2261
rect 15568 2252 15620 2304
rect 16304 2252 16356 2304
rect 16856 2295 16908 2304
rect 16856 2261 16865 2295
rect 16865 2261 16899 2295
rect 16899 2261 16908 2295
rect 16856 2252 16908 2261
rect 16948 2252 17000 2304
rect 18328 2320 18380 2372
rect 17776 2252 17828 2304
rect 18144 2252 18196 2304
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 18604 2252 18656 2304
rect 19156 2252 19208 2304
rect 19248 2295 19300 2304
rect 19248 2261 19257 2295
rect 19257 2261 19291 2295
rect 19291 2261 19300 2295
rect 19248 2252 19300 2261
rect 19708 2431 19760 2440
rect 19708 2397 19717 2431
rect 19717 2397 19751 2431
rect 19751 2397 19760 2431
rect 19708 2388 19760 2397
rect 20168 2388 20220 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 19984 2252 20036 2304
rect 20444 2320 20496 2372
rect 22376 2431 22428 2440
rect 22376 2397 22385 2431
rect 22385 2397 22419 2431
rect 22419 2397 22428 2431
rect 22376 2388 22428 2397
rect 22836 2431 22888 2440
rect 22836 2397 22845 2431
rect 22845 2397 22879 2431
rect 22879 2397 22888 2431
rect 22836 2388 22888 2397
rect 23296 2388 23348 2440
rect 23388 2431 23440 2440
rect 23388 2397 23397 2431
rect 23397 2397 23431 2431
rect 23431 2397 23440 2431
rect 23388 2388 23440 2397
rect 23940 2431 23992 2440
rect 23940 2397 23949 2431
rect 23949 2397 23983 2431
rect 23983 2397 23992 2431
rect 23940 2388 23992 2397
rect 24032 2388 24084 2440
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 20628 2295 20680 2304
rect 20628 2261 20637 2295
rect 20637 2261 20671 2295
rect 20671 2261 20680 2295
rect 20628 2252 20680 2261
rect 22744 2252 22796 2304
rect 24032 2295 24084 2304
rect 24032 2261 24041 2295
rect 24041 2261 24075 2295
rect 24075 2261 24084 2295
rect 24032 2252 24084 2261
rect 24216 2252 24268 2304
rect 6884 2150 6936 2202
rect 6948 2150 7000 2202
rect 7012 2150 7064 2202
rect 7076 2150 7128 2202
rect 7140 2150 7192 2202
rect 12818 2150 12870 2202
rect 12882 2150 12934 2202
rect 12946 2150 12998 2202
rect 13010 2150 13062 2202
rect 13074 2150 13126 2202
rect 18752 2150 18804 2202
rect 18816 2150 18868 2202
rect 18880 2150 18932 2202
rect 18944 2150 18996 2202
rect 19008 2150 19060 2202
rect 24686 2150 24738 2202
rect 24750 2150 24802 2202
rect 24814 2150 24866 2202
rect 24878 2150 24930 2202
rect 24942 2150 24994 2202
rect 2688 2091 2740 2100
rect 2688 2057 2697 2091
rect 2697 2057 2731 2091
rect 2731 2057 2740 2091
rect 2688 2048 2740 2057
rect 1768 1955 1820 1964
rect 1768 1921 1777 1955
rect 1777 1921 1811 1955
rect 1811 1921 1820 1955
rect 1768 1912 1820 1921
rect 2136 1955 2188 1964
rect 2136 1921 2145 1955
rect 2145 1921 2179 1955
rect 2179 1921 2188 1955
rect 2136 1912 2188 1921
rect 756 1844 808 1896
rect 1032 1776 1084 1828
rect 3148 1955 3200 1964
rect 3148 1921 3157 1955
rect 3157 1921 3191 1955
rect 3191 1921 3200 1955
rect 3148 1912 3200 1921
rect 3608 1912 3660 1964
rect 3792 1912 3844 1964
rect 3332 1776 3384 1828
rect 3608 1776 3660 1828
rect 1492 1751 1544 1760
rect 1492 1717 1501 1751
rect 1501 1717 1535 1751
rect 1535 1717 1544 1751
rect 1492 1708 1544 1717
rect 2228 1708 2280 1760
rect 2320 1751 2372 1760
rect 2320 1717 2329 1751
rect 2329 1717 2363 1751
rect 2363 1717 2372 1751
rect 2320 1708 2372 1717
rect 2964 1751 3016 1760
rect 2964 1717 2973 1751
rect 2973 1717 3007 1751
rect 3007 1717 3016 1751
rect 2964 1708 3016 1717
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 4712 1912 4764 1964
rect 4988 1912 5040 1964
rect 5264 1912 5316 1964
rect 4436 1844 4488 1896
rect 6552 1912 6604 1964
rect 6644 1955 6696 1964
rect 6644 1921 6653 1955
rect 6653 1921 6687 1955
rect 6687 1921 6696 1955
rect 6644 1912 6696 1921
rect 7472 2048 7524 2100
rect 7748 2048 7800 2100
rect 7840 2091 7892 2100
rect 7840 2057 7849 2091
rect 7849 2057 7883 2091
rect 7883 2057 7892 2091
rect 7840 2048 7892 2057
rect 8024 2048 8076 2100
rect 7380 1912 7432 1964
rect 7472 1955 7524 1964
rect 7472 1921 7481 1955
rect 7481 1921 7515 1955
rect 7515 1921 7524 1955
rect 7472 1912 7524 1921
rect 7748 1955 7800 1964
rect 7748 1921 7757 1955
rect 7757 1921 7791 1955
rect 7791 1921 7800 1955
rect 7748 1912 7800 1921
rect 8024 1955 8076 1964
rect 8024 1921 8033 1955
rect 8033 1921 8067 1955
rect 8067 1921 8076 1955
rect 8024 1912 8076 1921
rect 8300 1955 8352 1964
rect 8300 1921 8309 1955
rect 8309 1921 8343 1955
rect 8343 1921 8352 1955
rect 8300 1912 8352 1921
rect 6276 1844 6328 1896
rect 7564 1844 7616 1896
rect 7840 1844 7892 1896
rect 8760 1980 8812 2032
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 9128 1955 9180 1964
rect 9128 1921 9137 1955
rect 9137 1921 9171 1955
rect 9171 1921 9180 1955
rect 9128 1912 9180 1921
rect 9404 1955 9456 1964
rect 9404 1921 9405 1955
rect 9405 1921 9439 1955
rect 9439 1921 9456 1955
rect 9404 1912 9456 1921
rect 10416 2023 10468 2032
rect 10416 1989 10425 2023
rect 10425 1989 10459 2023
rect 10459 1989 10468 2023
rect 10416 1980 10468 1989
rect 12624 2048 12676 2100
rect 11244 1980 11296 2032
rect 10048 1912 10100 1964
rect 10324 1912 10376 1964
rect 11336 1912 11388 1964
rect 12348 1912 12400 1964
rect 13544 1912 13596 1964
rect 14004 2048 14056 2100
rect 15292 2048 15344 2100
rect 15384 2048 15436 2100
rect 17592 2048 17644 2100
rect 17868 2048 17920 2100
rect 18236 2048 18288 2100
rect 18328 2048 18380 2100
rect 14004 1912 14056 1964
rect 14280 1912 14332 1964
rect 14372 1955 14424 1964
rect 14372 1921 14381 1955
rect 14381 1921 14415 1955
rect 14415 1921 14424 1955
rect 14372 1912 14424 1921
rect 8116 1776 8168 1828
rect 12072 1844 12124 1896
rect 9036 1776 9088 1828
rect 4068 1751 4120 1760
rect 4068 1717 4077 1751
rect 4077 1717 4111 1751
rect 4111 1717 4120 1751
rect 4068 1708 4120 1717
rect 4252 1708 4304 1760
rect 5172 1751 5224 1760
rect 5172 1717 5181 1751
rect 5181 1717 5215 1751
rect 5215 1717 5224 1751
rect 5172 1708 5224 1717
rect 5540 1708 5592 1760
rect 6000 1751 6052 1760
rect 6000 1717 6009 1751
rect 6009 1717 6043 1751
rect 6043 1717 6052 1751
rect 6000 1708 6052 1717
rect 6460 1751 6512 1760
rect 6460 1717 6469 1751
rect 6469 1717 6503 1751
rect 6503 1717 6512 1751
rect 6460 1708 6512 1717
rect 6736 1751 6788 1760
rect 6736 1717 6745 1751
rect 6745 1717 6779 1751
rect 6779 1717 6788 1751
rect 6736 1708 6788 1717
rect 7104 1708 7156 1760
rect 8208 1708 8260 1760
rect 8668 1751 8720 1760
rect 8668 1717 8677 1751
rect 8677 1717 8711 1751
rect 8711 1717 8720 1751
rect 8668 1708 8720 1717
rect 9496 1819 9548 1828
rect 9496 1785 9505 1819
rect 9505 1785 9539 1819
rect 9539 1785 9548 1819
rect 9496 1776 9548 1785
rect 9680 1776 9732 1828
rect 13452 1776 13504 1828
rect 15108 1912 15160 1964
rect 16028 1980 16080 2032
rect 16120 1912 16172 1964
rect 17776 1980 17828 2032
rect 18420 1912 18472 1964
rect 19156 2048 19208 2100
rect 19248 2048 19300 2100
rect 20352 2048 20404 2100
rect 21088 2048 21140 2100
rect 21180 2048 21232 2100
rect 21640 2048 21692 2100
rect 22284 2091 22336 2100
rect 22284 2057 22293 2091
rect 22293 2057 22327 2091
rect 22327 2057 22336 2091
rect 22284 2048 22336 2057
rect 23112 2048 23164 2100
rect 24032 2048 24084 2100
rect 24400 2091 24452 2100
rect 24400 2057 24409 2091
rect 24409 2057 24443 2091
rect 24443 2057 24452 2091
rect 24400 2048 24452 2057
rect 19892 1980 19944 2032
rect 20628 1980 20680 2032
rect 23388 1980 23440 2032
rect 21088 1955 21140 1964
rect 21088 1921 21097 1955
rect 21097 1921 21131 1955
rect 21131 1921 21140 1955
rect 21088 1912 21140 1921
rect 21272 1912 21324 1964
rect 22008 1955 22060 1964
rect 22008 1921 22017 1955
rect 22017 1921 22051 1955
rect 22051 1921 22060 1955
rect 22008 1912 22060 1921
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 10968 1708 11020 1760
rect 11704 1751 11756 1760
rect 11704 1717 11713 1751
rect 11713 1717 11747 1751
rect 11747 1717 11756 1751
rect 11704 1708 11756 1717
rect 11796 1708 11848 1760
rect 12808 1708 12860 1760
rect 12900 1751 12952 1760
rect 12900 1717 12909 1751
rect 12909 1717 12943 1751
rect 12943 1717 12952 1751
rect 12900 1708 12952 1717
rect 13820 1708 13872 1760
rect 15384 1776 15436 1828
rect 17776 1776 17828 1828
rect 14280 1708 14332 1760
rect 14740 1708 14792 1760
rect 15476 1751 15528 1760
rect 15476 1717 15485 1751
rect 15485 1717 15519 1751
rect 15519 1717 15528 1751
rect 15476 1708 15528 1717
rect 15660 1708 15712 1760
rect 16580 1708 16632 1760
rect 16764 1708 16816 1760
rect 17960 1708 18012 1760
rect 18236 1708 18288 1760
rect 19432 1776 19484 1828
rect 19340 1708 19392 1760
rect 21180 1776 21232 1828
rect 20904 1751 20956 1760
rect 20904 1717 20913 1751
rect 20913 1717 20947 1751
rect 20947 1717 20956 1751
rect 20904 1708 20956 1717
rect 21732 1844 21784 1896
rect 22468 1912 22520 1964
rect 22744 1912 22796 1964
rect 23020 1955 23072 1964
rect 23020 1921 23029 1955
rect 23029 1921 23063 1955
rect 23063 1921 23072 1955
rect 23020 1912 23072 1921
rect 22192 1844 22244 1896
rect 22376 1844 22428 1896
rect 23112 1844 23164 1896
rect 24308 1844 24360 1896
rect 23480 1776 23532 1828
rect 23756 1776 23808 1828
rect 24124 1708 24176 1760
rect 3917 1606 3969 1658
rect 3981 1606 4033 1658
rect 4045 1606 4097 1658
rect 4109 1606 4161 1658
rect 4173 1606 4225 1658
rect 9851 1606 9903 1658
rect 9915 1606 9967 1658
rect 9979 1606 10031 1658
rect 10043 1606 10095 1658
rect 10107 1606 10159 1658
rect 15785 1606 15837 1658
rect 15849 1606 15901 1658
rect 15913 1606 15965 1658
rect 15977 1606 16029 1658
rect 16041 1606 16093 1658
rect 21719 1606 21771 1658
rect 21783 1606 21835 1658
rect 21847 1606 21899 1658
rect 21911 1606 21963 1658
rect 21975 1606 22027 1658
rect 2596 1547 2648 1556
rect 2596 1513 2605 1547
rect 2605 1513 2639 1547
rect 2639 1513 2648 1547
rect 2596 1504 2648 1513
rect 2872 1547 2924 1556
rect 2872 1513 2881 1547
rect 2881 1513 2915 1547
rect 2915 1513 2924 1547
rect 2872 1504 2924 1513
rect 1400 1300 1452 1352
rect 1492 1300 1544 1352
rect 3240 1368 3292 1420
rect 2780 1343 2832 1352
rect 2780 1309 2789 1343
rect 2789 1309 2823 1343
rect 2823 1309 2832 1343
rect 2780 1300 2832 1309
rect 3056 1343 3108 1352
rect 3056 1309 3065 1343
rect 3065 1309 3099 1343
rect 3099 1309 3108 1343
rect 3056 1300 3108 1309
rect 4344 1504 4396 1556
rect 5908 1504 5960 1556
rect 6000 1504 6052 1556
rect 6920 1504 6972 1556
rect 7104 1504 7156 1556
rect 3516 1300 3568 1352
rect 3884 1300 3936 1352
rect 1676 1164 1728 1216
rect 2044 1207 2096 1216
rect 2044 1173 2053 1207
rect 2053 1173 2087 1207
rect 2087 1173 2096 1207
rect 2044 1164 2096 1173
rect 2688 1232 2740 1284
rect 8484 1436 8536 1488
rect 8576 1479 8628 1488
rect 8576 1445 8585 1479
rect 8585 1445 8619 1479
rect 8619 1445 8628 1479
rect 8576 1436 8628 1445
rect 8944 1436 8996 1488
rect 5172 1300 5224 1352
rect 5540 1300 5592 1352
rect 6460 1300 6512 1352
rect 6736 1300 6788 1352
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 6920 1300 6972 1352
rect 7012 1300 7064 1352
rect 7840 1368 7892 1420
rect 8392 1368 8444 1420
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8484 1343 8536 1352
rect 8484 1309 8493 1343
rect 8493 1309 8527 1343
rect 8527 1309 8536 1343
rect 8484 1300 8536 1309
rect 9220 1300 9272 1352
rect 9496 1343 9548 1352
rect 9496 1309 9505 1343
rect 9505 1309 9539 1343
rect 9539 1309 9548 1343
rect 9496 1300 9548 1309
rect 2228 1164 2280 1216
rect 2320 1207 2372 1216
rect 2320 1173 2329 1207
rect 2329 1173 2363 1207
rect 2363 1173 2372 1207
rect 2320 1164 2372 1173
rect 3332 1164 3384 1216
rect 3516 1164 3568 1216
rect 3976 1164 4028 1216
rect 4344 1207 4396 1216
rect 4344 1173 4353 1207
rect 4353 1173 4387 1207
rect 4387 1173 4396 1207
rect 4344 1164 4396 1173
rect 4804 1207 4856 1216
rect 4804 1173 4813 1207
rect 4813 1173 4847 1207
rect 4847 1173 4856 1207
rect 4804 1164 4856 1173
rect 5172 1207 5224 1216
rect 5172 1173 5181 1207
rect 5181 1173 5215 1207
rect 5215 1173 5224 1207
rect 5172 1164 5224 1173
rect 5448 1207 5500 1216
rect 5448 1173 5457 1207
rect 5457 1173 5491 1207
rect 5491 1173 5500 1207
rect 5448 1164 5500 1173
rect 5540 1164 5592 1216
rect 6368 1207 6420 1216
rect 6368 1173 6377 1207
rect 6377 1173 6411 1207
rect 6411 1173 6420 1207
rect 6368 1164 6420 1173
rect 7840 1232 7892 1284
rect 7196 1164 7248 1216
rect 7656 1164 7708 1216
rect 7932 1164 7984 1216
rect 9128 1232 9180 1284
rect 9772 1300 9824 1352
rect 11060 1411 11112 1420
rect 11060 1377 11069 1411
rect 11069 1377 11103 1411
rect 11103 1377 11112 1411
rect 11060 1368 11112 1377
rect 9864 1232 9916 1284
rect 8208 1164 8260 1216
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 9680 1164 9732 1216
rect 10048 1164 10100 1216
rect 10692 1232 10744 1284
rect 10784 1275 10836 1284
rect 10784 1241 10793 1275
rect 10793 1241 10827 1275
rect 10827 1241 10836 1275
rect 10784 1232 10836 1241
rect 11152 1164 11204 1216
rect 11980 1436 12032 1488
rect 12532 1436 12584 1488
rect 13820 1504 13872 1556
rect 14924 1504 14976 1556
rect 11520 1368 11572 1420
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 11612 1164 11664 1216
rect 12440 1300 12492 1352
rect 12808 1368 12860 1420
rect 15292 1436 15344 1488
rect 16488 1504 16540 1556
rect 16028 1436 16080 1488
rect 13912 1300 13964 1352
rect 15384 1368 15436 1420
rect 16212 1368 16264 1420
rect 17592 1504 17644 1556
rect 19800 1504 19852 1556
rect 21180 1504 21232 1556
rect 22100 1504 22152 1556
rect 18696 1436 18748 1488
rect 17592 1368 17644 1420
rect 18144 1368 18196 1420
rect 18604 1368 18656 1420
rect 21548 1436 21600 1488
rect 21456 1368 21508 1420
rect 21824 1479 21876 1488
rect 21824 1445 21833 1479
rect 21833 1445 21867 1479
rect 21867 1445 21876 1479
rect 21824 1436 21876 1445
rect 22008 1436 22060 1488
rect 14648 1343 14700 1352
rect 14648 1309 14657 1343
rect 14657 1309 14691 1343
rect 14691 1309 14700 1343
rect 14648 1300 14700 1309
rect 15476 1300 15528 1352
rect 12072 1164 12124 1216
rect 12348 1207 12400 1216
rect 12348 1173 12357 1207
rect 12357 1173 12391 1207
rect 12391 1173 12400 1207
rect 12348 1164 12400 1173
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13452 1207 13504 1216
rect 13452 1173 13461 1207
rect 13461 1173 13495 1207
rect 13495 1173 13504 1207
rect 13452 1164 13504 1173
rect 14004 1164 14056 1216
rect 15016 1164 15068 1216
rect 16580 1300 16632 1352
rect 16856 1300 16908 1352
rect 16396 1232 16448 1284
rect 17408 1232 17460 1284
rect 18512 1232 18564 1284
rect 18696 1232 18748 1284
rect 19984 1300 20036 1352
rect 21732 1300 21784 1352
rect 16488 1164 16540 1216
rect 19616 1232 19668 1284
rect 19064 1164 19116 1216
rect 20536 1164 20588 1216
rect 21916 1164 21968 1216
rect 22560 1300 22612 1352
rect 22744 1300 22796 1352
rect 22928 1343 22980 1352
rect 22928 1309 22937 1343
rect 22937 1309 22971 1343
rect 22971 1309 22980 1343
rect 22928 1300 22980 1309
rect 23480 1436 23532 1488
rect 23756 1436 23808 1488
rect 25320 1436 25372 1488
rect 23848 1300 23900 1352
rect 24032 1343 24084 1352
rect 24032 1309 24041 1343
rect 24041 1309 24075 1343
rect 24075 1309 24084 1343
rect 24032 1300 24084 1309
rect 22284 1207 22336 1216
rect 22284 1173 22293 1207
rect 22293 1173 22327 1207
rect 22327 1173 22336 1207
rect 22284 1164 22336 1173
rect 23112 1207 23164 1216
rect 23112 1173 23121 1207
rect 23121 1173 23155 1207
rect 23155 1173 23164 1207
rect 23112 1164 23164 1173
rect 23664 1207 23716 1216
rect 23664 1173 23673 1207
rect 23673 1173 23707 1207
rect 23707 1173 23716 1207
rect 23664 1164 23716 1173
rect 23756 1164 23808 1216
rect 24308 1164 24360 1216
rect 6884 1062 6936 1114
rect 6948 1062 7000 1114
rect 7012 1062 7064 1114
rect 7076 1062 7128 1114
rect 7140 1062 7192 1114
rect 12818 1062 12870 1114
rect 12882 1062 12934 1114
rect 12946 1062 12998 1114
rect 13010 1062 13062 1114
rect 13074 1062 13126 1114
rect 18752 1062 18804 1114
rect 18816 1062 18868 1114
rect 18880 1062 18932 1114
rect 18944 1062 18996 1114
rect 19008 1062 19060 1114
rect 24686 1062 24738 1114
rect 24750 1062 24802 1114
rect 24814 1062 24866 1114
rect 24878 1062 24930 1114
rect 24942 1062 24994 1114
rect 2044 960 2096 1012
rect 2320 892 2372 944
rect 5448 960 5500 1012
rect 10784 960 10836 1012
rect 10876 960 10928 1012
rect 16396 960 16448 1012
rect 16948 960 17000 1012
rect 19616 960 19668 1012
rect 21916 960 21968 1012
rect 23112 960 23164 1012
rect 23664 960 23716 1012
rect 24308 960 24360 1012
rect 8576 892 8628 944
rect 9680 892 9732 944
rect 6368 824 6420 876
rect 11612 824 11664 876
rect 3424 756 3476 808
rect 6736 756 6788 808
rect 7564 756 7616 808
rect 8024 756 8076 808
rect 14648 892 14700 944
rect 16672 892 16724 944
rect 14188 824 14240 876
rect 3976 688 4028 740
rect 9220 620 9272 672
rect 20904 756 20956 808
rect 21732 756 21784 808
rect 12440 688 12492 740
rect 12900 688 12952 740
rect 14464 688 14516 740
rect 22284 756 22336 808
rect 22928 756 22980 808
rect 23296 756 23348 808
rect 25596 756 25648 808
rect 13544 620 13596 672
rect 15200 620 15252 672
rect 6920 552 6972 604
rect 16120 552 16172 604
rect 20352 620 20404 672
rect 21272 620 21324 672
rect 21456 620 21508 672
rect 23572 688 23624 740
rect 2780 484 2832 536
rect 3516 484 3568 536
rect 3608 484 3660 536
rect 5172 484 5224 536
rect 9864 484 9916 536
rect 11244 484 11296 536
rect 13360 484 13412 536
rect 21916 484 21968 536
rect 4344 416 4396 468
rect 12072 348 12124 400
rect 22652 348 22704 400
rect 24216 348 24268 400
rect 8944 280 8996 332
rect 9128 212 9180 264
rect 9680 212 9732 264
rect 16304 212 16356 264
<< metal2 >>
rect 938 7970 994 8000
rect 938 7942 1348 7970
rect 938 7840 994 7942
rect 1320 6458 1348 7942
rect 2134 7840 2190 8000
rect 3330 7970 3386 8000
rect 4526 7970 4582 8000
rect 5722 7970 5778 8000
rect 6918 7970 6974 8000
rect 8114 7970 8170 8000
rect 9310 7970 9366 8000
rect 10506 7970 10562 8000
rect 11702 7970 11758 8000
rect 12898 7970 12954 8000
rect 14094 7970 14150 8000
rect 15290 7970 15346 8000
rect 16486 7970 16542 8000
rect 17682 7970 17738 8000
rect 18878 7970 18934 8000
rect 20074 7970 20130 8000
rect 21270 7970 21326 8000
rect 22466 7970 22522 8000
rect 3330 7942 3832 7970
rect 3330 7840 3386 7942
rect 2148 6458 2176 7840
rect 3804 6458 3832 7942
rect 4526 7942 4660 7970
rect 4526 7840 4582 7942
rect 4632 6458 4660 7942
rect 5722 7942 6132 7970
rect 5722 7840 5778 7942
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 6104 6390 6132 7942
rect 6918 7942 7328 7970
rect 6918 7840 6974 7942
rect 6884 6556 7192 6565
rect 6884 6554 6890 6556
rect 6946 6554 6970 6556
rect 7026 6554 7050 6556
rect 7106 6554 7130 6556
rect 7186 6554 7192 6556
rect 6946 6502 6948 6554
rect 7128 6502 7130 6554
rect 6884 6500 6890 6502
rect 6946 6500 6970 6502
rect 7026 6500 7050 6502
rect 7106 6500 7130 6502
rect 7186 6500 7192 6502
rect 6884 6491 7192 6500
rect 7300 6458 7328 7942
rect 8114 7942 8432 7970
rect 8114 7840 8170 7942
rect 8404 6458 8432 7942
rect 9310 7942 9444 7970
rect 9310 7840 9366 7942
rect 9416 6458 9444 7942
rect 10506 7942 10640 7970
rect 10506 7840 10562 7942
rect 10612 6458 10640 7942
rect 11702 7942 12020 7970
rect 11702 7840 11758 7942
rect 11992 6458 12020 7942
rect 12898 7942 13216 7970
rect 12898 7840 12954 7942
rect 12818 6556 13126 6565
rect 12818 6554 12824 6556
rect 12880 6554 12904 6556
rect 12960 6554 12984 6556
rect 13040 6554 13064 6556
rect 13120 6554 13126 6556
rect 12880 6502 12882 6554
rect 13062 6502 13064 6554
rect 12818 6500 12824 6502
rect 12880 6500 12904 6502
rect 12960 6500 12984 6502
rect 13040 6500 13064 6502
rect 13120 6500 13126 6502
rect 12818 6491 13126 6500
rect 13188 6458 13216 7942
rect 14094 7942 14320 7970
rect 14094 7840 14150 7942
rect 14292 6458 14320 7942
rect 15290 7942 15424 7970
rect 15290 7840 15346 7942
rect 15396 6458 15424 7942
rect 16486 7942 16896 7970
rect 16486 7840 16542 7942
rect 16868 6458 16896 7942
rect 17682 7942 18000 7970
rect 17682 7840 17738 7942
rect 17972 6458 18000 7942
rect 18878 7942 19472 7970
rect 18878 7840 18934 7942
rect 18752 6556 19060 6565
rect 18752 6554 18758 6556
rect 18814 6554 18838 6556
rect 18894 6554 18918 6556
rect 18974 6554 18998 6556
rect 19054 6554 19060 6556
rect 18814 6502 18816 6554
rect 18996 6502 18998 6554
rect 18752 6500 18758 6502
rect 18814 6500 18838 6502
rect 18894 6500 18918 6502
rect 18974 6500 18998 6502
rect 19054 6500 19060 6502
rect 18752 6491 19060 6500
rect 19444 6458 19472 7942
rect 20074 7942 20392 7970
rect 20074 7840 20130 7942
rect 20364 6458 20392 7942
rect 21270 7942 21588 7970
rect 21270 7840 21326 7942
rect 21560 6458 21588 7942
rect 22466 7942 22600 7970
rect 22466 7840 22522 7942
rect 22572 6458 22600 7942
rect 23662 7840 23718 8000
rect 24858 7970 24914 8000
rect 24504 7942 24914 7970
rect 23676 7018 23704 7840
rect 23676 6990 23980 7018
rect 23952 6458 23980 6990
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 22560 6452 22612 6458
rect 22560 6394 22612 6400
rect 23940 6452 23992 6458
rect 23940 6394 23992 6400
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 480 2508 532 2514
rect 480 2450 532 2456
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 160 244 2314
rect 492 160 520 2450
rect 1308 2440 1360 2446
rect 1308 2382 1360 2388
rect 756 1896 808 1902
rect 756 1838 808 1844
rect 768 160 796 1838
rect 1032 1828 1084 1834
rect 1032 1770 1084 1776
rect 1044 160 1072 1770
rect 1320 160 1348 2382
rect 1412 1358 1440 2994
rect 1504 1873 1532 6258
rect 5644 6186 5672 6326
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 3917 6012 4225 6021
rect 3917 6010 3923 6012
rect 3979 6010 4003 6012
rect 4059 6010 4083 6012
rect 4139 6010 4163 6012
rect 4219 6010 4225 6012
rect 3979 5958 3981 6010
rect 4161 5958 4163 6010
rect 3917 5956 3923 5958
rect 3979 5956 4003 5958
rect 4059 5956 4083 5958
rect 4139 5956 4163 5958
rect 4219 5956 4225 5958
rect 3917 5947 4225 5956
rect 6564 5914 6592 6258
rect 7576 5914 7604 6258
rect 8772 5914 8800 6258
rect 9692 5914 9720 6258
rect 9851 6012 10159 6021
rect 9851 6010 9857 6012
rect 9913 6010 9937 6012
rect 9993 6010 10017 6012
rect 10073 6010 10097 6012
rect 10153 6010 10159 6012
rect 9913 5958 9915 6010
rect 10095 5958 10097 6010
rect 9851 5956 9857 5958
rect 9913 5956 9937 5958
rect 9993 5956 10017 5958
rect 10073 5956 10097 5958
rect 10153 5956 10159 5958
rect 9851 5947 10159 5956
rect 11164 5914 11192 6258
rect 12360 5914 12388 6258
rect 12636 5914 12664 6258
rect 13556 5914 13584 6258
rect 14660 5914 14688 6258
rect 15120 5914 15148 6258
rect 15672 5914 15700 6258
rect 15785 6012 16093 6021
rect 15785 6010 15791 6012
rect 15847 6010 15871 6012
rect 15927 6010 15951 6012
rect 16007 6010 16031 6012
rect 16087 6010 16093 6012
rect 15847 5958 15849 6010
rect 16029 5958 16031 6010
rect 15785 5956 15791 5958
rect 15847 5956 15871 5958
rect 15927 5956 15951 5958
rect 16007 5956 16031 5958
rect 16087 5956 16093 5958
rect 15785 5947 16093 5956
rect 17420 5914 17448 6258
rect 18340 5914 18368 6258
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 12348 5908 12400 5914
rect 12348 5850 12400 5856
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 18328 5908 18380 5914
rect 18328 5850 18380 5856
rect 19996 5846 20024 6258
rect 20548 5914 20576 6258
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 18420 5704 18472 5710
rect 18420 5646 18472 5652
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 6288 5370 6316 5646
rect 6884 5468 7192 5477
rect 6884 5466 6890 5468
rect 6946 5466 6970 5468
rect 7026 5466 7050 5468
rect 7106 5466 7130 5468
rect 7186 5466 7192 5468
rect 6946 5414 6948 5466
rect 7128 5414 7130 5466
rect 6884 5412 6890 5414
rect 6946 5412 6970 5414
rect 7026 5412 7050 5414
rect 7106 5412 7130 5414
rect 7186 5412 7192 5414
rect 6884 5403 7192 5412
rect 7576 5370 7604 5646
rect 8772 5370 8800 5646
rect 9876 5370 9904 5646
rect 11072 5370 11100 5646
rect 11992 5370 12020 5646
rect 12452 5370 12480 5646
rect 12818 5468 13126 5477
rect 12818 5466 12824 5468
rect 12880 5466 12904 5468
rect 12960 5466 12984 5468
rect 13040 5466 13064 5468
rect 13120 5466 13126 5468
rect 12880 5414 12882 5466
rect 13062 5414 13064 5466
rect 12818 5412 12824 5414
rect 12880 5412 12904 5414
rect 12960 5412 12984 5414
rect 13040 5412 13064 5414
rect 13120 5412 13126 5414
rect 12818 5403 13126 5412
rect 13464 5370 13492 5646
rect 14568 5370 14596 5646
rect 14844 5370 14872 5646
rect 15948 5370 15976 5646
rect 17144 5370 17172 5646
rect 18432 5370 18460 5646
rect 18752 5468 19060 5477
rect 18752 5466 18758 5468
rect 18814 5466 18838 5468
rect 18894 5466 18918 5468
rect 18974 5466 18998 5468
rect 19054 5466 19060 5468
rect 18814 5414 18816 5466
rect 18996 5414 18998 5466
rect 18752 5412 18758 5414
rect 18814 5412 18838 5414
rect 18894 5412 18918 5414
rect 18974 5412 18998 5414
rect 19054 5412 19060 5414
rect 18752 5403 19060 5412
rect 19996 5370 20024 5646
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 18420 5364 18472 5370
rect 18420 5306 18472 5312
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 13176 5296 13228 5302
rect 13176 5238 13228 5244
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 8208 5024 8260 5030
rect 8208 4966 8260 4972
rect 3917 4924 4225 4933
rect 3917 4922 3923 4924
rect 3979 4922 4003 4924
rect 4059 4922 4083 4924
rect 4139 4922 4163 4924
rect 4219 4922 4225 4924
rect 3979 4870 3981 4922
rect 4161 4870 4163 4922
rect 3917 4868 3923 4870
rect 3979 4868 4003 4870
rect 4059 4868 4083 4870
rect 4139 4868 4163 4870
rect 4219 4868 4225 4870
rect 3917 4859 4225 4868
rect 6884 4380 7192 4389
rect 6884 4378 6890 4380
rect 6946 4378 6970 4380
rect 7026 4378 7050 4380
rect 7106 4378 7130 4380
rect 7186 4378 7192 4380
rect 6946 4326 6948 4378
rect 7128 4326 7130 4378
rect 6884 4324 6890 4326
rect 6946 4324 6970 4326
rect 7026 4324 7050 4326
rect 7106 4324 7130 4326
rect 7186 4324 7192 4326
rect 6884 4315 7192 4324
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 3917 3836 4225 3845
rect 3917 3834 3923 3836
rect 3979 3834 4003 3836
rect 4059 3834 4083 3836
rect 4139 3834 4163 3836
rect 4219 3834 4225 3836
rect 3979 3782 3981 3834
rect 4161 3782 4163 3834
rect 3917 3780 3923 3782
rect 3979 3780 4003 3782
rect 4059 3780 4083 3782
rect 4139 3780 4163 3782
rect 4219 3780 4225 3782
rect 3917 3771 4225 3780
rect 6884 3292 7192 3301
rect 6884 3290 6890 3292
rect 6946 3290 6970 3292
rect 7026 3290 7050 3292
rect 7106 3290 7130 3292
rect 7186 3290 7192 3292
rect 6946 3238 6948 3290
rect 7128 3238 7130 3290
rect 6884 3236 6890 3238
rect 6946 3236 6970 3238
rect 7026 3236 7050 3238
rect 7106 3236 7130 3238
rect 7186 3236 7192 3238
rect 6884 3227 7192 3236
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 1952 2848 2004 2854
rect 1952 2790 2004 2796
rect 1964 2582 1992 2790
rect 1584 2576 1636 2582
rect 1582 2544 1584 2553
rect 1952 2576 2004 2582
rect 1636 2544 1638 2553
rect 1952 2518 2004 2524
rect 1582 2479 1638 2488
rect 2596 2508 2648 2514
rect 2596 2450 2648 2456
rect 1952 2372 2004 2378
rect 1952 2314 2004 2320
rect 1768 1964 1820 1970
rect 1768 1906 1820 1912
rect 1490 1864 1546 1873
rect 1490 1799 1546 1808
rect 1492 1760 1544 1766
rect 1492 1702 1544 1708
rect 1504 1358 1532 1702
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 1676 1216 1728 1222
rect 1676 1158 1728 1164
rect 1688 1057 1716 1158
rect 1674 1048 1730 1057
rect 1674 983 1730 992
rect 202 0 258 160
rect 478 0 534 160
rect 754 0 810 160
rect 1030 0 1086 160
rect 1306 0 1362 160
rect 1582 82 1638 160
rect 1780 82 1808 1906
rect 1964 1272 1992 2314
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 1872 1244 1992 1272
rect 1872 160 1900 1244
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 2056 1018 2084 1158
rect 2044 1012 2096 1018
rect 2044 954 2096 960
rect 2148 160 2176 1906
rect 2228 1760 2280 1766
rect 2228 1702 2280 1708
rect 2320 1760 2372 1766
rect 2320 1702 2372 1708
rect 2240 1465 2268 1702
rect 2226 1456 2282 1465
rect 2226 1391 2282 1400
rect 2332 1329 2360 1702
rect 2608 1562 2636 2450
rect 2700 2106 2728 2858
rect 3917 2748 4225 2757
rect 3917 2746 3923 2748
rect 3979 2746 4003 2748
rect 4059 2746 4083 2748
rect 4139 2746 4163 2748
rect 4219 2746 4225 2748
rect 3979 2694 3981 2746
rect 4161 2694 4163 2746
rect 3917 2692 3923 2694
rect 3979 2692 4003 2694
rect 4059 2692 4083 2694
rect 4139 2692 4163 2694
rect 4219 2692 4225 2694
rect 3917 2683 4225 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 2884 1562 2912 2246
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 2964 1760 3016 1766
rect 2964 1702 3016 1708
rect 2596 1556 2648 1562
rect 2596 1498 2648 1504
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 2780 1352 2832 1358
rect 2318 1320 2374 1329
rect 2780 1294 2832 1300
rect 2318 1255 2374 1264
rect 2688 1284 2740 1290
rect 2688 1226 2740 1232
rect 2228 1216 2280 1222
rect 2228 1158 2280 1164
rect 2320 1216 2372 1222
rect 2320 1158 2372 1164
rect 1582 54 1808 82
rect 1582 0 1638 54
rect 1858 0 1914 160
rect 2134 0 2190 160
rect 2240 82 2268 1158
rect 2332 950 2360 1158
rect 2320 944 2372 950
rect 2320 886 2372 892
rect 2700 160 2728 1226
rect 2792 542 2820 1294
rect 2976 1057 3004 1702
rect 3054 1592 3110 1601
rect 3054 1527 3110 1536
rect 3068 1358 3096 1527
rect 3056 1352 3108 1358
rect 3056 1294 3108 1300
rect 2962 1048 3018 1057
rect 2962 983 3018 992
rect 2780 536 2832 542
rect 2780 478 2832 484
rect 2410 82 2466 160
rect 2240 54 2466 82
rect 2410 0 2466 54
rect 2686 0 2742 160
rect 2962 82 3018 160
rect 3160 82 3188 1906
rect 3332 1828 3384 1834
rect 3332 1770 3384 1776
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3252 160 3280 1362
rect 3344 1222 3372 1770
rect 3332 1216 3384 1222
rect 3332 1158 3384 1164
rect 3436 814 3464 2586
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 3528 2060 3924 2088
rect 3528 1442 3556 2060
rect 3608 1964 3660 1970
rect 3792 1964 3844 1970
rect 3660 1924 3740 1952
rect 3608 1906 3660 1912
rect 3608 1828 3660 1834
rect 3608 1770 3660 1776
rect 3620 1601 3648 1770
rect 3606 1592 3662 1601
rect 3606 1527 3662 1536
rect 3528 1414 3648 1442
rect 3516 1352 3568 1358
rect 3516 1294 3568 1300
rect 3528 1222 3556 1294
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3424 808 3476 814
rect 3424 750 3476 756
rect 3620 542 3648 1414
rect 3516 536 3568 542
rect 3516 478 3568 484
rect 3608 536 3660 542
rect 3608 478 3660 484
rect 3528 160 3556 478
rect 2962 54 3188 82
rect 2962 0 3018 54
rect 3238 0 3294 160
rect 3514 0 3570 160
rect 3712 82 3740 1924
rect 3792 1906 3844 1912
rect 3804 490 3832 1906
rect 3896 1748 3924 2060
rect 4264 1970 4292 2246
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4068 1760 4120 1766
rect 3896 1720 4068 1748
rect 4068 1702 4120 1708
rect 4252 1760 4304 1766
rect 4252 1702 4304 1708
rect 3917 1660 4225 1669
rect 3917 1658 3923 1660
rect 3979 1658 4003 1660
rect 4059 1658 4083 1660
rect 4139 1658 4163 1660
rect 4219 1658 4225 1660
rect 3979 1606 3981 1658
rect 4161 1606 4163 1658
rect 3917 1604 3923 1606
rect 3979 1604 4003 1606
rect 4059 1604 4083 1606
rect 4139 1604 4163 1606
rect 4219 1604 4225 1606
rect 3917 1595 4225 1604
rect 3884 1352 3936 1358
rect 4264 1340 4292 1702
rect 4356 1562 4384 2246
rect 4436 1896 4488 1902
rect 4436 1838 4488 1844
rect 4344 1556 4396 1562
rect 4344 1498 4396 1504
rect 3936 1312 4292 1340
rect 3884 1294 3936 1300
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 4344 1216 4396 1222
rect 4344 1158 4396 1164
rect 3988 746 4016 1158
rect 3976 740 4028 746
rect 3976 682 4028 688
rect 3804 462 3924 490
rect 4356 474 4384 1158
rect 3790 82 3846 160
rect 3712 54 3846 82
rect 3896 82 3924 462
rect 4344 468 4396 474
rect 4344 410 4396 416
rect 4066 82 4122 160
rect 3896 54 4122 82
rect 3790 0 3846 54
rect 4066 0 4122 54
rect 4342 82 4398 160
rect 4448 82 4476 1838
rect 4632 160 4660 2382
rect 4712 1964 4764 1970
rect 4712 1906 4764 1912
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 5264 1964 5316 1970
rect 5264 1906 5316 1912
rect 4724 1034 4752 1906
rect 5000 1850 5028 1906
rect 5000 1822 5120 1850
rect 4802 1320 4858 1329
rect 4802 1255 4858 1264
rect 4816 1222 4844 1255
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4724 1006 4936 1034
rect 4908 160 4936 1006
rect 4342 54 4476 82
rect 4342 0 4398 54
rect 4618 0 4674 160
rect 4894 0 4950 160
rect 5092 82 5120 1822
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5184 1358 5212 1702
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 5184 542 5212 1158
rect 5172 536 5224 542
rect 5172 478 5224 484
rect 5170 82 5226 160
rect 5092 54 5226 82
rect 5276 82 5304 1906
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5552 1358 5580 1702
rect 5920 1562 5948 2926
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6274 2408 6330 2417
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 6012 1562 6040 1702
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5448 1216 5500 1222
rect 5448 1158 5500 1164
rect 5540 1216 5592 1222
rect 5592 1176 5764 1204
rect 5540 1158 5592 1164
rect 5460 1018 5488 1158
rect 5448 1012 5500 1018
rect 5448 954 5500 960
rect 5736 160 5764 1176
rect 6104 490 6132 2382
rect 6274 2343 6330 2352
rect 6288 2310 6316 2343
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6748 2088 6776 2790
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7208 2446 7236 2586
rect 7196 2440 7248 2446
rect 7380 2440 7432 2446
rect 7196 2382 7248 2388
rect 7300 2400 7380 2428
rect 6884 2204 7192 2213
rect 6884 2202 6890 2204
rect 6946 2202 6970 2204
rect 7026 2202 7050 2204
rect 7106 2202 7130 2204
rect 7186 2202 7192 2204
rect 6946 2150 6948 2202
rect 7128 2150 7130 2202
rect 6884 2148 6890 2150
rect 6946 2148 6970 2150
rect 7026 2148 7050 2150
rect 7106 2148 7130 2150
rect 7186 2148 7192 2150
rect 6884 2139 7192 2148
rect 6748 2060 7052 2088
rect 6918 2000 6974 2009
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6644 1964 6696 1970
rect 6918 1935 6974 1944
rect 6644 1906 6696 1912
rect 6276 1896 6328 1902
rect 6276 1838 6328 1844
rect 6012 462 6132 490
rect 6012 160 6040 462
rect 6288 160 6316 1838
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6472 1358 6500 1702
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 6368 1216 6420 1222
rect 6368 1158 6420 1164
rect 6380 882 6408 1158
rect 6368 876 6420 882
rect 6368 818 6420 824
rect 6564 160 6592 1906
rect 6656 660 6684 1906
rect 6736 1760 6788 1766
rect 6736 1702 6788 1708
rect 6748 1358 6776 1702
rect 6932 1562 6960 1935
rect 6920 1556 6972 1562
rect 6920 1498 6972 1504
rect 7024 1358 7052 2060
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 7116 1562 7144 1702
rect 7104 1556 7156 1562
rect 7104 1498 7156 1504
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6920 1352 6972 1358
rect 6920 1294 6972 1300
rect 7012 1352 7064 1358
rect 7012 1294 7064 1300
rect 6840 1204 6868 1294
rect 6748 1176 6868 1204
rect 6932 1204 6960 1294
rect 7196 1216 7248 1222
rect 6932 1176 7196 1204
rect 6748 814 6776 1176
rect 7196 1158 7248 1164
rect 6884 1116 7192 1125
rect 6884 1114 6890 1116
rect 6946 1114 6970 1116
rect 7026 1114 7050 1116
rect 7106 1114 7130 1116
rect 7186 1114 7192 1116
rect 6946 1062 6948 1114
rect 7128 1062 7130 1114
rect 6884 1060 6890 1062
rect 6946 1060 6970 1062
rect 7026 1060 7050 1062
rect 7106 1060 7130 1062
rect 7186 1060 7192 1062
rect 6884 1051 7192 1060
rect 7300 932 7328 2400
rect 7380 2382 7432 2388
rect 7484 2106 7512 2858
rect 7562 2136 7618 2145
rect 7472 2100 7524 2106
rect 7562 2071 7618 2080
rect 7472 2042 7524 2048
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7116 904 7328 932
rect 6736 808 6788 814
rect 6736 750 6788 756
rect 6656 632 6868 660
rect 6840 160 6868 632
rect 6918 640 6974 649
rect 6918 575 6920 584
rect 6972 575 6974 584
rect 6920 546 6972 552
rect 7116 160 7144 904
rect 7392 160 7420 1906
rect 7484 1034 7512 1906
rect 7576 1902 7604 2071
rect 7564 1896 7616 1902
rect 7564 1838 7616 1844
rect 7668 1222 7696 4218
rect 8220 4185 8248 4966
rect 9851 4924 10159 4933
rect 9851 4922 9857 4924
rect 9913 4922 9937 4924
rect 9993 4922 10017 4924
rect 10073 4922 10097 4924
rect 10153 4922 10159 4924
rect 9913 4870 9915 4922
rect 10095 4870 10097 4922
rect 9851 4868 9857 4870
rect 9913 4868 9937 4870
rect 9993 4868 10017 4870
rect 10073 4868 10097 4870
rect 10153 4868 10159 4870
rect 9851 4859 10159 4868
rect 8206 4176 8262 4185
rect 8206 4111 8262 4120
rect 9851 3836 10159 3845
rect 9851 3834 9857 3836
rect 9913 3834 9937 3836
rect 9993 3834 10017 3836
rect 10073 3834 10097 3836
rect 10153 3834 10159 3836
rect 9913 3782 9915 3834
rect 10095 3782 10097 3834
rect 9851 3780 9857 3782
rect 9913 3780 9937 3782
rect 9993 3780 10017 3782
rect 10073 3780 10097 3782
rect 10153 3780 10159 3782
rect 9851 3771 10159 3780
rect 10980 3126 11008 5170
rect 10968 3120 11020 3126
rect 8206 3088 8262 3097
rect 10968 3062 11020 3068
rect 11256 3058 11284 5170
rect 12818 4380 13126 4389
rect 12818 4378 12824 4380
rect 12880 4378 12904 4380
rect 12960 4378 12984 4380
rect 13040 4378 13064 4380
rect 13120 4378 13126 4380
rect 12880 4326 12882 4378
rect 13062 4326 13064 4378
rect 12818 4324 12824 4326
rect 12880 4324 12904 4326
rect 12960 4324 12984 4326
rect 13040 4324 13064 4326
rect 13120 4324 13126 4326
rect 12818 4315 13126 4324
rect 12818 3292 13126 3301
rect 12818 3290 12824 3292
rect 12880 3290 12904 3292
rect 12960 3290 12984 3292
rect 13040 3290 13064 3292
rect 13120 3290 13126 3292
rect 12880 3238 12882 3290
rect 13062 3238 13064 3290
rect 12818 3236 12824 3238
rect 12880 3236 12904 3238
rect 12960 3236 12984 3238
rect 13040 3236 13064 3238
rect 13120 3236 13126 3238
rect 12818 3227 13126 3236
rect 8206 3023 8262 3032
rect 10416 3052 10468 3058
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7760 2106 7788 2382
rect 7852 2106 7880 2518
rect 8036 2106 8064 2858
rect 8116 2304 8168 2310
rect 8114 2272 8116 2281
rect 8168 2272 8170 2281
rect 8114 2207 8170 2216
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8220 1986 8248 3023
rect 10416 2994 10468 3000
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9312 2440 9364 2446
rect 9048 2378 9260 2394
rect 9312 2382 9364 2388
rect 9048 2372 9272 2378
rect 9048 2366 9220 2372
rect 8760 2032 8812 2038
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 8128 1958 8248 1986
rect 8588 1992 8760 2020
rect 8300 1964 8352 1970
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7484 1006 7696 1034
rect 7564 808 7616 814
rect 7562 776 7564 785
rect 7616 776 7618 785
rect 7562 711 7618 720
rect 7668 160 7696 1006
rect 7760 728 7788 1906
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 7852 1426 7880 1838
rect 7930 1728 7986 1737
rect 7930 1663 7986 1672
rect 7840 1420 7892 1426
rect 7840 1362 7892 1368
rect 7944 1306 7972 1663
rect 7852 1290 7972 1306
rect 7840 1284 7972 1290
rect 7892 1278 7972 1284
rect 7840 1226 7892 1232
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7944 898 7972 1158
rect 8036 1034 8064 1906
rect 8128 1834 8156 1958
rect 8300 1906 8352 1912
rect 8116 1828 8168 1834
rect 8116 1770 8168 1776
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 8220 1358 8248 1702
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8208 1216 8260 1222
rect 8206 1184 8208 1193
rect 8260 1184 8262 1193
rect 8206 1119 8262 1128
rect 8312 1034 8340 1906
rect 8482 1592 8538 1601
rect 8482 1527 8538 1536
rect 8496 1494 8524 1527
rect 8588 1494 8616 1992
rect 8760 1974 8812 1980
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8484 1488 8536 1494
rect 8484 1430 8536 1436
rect 8576 1488 8628 1494
rect 8576 1430 8628 1436
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8404 1170 8432 1362
rect 8484 1352 8536 1358
rect 8680 1340 8708 1702
rect 8536 1312 8708 1340
rect 8484 1294 8536 1300
rect 8404 1142 8800 1170
rect 8574 1048 8630 1057
rect 8036 1006 8248 1034
rect 8312 1006 8524 1034
rect 7944 870 8064 898
rect 8036 814 8064 870
rect 8024 808 8076 814
rect 8024 750 8076 756
rect 7760 700 7972 728
rect 7944 160 7972 700
rect 8220 160 8248 1006
rect 8496 160 8524 1006
rect 8574 983 8630 992
rect 8588 950 8616 983
rect 8576 944 8628 950
rect 8576 886 8628 892
rect 8772 160 8800 1142
rect 8864 218 8892 1906
rect 9048 1834 9076 2366
rect 9220 2314 9272 2320
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 1970 9168 2246
rect 9128 1964 9180 1970
rect 9128 1906 9180 1912
rect 9036 1828 9088 1834
rect 9036 1770 9088 1776
rect 9218 1728 9274 1737
rect 9218 1663 9274 1672
rect 8942 1592 8998 1601
rect 8942 1527 8998 1536
rect 8956 1494 8984 1527
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 9232 1358 9260 1663
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 9128 1284 9180 1290
rect 9128 1226 9180 1232
rect 8942 1184 8998 1193
rect 8942 1119 8998 1128
rect 8956 338 8984 1119
rect 8944 332 8996 338
rect 8944 274 8996 280
rect 9140 270 9168 1226
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9232 678 9260 1158
rect 9220 672 9272 678
rect 9220 614 9272 620
rect 9128 264 9180 270
rect 8864 190 9076 218
rect 9128 206 9180 212
rect 9048 160 9076 190
rect 9324 160 9352 2382
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 1970 9444 2246
rect 9404 1964 9456 1970
rect 9404 1906 9456 1912
rect 9508 1834 9536 2790
rect 9600 2530 9628 2926
rect 9851 2748 10159 2757
rect 9851 2746 9857 2748
rect 9913 2746 9937 2748
rect 9993 2746 10017 2748
rect 10073 2746 10097 2748
rect 10153 2746 10159 2748
rect 9913 2694 9915 2746
rect 10095 2694 10097 2746
rect 9851 2692 9857 2694
rect 9913 2692 9937 2694
rect 9993 2692 10017 2694
rect 10073 2692 10097 2694
rect 10153 2692 10159 2694
rect 9851 2683 10159 2692
rect 9600 2502 10088 2530
rect 9680 2440 9732 2446
rect 9600 2400 9680 2428
rect 9496 1828 9548 1834
rect 9496 1770 9548 1776
rect 9600 1544 9628 2400
rect 9680 2382 9732 2388
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 9416 1516 9628 1544
rect 9416 1204 9444 1516
rect 9692 1442 9720 1770
rect 9508 1414 9720 1442
rect 9508 1358 9536 1414
rect 9784 1358 9812 2246
rect 10060 1970 10088 2502
rect 10428 2038 10456 2994
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 2394 10732 2586
rect 10796 2582 10824 2926
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 11060 2644 11112 2650
rect 10888 2604 11060 2632
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10888 2514 10916 2604
rect 11060 2586 11112 2592
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 12254 2544 12310 2553
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10980 2394 11008 2450
rect 10416 2032 10468 2038
rect 10230 2000 10286 2009
rect 10048 1964 10100 1970
rect 10416 1974 10468 1980
rect 10230 1935 10286 1944
rect 10324 1964 10376 1970
rect 10048 1906 10100 1912
rect 10244 1737 10272 1935
rect 10324 1906 10376 1912
rect 10230 1728 10286 1737
rect 9851 1660 10159 1669
rect 10230 1663 10286 1672
rect 9851 1658 9857 1660
rect 9913 1658 9937 1660
rect 9993 1658 10017 1660
rect 10073 1658 10097 1660
rect 10153 1658 10159 1660
rect 9913 1606 9915 1658
rect 10095 1606 10097 1658
rect 9851 1604 9857 1606
rect 9913 1604 9937 1606
rect 9993 1604 10017 1606
rect 10073 1604 10097 1606
rect 10153 1604 10159 1606
rect 9851 1595 10159 1604
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9772 1352 9824 1358
rect 9772 1294 9824 1300
rect 9864 1284 9916 1290
rect 9864 1226 9916 1232
rect 9680 1216 9732 1222
rect 9416 1176 9628 1204
rect 9600 160 9628 1176
rect 9680 1158 9732 1164
rect 9692 950 9720 1158
rect 9680 944 9732 950
rect 9680 886 9732 892
rect 9876 542 9904 1226
rect 10048 1216 10100 1222
rect 10048 1158 10100 1164
rect 9864 536 9916 542
rect 9864 478 9916 484
rect 9680 264 9732 270
rect 9732 212 9904 218
rect 9680 206 9904 212
rect 9692 190 9904 206
rect 9876 160 9904 190
rect 5446 82 5502 160
rect 5276 54 5502 82
rect 5170 0 5226 54
rect 5446 0 5502 54
rect 5722 0 5778 160
rect 5998 0 6054 160
rect 6274 0 6330 160
rect 6550 0 6606 160
rect 6826 0 6882 160
rect 7102 0 7158 160
rect 7378 0 7434 160
rect 7654 0 7710 160
rect 7930 0 7986 160
rect 8206 0 8262 160
rect 8482 0 8538 160
rect 8758 0 8814 160
rect 9034 0 9090 160
rect 9310 0 9366 160
rect 9586 0 9642 160
rect 9862 0 9918 160
rect 10060 82 10088 1158
rect 10336 1057 10364 1906
rect 10508 1760 10560 1766
rect 10428 1720 10508 1748
rect 10322 1048 10378 1057
rect 10322 983 10378 992
rect 10428 160 10456 1720
rect 10508 1702 10560 1708
rect 10612 649 10640 2382
rect 10704 2366 11008 2394
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 10692 1284 10744 1290
rect 10692 1226 10744 1232
rect 10784 1284 10836 1290
rect 10784 1226 10836 1232
rect 10598 640 10654 649
rect 10598 575 10654 584
rect 10704 160 10732 1226
rect 10796 1018 10824 1226
rect 10888 1018 10916 2246
rect 11244 2032 11296 2038
rect 11244 1974 11296 1980
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 10784 1012 10836 1018
rect 10784 954 10836 960
rect 10876 1012 10928 1018
rect 10876 954 10928 960
rect 10980 160 11008 1702
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 10138 82 10194 160
rect 10060 54 10194 82
rect 10138 0 10194 54
rect 10414 0 10470 160
rect 10690 0 10746 160
rect 10966 0 11022 160
rect 11072 82 11100 1362
rect 11152 1216 11204 1222
rect 11152 1158 11204 1164
rect 11164 354 11192 1158
rect 11256 542 11284 1974
rect 11336 1964 11388 1970
rect 11336 1906 11388 1912
rect 11348 785 11376 1906
rect 11532 1426 11560 2246
rect 11808 2009 11836 2382
rect 11794 2000 11850 2009
rect 11794 1935 11850 1944
rect 11716 1822 11928 1850
rect 11716 1766 11744 1822
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 11704 1352 11756 1358
rect 11702 1320 11704 1329
rect 11756 1320 11758 1329
rect 11702 1255 11758 1264
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11624 882 11652 1158
rect 11612 876 11664 882
rect 11612 818 11664 824
rect 11334 776 11390 785
rect 11334 711 11390 720
rect 11244 536 11296 542
rect 11244 478 11296 484
rect 11164 326 11560 354
rect 11532 160 11560 326
rect 11808 160 11836 1702
rect 11242 82 11298 160
rect 11072 54 11298 82
rect 11242 0 11298 54
rect 11518 0 11574 160
rect 11794 0 11850 160
rect 11900 82 11928 1822
rect 11992 1494 12020 2518
rect 12254 2479 12310 2488
rect 12072 2304 12124 2310
rect 12268 2281 12296 2479
rect 12348 2304 12400 2310
rect 12072 2246 12124 2252
rect 12254 2272 12310 2281
rect 12084 1902 12112 2246
rect 12348 2246 12400 2252
rect 12254 2207 12310 2216
rect 12360 1970 12388 2246
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12452 1714 12480 2790
rect 12532 2440 12584 2446
rect 12584 2400 12756 2428
rect 12532 2382 12584 2388
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12636 2106 12664 2246
rect 12624 2100 12676 2106
rect 12624 2042 12676 2048
rect 12452 1686 12572 1714
rect 12544 1494 12572 1686
rect 11980 1488 12032 1494
rect 11980 1430 12032 1436
rect 12532 1488 12584 1494
rect 12532 1430 12584 1436
rect 12440 1352 12492 1358
rect 12728 1329 12756 2400
rect 12818 2204 13126 2213
rect 12818 2202 12824 2204
rect 12880 2202 12904 2204
rect 12960 2202 12984 2204
rect 13040 2202 13064 2204
rect 13120 2202 13126 2204
rect 12880 2150 12882 2202
rect 13062 2150 13064 2202
rect 12818 2148 12824 2150
rect 12880 2148 12904 2150
rect 12960 2148 12984 2150
rect 13040 2148 13064 2150
rect 13120 2148 13126 2150
rect 12818 2139 13126 2148
rect 13188 1884 13216 5238
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 13648 3466 13676 5170
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13452 2508 13504 2514
rect 13452 2450 13504 2456
rect 13188 1856 13400 1884
rect 12808 1760 12860 1766
rect 12808 1702 12860 1708
rect 12900 1760 12952 1766
rect 12900 1702 12952 1708
rect 12820 1426 12848 1702
rect 12808 1420 12860 1426
rect 12808 1362 12860 1368
rect 12440 1294 12492 1300
rect 12714 1320 12770 1329
rect 12072 1216 12124 1222
rect 12072 1158 12124 1164
rect 12348 1216 12400 1222
rect 12348 1158 12400 1164
rect 12084 406 12112 1158
rect 12072 400 12124 406
rect 12072 342 12124 348
rect 12360 160 12388 1158
rect 12452 746 12480 1294
rect 12714 1255 12770 1264
rect 12912 1204 12940 1702
rect 12636 1176 12940 1204
rect 13084 1216 13136 1222
rect 12440 740 12492 746
rect 12440 682 12492 688
rect 12636 160 12664 1176
rect 13136 1176 13216 1204
rect 13084 1158 13136 1164
rect 12818 1116 13126 1125
rect 12818 1114 12824 1116
rect 12880 1114 12904 1116
rect 12960 1114 12984 1116
rect 13040 1114 13064 1116
rect 13120 1114 13126 1116
rect 12880 1062 12882 1114
rect 13062 1062 13064 1114
rect 12818 1060 12824 1062
rect 12880 1060 12904 1062
rect 12960 1060 12984 1062
rect 13040 1060 13064 1062
rect 13120 1060 13126 1062
rect 12818 1051 13126 1060
rect 12900 740 12952 746
rect 12900 682 12952 688
rect 12912 160 12940 682
rect 13188 160 13216 1176
rect 13372 542 13400 1856
rect 13464 1834 13492 2450
rect 14004 2304 14056 2310
rect 14004 2246 14056 2252
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14016 2106 14044 2246
rect 14004 2100 14056 2106
rect 14004 2042 14056 2048
rect 14108 1986 14136 2246
rect 14016 1970 14136 1986
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 14004 1964 14136 1970
rect 14056 1958 14136 1964
rect 14004 1906 14056 1912
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13452 1216 13504 1222
rect 13452 1158 13504 1164
rect 13360 536 13412 542
rect 13360 478 13412 484
rect 13464 160 13492 1158
rect 13556 678 13584 1906
rect 13820 1760 13872 1766
rect 13872 1708 13952 1714
rect 13820 1702 13952 1708
rect 13832 1686 13952 1702
rect 13820 1556 13872 1562
rect 13740 1516 13820 1544
rect 13544 672 13596 678
rect 13544 614 13596 620
rect 13740 160 13768 1516
rect 13820 1498 13872 1504
rect 13924 1358 13952 1686
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 14016 160 14044 1158
rect 14200 882 14228 5102
rect 14370 2680 14426 2689
rect 14370 2615 14426 2624
rect 14384 1970 14412 2615
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14292 1850 14320 1906
rect 14292 1822 14412 1850
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 14188 876 14240 882
rect 14188 818 14240 824
rect 14292 160 14320 1702
rect 14384 1465 14412 1822
rect 14370 1456 14426 1465
rect 14370 1391 14426 1400
rect 14476 746 14504 5170
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 15785 4924 16093 4933
rect 15785 4922 15791 4924
rect 15847 4922 15871 4924
rect 15927 4922 15951 4924
rect 16007 4922 16031 4924
rect 16087 4922 16093 4924
rect 15847 4870 15849 4922
rect 16029 4870 16031 4922
rect 15785 4868 15791 4870
rect 15847 4868 15871 4870
rect 15927 4868 15951 4870
rect 16007 4868 16031 4870
rect 16087 4868 16093 4870
rect 15785 4859 16093 4868
rect 17144 4214 17172 5102
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 15785 3836 16093 3845
rect 15785 3834 15791 3836
rect 15847 3834 15871 3836
rect 15927 3834 15951 3836
rect 16007 3834 16031 3836
rect 16087 3834 16093 3836
rect 15847 3782 15849 3834
rect 16029 3782 16031 3834
rect 15785 3780 15791 3782
rect 15847 3780 15871 3782
rect 15927 3780 15951 3782
rect 16007 3780 16031 3782
rect 16087 3780 16093 3782
rect 15785 3771 16093 3780
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 14660 950 14688 1294
rect 14648 944 14700 950
rect 14648 886 14700 892
rect 14464 740 14516 746
rect 14464 682 14516 688
rect 12070 82 12126 160
rect 11900 54 12126 82
rect 12070 0 12126 54
rect 12346 0 12402 160
rect 12622 0 12678 160
rect 12898 0 12954 160
rect 13174 0 13230 160
rect 13450 0 13506 160
rect 13726 0 13782 160
rect 14002 0 14058 160
rect 14278 0 14334 160
rect 14554 82 14610 160
rect 14752 82 14780 1702
rect 14924 1556 14976 1562
rect 14844 1516 14924 1544
rect 14844 160 14872 1516
rect 14924 1498 14976 1504
rect 15028 1222 15056 2858
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 1970 15148 2246
rect 15108 1964 15160 1970
rect 15108 1906 15160 1912
rect 15212 1544 15240 2994
rect 15785 2748 16093 2757
rect 15785 2746 15791 2748
rect 15847 2746 15871 2748
rect 15927 2746 15951 2748
rect 16007 2746 16031 2748
rect 16087 2746 16093 2748
rect 15847 2694 15849 2746
rect 16029 2694 16031 2746
rect 15785 2692 15791 2694
rect 15847 2692 15871 2694
rect 15927 2692 15951 2694
rect 16007 2692 16031 2694
rect 16087 2692 16093 2694
rect 15785 2683 16093 2692
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15304 2106 15332 2382
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15396 2106 15424 2246
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15384 1828 15436 1834
rect 15384 1770 15436 1776
rect 15120 1516 15240 1544
rect 15120 1306 15148 1516
rect 15292 1488 15344 1494
rect 15292 1430 15344 1436
rect 15120 1278 15240 1306
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15212 678 15240 1278
rect 15200 672 15252 678
rect 15200 614 15252 620
rect 15304 524 15332 1430
rect 15396 1426 15424 1770
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15384 1420 15436 1426
rect 15384 1362 15436 1368
rect 15488 1358 15516 1702
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 15580 1170 15608 2246
rect 16040 2038 16068 2450
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 16304 2304 16356 2310
rect 16304 2246 16356 2252
rect 16028 2032 16080 2038
rect 16028 1974 16080 1980
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 15660 1760 15712 1766
rect 15660 1702 15712 1708
rect 15120 496 15332 524
rect 15396 1142 15608 1170
rect 15120 160 15148 496
rect 15396 160 15424 1142
rect 15672 160 15700 1702
rect 15785 1660 16093 1669
rect 15785 1658 15791 1660
rect 15847 1658 15871 1660
rect 15927 1658 15951 1660
rect 16007 1658 16031 1660
rect 16087 1658 16093 1660
rect 15847 1606 15849 1658
rect 16029 1606 16031 1658
rect 15785 1604 15791 1606
rect 15847 1604 15871 1606
rect 15927 1604 15951 1606
rect 16007 1604 16031 1606
rect 16087 1604 16093 1606
rect 15785 1595 16093 1604
rect 16028 1488 16080 1494
rect 16028 1430 16080 1436
rect 16040 626 16068 1430
rect 15948 598 16068 626
rect 16132 610 16160 1906
rect 16212 1420 16264 1426
rect 16212 1362 16264 1368
rect 16120 604 16172 610
rect 15948 160 15976 598
rect 16120 546 16172 552
rect 16224 160 16252 1362
rect 16316 270 16344 2246
rect 16500 1562 16528 2382
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 16592 1358 16620 1702
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16396 1284 16448 1290
rect 16396 1226 16448 1232
rect 16408 1018 16436 1226
rect 16488 1216 16540 1222
rect 16488 1158 16540 1164
rect 16396 1012 16448 1018
rect 16396 954 16448 960
rect 16304 264 16356 270
rect 16304 206 16356 212
rect 16500 160 16528 1158
rect 16684 950 16712 3062
rect 17236 2990 17264 4966
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16764 2848 16816 2854
rect 16764 2790 16816 2796
rect 16776 2446 16804 2790
rect 17880 2650 17908 4150
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17868 2644 17920 2650
rect 17868 2586 17920 2592
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16856 2304 16908 2310
rect 16856 2246 16908 2252
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16764 1760 16816 1766
rect 16764 1702 16816 1708
rect 16672 944 16724 950
rect 16672 886 16724 892
rect 16776 160 16804 1702
rect 16868 1358 16896 2246
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16960 1018 16988 2246
rect 17420 1290 17448 2586
rect 17972 2514 18000 4150
rect 18616 2582 18644 5170
rect 18752 4380 19060 4389
rect 18752 4378 18758 4380
rect 18814 4378 18838 4380
rect 18894 4378 18918 4380
rect 18974 4378 18998 4380
rect 19054 4378 19060 4380
rect 18814 4326 18816 4378
rect 18996 4326 18998 4378
rect 18752 4324 18758 4326
rect 18814 4324 18838 4326
rect 18894 4324 18918 4326
rect 18974 4324 18998 4326
rect 19054 4324 19060 4326
rect 18752 4315 19060 4324
rect 18752 3292 19060 3301
rect 18752 3290 18758 3292
rect 18814 3290 18838 3292
rect 18894 3290 18918 3292
rect 18974 3290 18998 3292
rect 19054 3290 19060 3292
rect 18814 3238 18816 3290
rect 18996 3238 18998 3290
rect 18752 3236 18758 3238
rect 18814 3236 18838 3238
rect 18894 3236 18918 3238
rect 18974 3236 18998 3238
rect 19054 3236 19060 3238
rect 18752 3227 19060 3236
rect 18604 2576 18656 2582
rect 18142 2544 18198 2553
rect 17960 2508 18012 2514
rect 18604 2518 18656 2524
rect 18142 2479 18198 2488
rect 20088 2502 20484 2530
rect 17960 2450 18012 2456
rect 18156 2446 18184 2479
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18420 2440 18472 2446
rect 18696 2440 18748 2446
rect 18420 2382 18472 2388
rect 18524 2400 18696 2428
rect 17604 2106 17632 2382
rect 17776 2304 17828 2310
rect 17776 2246 17828 2252
rect 17592 2100 17644 2106
rect 17592 2042 17644 2048
rect 17788 2038 17816 2246
rect 17880 2106 17908 2382
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18236 2304 18288 2310
rect 18236 2246 18288 2252
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17776 1828 17828 1834
rect 17696 1788 17776 1816
rect 17592 1556 17644 1562
rect 17512 1516 17592 1544
rect 17408 1284 17460 1290
rect 17408 1226 17460 1232
rect 16948 1012 17000 1018
rect 16948 954 17000 960
rect 17512 728 17540 1516
rect 17592 1498 17644 1504
rect 17592 1420 17644 1426
rect 17592 1362 17644 1368
rect 17052 700 17540 728
rect 17052 160 17080 700
rect 17604 626 17632 1362
rect 17328 598 17632 626
rect 17328 160 17356 598
rect 17696 524 17724 1788
rect 17776 1770 17828 1776
rect 17880 1822 18000 1850
rect 17604 496 17724 524
rect 17604 160 17632 496
rect 17880 160 17908 1822
rect 17972 1766 18000 1822
rect 17960 1760 18012 1766
rect 17960 1702 18012 1708
rect 18156 1426 18184 2246
rect 18248 2106 18276 2246
rect 18340 2106 18368 2314
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18328 2100 18380 2106
rect 18328 2042 18380 2048
rect 18432 1970 18460 2382
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18236 1760 18288 1766
rect 18236 1702 18288 1708
rect 18144 1420 18196 1426
rect 18144 1362 18196 1368
rect 18248 898 18276 1702
rect 18524 1465 18552 2400
rect 19708 2440 19760 2446
rect 18696 2382 18748 2388
rect 19706 2408 19708 2417
rect 19760 2408 19762 2417
rect 19706 2343 19762 2352
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 18616 1578 18644 2246
rect 18752 2204 19060 2213
rect 18752 2202 18758 2204
rect 18814 2202 18838 2204
rect 18894 2202 18918 2204
rect 18974 2202 18998 2204
rect 19054 2202 19060 2204
rect 18814 2150 18816 2202
rect 18996 2150 18998 2202
rect 18752 2148 18758 2150
rect 18814 2148 18838 2150
rect 18894 2148 18918 2150
rect 18974 2148 18998 2150
rect 19054 2148 19060 2150
rect 18752 2139 19060 2148
rect 19168 2106 19196 2246
rect 19260 2106 19288 2246
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19892 2032 19944 2038
rect 19892 1974 19944 1980
rect 19432 1828 19484 1834
rect 19432 1770 19484 1776
rect 19340 1760 19392 1766
rect 19340 1702 19392 1708
rect 18616 1550 18828 1578
rect 18696 1488 18748 1494
rect 18510 1456 18566 1465
rect 18696 1430 18748 1436
rect 18510 1391 18566 1400
rect 18604 1420 18656 1426
rect 18604 1362 18656 1368
rect 18512 1284 18564 1290
rect 18156 870 18276 898
rect 18432 1244 18512 1272
rect 18156 160 18184 870
rect 18432 160 18460 1244
rect 18512 1226 18564 1232
rect 18616 728 18644 1362
rect 18708 1290 18736 1430
rect 18696 1284 18748 1290
rect 18696 1226 18748 1232
rect 18800 1204 18828 1550
rect 19352 1442 19380 1702
rect 19168 1414 19380 1442
rect 19064 1216 19116 1222
rect 18800 1176 19064 1204
rect 19064 1158 19116 1164
rect 18752 1116 19060 1125
rect 18752 1114 18758 1116
rect 18814 1114 18838 1116
rect 18894 1114 18918 1116
rect 18974 1114 18998 1116
rect 19054 1114 19060 1116
rect 18814 1062 18816 1114
rect 18996 1062 18998 1114
rect 18752 1060 18758 1062
rect 18814 1060 18838 1062
rect 18894 1060 18918 1062
rect 18974 1060 18998 1062
rect 19054 1060 19060 1062
rect 18752 1051 19060 1060
rect 19168 898 19196 1414
rect 19444 1306 19472 1770
rect 19904 1714 19932 1974
rect 18984 870 19196 898
rect 19260 1278 19472 1306
rect 19720 1686 19932 1714
rect 19616 1284 19668 1290
rect 18616 700 18736 728
rect 18708 160 18736 700
rect 18984 160 19012 870
rect 19260 160 19288 1278
rect 19616 1226 19668 1232
rect 19628 1018 19656 1226
rect 19616 1012 19668 1018
rect 19616 954 19668 960
rect 14554 54 14780 82
rect 14554 0 14610 54
rect 14830 0 14886 160
rect 15106 0 15162 160
rect 15382 0 15438 160
rect 15658 0 15714 160
rect 15934 0 15990 160
rect 16210 0 16266 160
rect 16486 0 16542 160
rect 16762 0 16818 160
rect 17038 0 17094 160
rect 17314 0 17370 160
rect 17590 0 17646 160
rect 17866 0 17922 160
rect 18142 0 18198 160
rect 18418 0 18474 160
rect 18694 0 18750 160
rect 18970 0 19026 160
rect 19246 0 19302 160
rect 19522 82 19578 160
rect 19720 82 19748 1686
rect 19800 1556 19852 1562
rect 19800 1498 19852 1504
rect 19812 160 19840 1498
rect 19996 1358 20024 2246
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 20088 160 20116 2502
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20180 1465 20208 2382
rect 20272 2009 20300 2382
rect 20456 2378 20484 2502
rect 20444 2372 20496 2378
rect 20444 2314 20496 2320
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20364 2106 20392 2246
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20640 2038 20668 2246
rect 21192 2106 21220 5170
rect 21652 2106 21680 6190
rect 21719 6012 22027 6021
rect 21719 6010 21725 6012
rect 21781 6010 21805 6012
rect 21861 6010 21885 6012
rect 21941 6010 21965 6012
rect 22021 6010 22027 6012
rect 21781 5958 21783 6010
rect 21963 5958 21965 6010
rect 21719 5956 21725 5958
rect 21781 5956 21805 5958
rect 21861 5956 21885 5958
rect 21941 5956 21965 5958
rect 22021 5956 22027 5958
rect 21719 5947 22027 5956
rect 22560 5092 22612 5098
rect 22560 5034 22612 5040
rect 21719 4924 22027 4933
rect 21719 4922 21725 4924
rect 21781 4922 21805 4924
rect 21861 4922 21885 4924
rect 21941 4922 21965 4924
rect 22021 4922 22027 4924
rect 21781 4870 21783 4922
rect 21963 4870 21965 4922
rect 21719 4868 21725 4870
rect 21781 4868 21805 4870
rect 21861 4868 21885 4870
rect 21941 4868 21965 4870
rect 22021 4868 22027 4870
rect 21719 4859 22027 4868
rect 21719 3836 22027 3845
rect 21719 3834 21725 3836
rect 21781 3834 21805 3836
rect 21861 3834 21885 3836
rect 21941 3834 21965 3836
rect 22021 3834 22027 3836
rect 21781 3782 21783 3834
rect 21963 3782 21965 3834
rect 21719 3780 21725 3782
rect 21781 3780 21805 3782
rect 21861 3780 21885 3782
rect 21941 3780 21965 3782
rect 22021 3780 22027 3782
rect 21719 3771 22027 3780
rect 22192 3460 22244 3466
rect 22192 3402 22244 3408
rect 21719 2748 22027 2757
rect 21719 2746 21725 2748
rect 21781 2746 21805 2748
rect 21861 2746 21885 2748
rect 21941 2746 21965 2748
rect 22021 2746 22027 2748
rect 21781 2694 21783 2746
rect 21963 2694 21965 2746
rect 21719 2692 21725 2694
rect 21781 2692 21805 2694
rect 21861 2692 21885 2694
rect 21941 2692 21965 2694
rect 22021 2692 22027 2694
rect 21719 2683 22027 2692
rect 21088 2100 21140 2106
rect 21088 2042 21140 2048
rect 21180 2100 21232 2106
rect 21180 2042 21232 2048
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 20628 2032 20680 2038
rect 20258 2000 20314 2009
rect 20628 1974 20680 1980
rect 21100 1970 21128 2042
rect 20258 1935 20314 1944
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 21272 1964 21324 1970
rect 21272 1906 21324 1912
rect 22008 1964 22060 1970
rect 22008 1906 22060 1912
rect 20902 1864 20958 1873
rect 20902 1799 20958 1808
rect 21180 1828 21232 1834
rect 20916 1766 20944 1799
rect 21180 1770 21232 1776
rect 20904 1760 20956 1766
rect 20904 1702 20956 1708
rect 21192 1562 21220 1770
rect 21180 1556 21232 1562
rect 21180 1498 21232 1504
rect 20166 1456 20222 1465
rect 20166 1391 20222 1400
rect 20536 1216 20588 1222
rect 20536 1158 20588 1164
rect 20352 672 20404 678
rect 20352 614 20404 620
rect 20364 160 20392 614
rect 19522 54 19748 82
rect 19522 0 19578 54
rect 19798 0 19854 160
rect 20074 0 20130 160
rect 20350 0 20406 160
rect 20548 82 20576 1158
rect 20904 808 20956 814
rect 20904 750 20956 756
rect 20916 160 20944 750
rect 21284 678 21312 1906
rect 21732 1896 21784 1902
rect 21652 1856 21732 1884
rect 21548 1488 21600 1494
rect 21548 1430 21600 1436
rect 21456 1420 21508 1426
rect 21456 1362 21508 1368
rect 21468 1193 21496 1362
rect 21454 1184 21510 1193
rect 21454 1119 21510 1128
rect 21560 762 21588 1430
rect 21376 734 21588 762
rect 21272 672 21324 678
rect 21272 614 21324 620
rect 20626 82 20682 160
rect 20548 54 20682 82
rect 20626 0 20682 54
rect 20902 0 20958 160
rect 21178 82 21234 160
rect 21376 82 21404 734
rect 21456 672 21508 678
rect 21456 614 21508 620
rect 21468 160 21496 614
rect 21178 54 21404 82
rect 21178 0 21234 54
rect 21454 0 21510 160
rect 21652 82 21680 1856
rect 21732 1838 21784 1844
rect 22020 1850 22048 1906
rect 22204 1902 22232 3402
rect 22284 2984 22336 2990
rect 22284 2926 22336 2932
rect 22296 2106 22324 2926
rect 22376 2440 22428 2446
rect 22376 2382 22428 2388
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 22388 1902 22416 2382
rect 22468 1964 22520 1970
rect 22468 1906 22520 1912
rect 22192 1896 22244 1902
rect 22020 1822 22140 1850
rect 22192 1838 22244 1844
rect 22376 1896 22428 1902
rect 22376 1838 22428 1844
rect 21719 1660 22027 1669
rect 21719 1658 21725 1660
rect 21781 1658 21805 1660
rect 21861 1658 21885 1660
rect 21941 1658 21965 1660
rect 22021 1658 22027 1660
rect 21781 1606 21783 1658
rect 21963 1606 21965 1658
rect 21719 1604 21725 1606
rect 21781 1604 21805 1606
rect 21861 1604 21885 1606
rect 21941 1604 21965 1606
rect 22021 1604 22027 1606
rect 21719 1595 22027 1604
rect 22112 1562 22140 1822
rect 22100 1556 22152 1562
rect 22100 1498 22152 1504
rect 21824 1488 21876 1494
rect 21822 1456 21824 1465
rect 22008 1488 22060 1494
rect 21876 1456 21878 1465
rect 22008 1430 22060 1436
rect 21822 1391 21878 1400
rect 21732 1352 21784 1358
rect 21730 1320 21732 1329
rect 21784 1320 21786 1329
rect 21730 1255 21786 1264
rect 21916 1216 21968 1222
rect 21744 1176 21916 1204
rect 21744 814 21772 1176
rect 21916 1158 21968 1164
rect 21916 1012 21968 1018
rect 21916 954 21968 960
rect 21732 808 21784 814
rect 21732 750 21784 756
rect 21928 542 21956 954
rect 21916 536 21968 542
rect 21916 478 21968 484
rect 22020 160 22048 1430
rect 22284 1216 22336 1222
rect 22284 1158 22336 1164
rect 22296 814 22324 1158
rect 22374 1048 22430 1057
rect 22374 983 22430 992
rect 22284 808 22336 814
rect 22284 750 22336 756
rect 21730 82 21786 160
rect 21652 54 21786 82
rect 21730 0 21786 54
rect 22006 0 22062 160
rect 22282 82 22338 160
rect 22388 82 22416 983
rect 22480 762 22508 1906
rect 22572 1358 22600 5034
rect 22928 4616 22980 4622
rect 22928 4558 22980 4564
rect 22836 2848 22888 2854
rect 22836 2790 22888 2796
rect 22848 2446 22876 2790
rect 22940 2650 22968 4558
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 22836 2440 22888 2446
rect 22836 2382 22888 2388
rect 22744 2304 22796 2310
rect 22744 2246 22796 2252
rect 22756 1970 22784 2246
rect 23124 2106 23152 6258
rect 23676 3738 23704 6258
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 24032 5840 24084 5846
rect 24032 5782 24084 5788
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23860 5370 23888 5578
rect 23848 5364 23900 5370
rect 23848 5306 23900 5312
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23388 2440 23440 2446
rect 23440 2388 23520 2394
rect 23388 2382 23520 2388
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 22744 1964 22796 1970
rect 23020 1964 23072 1970
rect 22744 1906 22796 1912
rect 22848 1924 23020 1952
rect 22560 1352 22612 1358
rect 22744 1352 22796 1358
rect 22560 1294 22612 1300
rect 22650 1320 22706 1329
rect 22706 1300 22744 1306
rect 22706 1294 22796 1300
rect 22706 1278 22784 1294
rect 22650 1255 22706 1264
rect 22742 1184 22798 1193
rect 22742 1119 22798 1128
rect 22480 734 22692 762
rect 22664 406 22692 734
rect 22652 400 22704 406
rect 22652 342 22704 348
rect 22282 54 22416 82
rect 22558 82 22614 160
rect 22756 82 22784 1119
rect 22848 160 22876 1924
rect 23020 1906 23072 1912
rect 23112 1896 23164 1902
rect 23164 1856 23244 1884
rect 23112 1838 23164 1844
rect 22928 1352 22980 1358
rect 22928 1294 22980 1300
rect 22940 814 22968 1294
rect 23112 1216 23164 1222
rect 23112 1158 23164 1164
rect 23124 1018 23152 1158
rect 23112 1012 23164 1018
rect 23112 954 23164 960
rect 23216 898 23244 1856
rect 23124 870 23244 898
rect 22928 808 22980 814
rect 22928 750 22980 756
rect 23124 160 23152 870
rect 23308 814 23336 2382
rect 23400 2366 23520 2382
rect 23388 2032 23440 2038
rect 23388 1974 23440 1980
rect 23296 808 23348 814
rect 23296 750 23348 756
rect 23400 160 23428 1974
rect 23492 1834 23520 2366
rect 23480 1828 23532 1834
rect 23480 1770 23532 1776
rect 23676 1578 23704 2790
rect 23768 2650 23796 5102
rect 24044 3074 24072 5782
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 24136 3194 24164 3470
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 24044 3046 24164 3074
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 24044 2446 24072 2790
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24032 2440 24084 2446
rect 24032 2382 24084 2388
rect 23756 1828 23808 1834
rect 23756 1770 23808 1776
rect 23492 1550 23704 1578
rect 23492 1494 23520 1550
rect 23768 1494 23796 1770
rect 23480 1488 23532 1494
rect 23480 1430 23532 1436
rect 23756 1488 23808 1494
rect 23756 1430 23808 1436
rect 23848 1352 23900 1358
rect 23584 1278 23796 1306
rect 23848 1294 23900 1300
rect 23584 746 23612 1278
rect 23768 1222 23796 1278
rect 23664 1216 23716 1222
rect 23664 1158 23716 1164
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23676 1018 23704 1158
rect 23860 1057 23888 1294
rect 23846 1048 23902 1057
rect 23664 1012 23716 1018
rect 23846 983 23902 992
rect 23664 954 23716 960
rect 23952 898 23980 2382
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24044 2106 24072 2246
rect 24032 2100 24084 2106
rect 24032 2042 24084 2048
rect 24136 1766 24164 3046
rect 24228 2394 24256 6122
rect 24504 5914 24532 7942
rect 24858 7840 24914 7942
rect 24686 6556 24994 6565
rect 24686 6554 24692 6556
rect 24748 6554 24772 6556
rect 24828 6554 24852 6556
rect 24908 6554 24932 6556
rect 24988 6554 24994 6556
rect 24748 6502 24750 6554
rect 24930 6502 24932 6554
rect 24686 6500 24692 6502
rect 24748 6500 24772 6502
rect 24828 6500 24852 6502
rect 24908 6500 24932 6502
rect 24988 6500 24994 6502
rect 24686 6491 24994 6500
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24686 5468 24994 5477
rect 24686 5466 24692 5468
rect 24748 5466 24772 5468
rect 24828 5466 24852 5468
rect 24908 5466 24932 5468
rect 24988 5466 24994 5468
rect 24748 5414 24750 5466
rect 24930 5414 24932 5466
rect 24686 5412 24692 5414
rect 24748 5412 24772 5414
rect 24828 5412 24852 5414
rect 24908 5412 24932 5414
rect 24988 5412 24994 5414
rect 24686 5403 24994 5412
rect 24400 5296 24452 5302
rect 24400 5238 24452 5244
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24320 4826 24348 5170
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24308 3052 24360 3058
rect 24308 2994 24360 3000
rect 24320 2650 24348 2994
rect 24308 2644 24360 2650
rect 24308 2586 24360 2592
rect 24228 2366 24348 2394
rect 24216 2304 24268 2310
rect 24216 2246 24268 2252
rect 24124 1760 24176 1766
rect 24124 1702 24176 1708
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 24044 1193 24072 1294
rect 24030 1184 24086 1193
rect 24030 1119 24086 1128
rect 24228 1034 24256 2246
rect 24320 1902 24348 2366
rect 24412 2106 24440 5238
rect 24686 4380 24994 4389
rect 24686 4378 24692 4380
rect 24748 4378 24772 4380
rect 24828 4378 24852 4380
rect 24908 4378 24932 4380
rect 24988 4378 24994 4380
rect 24748 4326 24750 4378
rect 24930 4326 24932 4378
rect 24686 4324 24692 4326
rect 24748 4324 24772 4326
rect 24828 4324 24852 4326
rect 24908 4324 24932 4326
rect 24988 4324 24994 4326
rect 24686 4315 24994 4324
rect 24686 3292 24994 3301
rect 24686 3290 24692 3292
rect 24748 3290 24772 3292
rect 24828 3290 24852 3292
rect 24908 3290 24932 3292
rect 24988 3290 24994 3292
rect 24748 3238 24750 3290
rect 24930 3238 24932 3290
rect 24686 3236 24692 3238
rect 24748 3236 24772 3238
rect 24828 3236 24852 3238
rect 24908 3236 24932 3238
rect 24988 3236 24994 3238
rect 24686 3227 24994 3236
rect 25044 3120 25096 3126
rect 25044 3062 25096 3068
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24400 2100 24452 2106
rect 24400 2042 24452 2048
rect 24308 1896 24360 1902
rect 24308 1838 24360 1844
rect 24308 1216 24360 1222
rect 24308 1158 24360 1164
rect 23676 870 23980 898
rect 24044 1006 24256 1034
rect 24320 1018 24348 1158
rect 24308 1012 24360 1018
rect 23572 740 23624 746
rect 23572 682 23624 688
rect 23676 160 23704 870
rect 24044 796 24072 1006
rect 24308 954 24360 960
rect 23952 768 24072 796
rect 23952 160 23980 768
rect 24216 400 24268 406
rect 24216 342 24268 348
rect 24228 160 24256 342
rect 24504 160 24532 2926
rect 24584 2916 24636 2922
rect 24584 2858 24636 2864
rect 22558 54 22784 82
rect 22282 0 22338 54
rect 22558 0 22614 54
rect 22834 0 22890 160
rect 23110 0 23166 160
rect 23386 0 23442 160
rect 23662 0 23718 160
rect 23938 0 23994 160
rect 24214 0 24270 160
rect 24490 0 24546 160
rect 24596 82 24624 2858
rect 24686 2204 24994 2213
rect 24686 2202 24692 2204
rect 24748 2202 24772 2204
rect 24828 2202 24852 2204
rect 24908 2202 24932 2204
rect 24988 2202 24994 2204
rect 24748 2150 24750 2202
rect 24930 2150 24932 2202
rect 24686 2148 24692 2150
rect 24748 2148 24772 2150
rect 24828 2148 24852 2150
rect 24908 2148 24932 2150
rect 24988 2148 24994 2150
rect 24686 2139 24994 2148
rect 24686 1116 24994 1125
rect 24686 1114 24692 1116
rect 24748 1114 24772 1116
rect 24828 1114 24852 1116
rect 24908 1114 24932 1116
rect 24988 1114 24994 1116
rect 24748 1062 24750 1114
rect 24930 1062 24932 1114
rect 24686 1060 24692 1062
rect 24748 1060 24772 1062
rect 24828 1060 24852 1062
rect 24908 1060 24932 1062
rect 24988 1060 24994 1062
rect 24686 1051 24994 1060
rect 25056 160 25084 3062
rect 25320 1488 25372 1494
rect 25320 1430 25372 1436
rect 25332 160 25360 1430
rect 25596 808 25648 814
rect 25596 750 25648 756
rect 25608 160 25636 750
rect 24766 82 24822 160
rect 24596 54 24822 82
rect 24766 0 24822 54
rect 25042 0 25098 160
rect 25318 0 25374 160
rect 25594 0 25650 160
<< via2 >>
rect 6890 6554 6946 6556
rect 6970 6554 7026 6556
rect 7050 6554 7106 6556
rect 7130 6554 7186 6556
rect 6890 6502 6936 6554
rect 6936 6502 6946 6554
rect 6970 6502 7000 6554
rect 7000 6502 7012 6554
rect 7012 6502 7026 6554
rect 7050 6502 7064 6554
rect 7064 6502 7076 6554
rect 7076 6502 7106 6554
rect 7130 6502 7140 6554
rect 7140 6502 7186 6554
rect 6890 6500 6946 6502
rect 6970 6500 7026 6502
rect 7050 6500 7106 6502
rect 7130 6500 7186 6502
rect 12824 6554 12880 6556
rect 12904 6554 12960 6556
rect 12984 6554 13040 6556
rect 13064 6554 13120 6556
rect 12824 6502 12870 6554
rect 12870 6502 12880 6554
rect 12904 6502 12934 6554
rect 12934 6502 12946 6554
rect 12946 6502 12960 6554
rect 12984 6502 12998 6554
rect 12998 6502 13010 6554
rect 13010 6502 13040 6554
rect 13064 6502 13074 6554
rect 13074 6502 13120 6554
rect 12824 6500 12880 6502
rect 12904 6500 12960 6502
rect 12984 6500 13040 6502
rect 13064 6500 13120 6502
rect 18758 6554 18814 6556
rect 18838 6554 18894 6556
rect 18918 6554 18974 6556
rect 18998 6554 19054 6556
rect 18758 6502 18804 6554
rect 18804 6502 18814 6554
rect 18838 6502 18868 6554
rect 18868 6502 18880 6554
rect 18880 6502 18894 6554
rect 18918 6502 18932 6554
rect 18932 6502 18944 6554
rect 18944 6502 18974 6554
rect 18998 6502 19008 6554
rect 19008 6502 19054 6554
rect 18758 6500 18814 6502
rect 18838 6500 18894 6502
rect 18918 6500 18974 6502
rect 18998 6500 19054 6502
rect 3923 6010 3979 6012
rect 4003 6010 4059 6012
rect 4083 6010 4139 6012
rect 4163 6010 4219 6012
rect 3923 5958 3969 6010
rect 3969 5958 3979 6010
rect 4003 5958 4033 6010
rect 4033 5958 4045 6010
rect 4045 5958 4059 6010
rect 4083 5958 4097 6010
rect 4097 5958 4109 6010
rect 4109 5958 4139 6010
rect 4163 5958 4173 6010
rect 4173 5958 4219 6010
rect 3923 5956 3979 5958
rect 4003 5956 4059 5958
rect 4083 5956 4139 5958
rect 4163 5956 4219 5958
rect 9857 6010 9913 6012
rect 9937 6010 9993 6012
rect 10017 6010 10073 6012
rect 10097 6010 10153 6012
rect 9857 5958 9903 6010
rect 9903 5958 9913 6010
rect 9937 5958 9967 6010
rect 9967 5958 9979 6010
rect 9979 5958 9993 6010
rect 10017 5958 10031 6010
rect 10031 5958 10043 6010
rect 10043 5958 10073 6010
rect 10097 5958 10107 6010
rect 10107 5958 10153 6010
rect 9857 5956 9913 5958
rect 9937 5956 9993 5958
rect 10017 5956 10073 5958
rect 10097 5956 10153 5958
rect 15791 6010 15847 6012
rect 15871 6010 15927 6012
rect 15951 6010 16007 6012
rect 16031 6010 16087 6012
rect 15791 5958 15837 6010
rect 15837 5958 15847 6010
rect 15871 5958 15901 6010
rect 15901 5958 15913 6010
rect 15913 5958 15927 6010
rect 15951 5958 15965 6010
rect 15965 5958 15977 6010
rect 15977 5958 16007 6010
rect 16031 5958 16041 6010
rect 16041 5958 16087 6010
rect 15791 5956 15847 5958
rect 15871 5956 15927 5958
rect 15951 5956 16007 5958
rect 16031 5956 16087 5958
rect 6890 5466 6946 5468
rect 6970 5466 7026 5468
rect 7050 5466 7106 5468
rect 7130 5466 7186 5468
rect 6890 5414 6936 5466
rect 6936 5414 6946 5466
rect 6970 5414 7000 5466
rect 7000 5414 7012 5466
rect 7012 5414 7026 5466
rect 7050 5414 7064 5466
rect 7064 5414 7076 5466
rect 7076 5414 7106 5466
rect 7130 5414 7140 5466
rect 7140 5414 7186 5466
rect 6890 5412 6946 5414
rect 6970 5412 7026 5414
rect 7050 5412 7106 5414
rect 7130 5412 7186 5414
rect 12824 5466 12880 5468
rect 12904 5466 12960 5468
rect 12984 5466 13040 5468
rect 13064 5466 13120 5468
rect 12824 5414 12870 5466
rect 12870 5414 12880 5466
rect 12904 5414 12934 5466
rect 12934 5414 12946 5466
rect 12946 5414 12960 5466
rect 12984 5414 12998 5466
rect 12998 5414 13010 5466
rect 13010 5414 13040 5466
rect 13064 5414 13074 5466
rect 13074 5414 13120 5466
rect 12824 5412 12880 5414
rect 12904 5412 12960 5414
rect 12984 5412 13040 5414
rect 13064 5412 13120 5414
rect 18758 5466 18814 5468
rect 18838 5466 18894 5468
rect 18918 5466 18974 5468
rect 18998 5466 19054 5468
rect 18758 5414 18804 5466
rect 18804 5414 18814 5466
rect 18838 5414 18868 5466
rect 18868 5414 18880 5466
rect 18880 5414 18894 5466
rect 18918 5414 18932 5466
rect 18932 5414 18944 5466
rect 18944 5414 18974 5466
rect 18998 5414 19008 5466
rect 19008 5414 19054 5466
rect 18758 5412 18814 5414
rect 18838 5412 18894 5414
rect 18918 5412 18974 5414
rect 18998 5412 19054 5414
rect 3923 4922 3979 4924
rect 4003 4922 4059 4924
rect 4083 4922 4139 4924
rect 4163 4922 4219 4924
rect 3923 4870 3969 4922
rect 3969 4870 3979 4922
rect 4003 4870 4033 4922
rect 4033 4870 4045 4922
rect 4045 4870 4059 4922
rect 4083 4870 4097 4922
rect 4097 4870 4109 4922
rect 4109 4870 4139 4922
rect 4163 4870 4173 4922
rect 4173 4870 4219 4922
rect 3923 4868 3979 4870
rect 4003 4868 4059 4870
rect 4083 4868 4139 4870
rect 4163 4868 4219 4870
rect 6890 4378 6946 4380
rect 6970 4378 7026 4380
rect 7050 4378 7106 4380
rect 7130 4378 7186 4380
rect 6890 4326 6936 4378
rect 6936 4326 6946 4378
rect 6970 4326 7000 4378
rect 7000 4326 7012 4378
rect 7012 4326 7026 4378
rect 7050 4326 7064 4378
rect 7064 4326 7076 4378
rect 7076 4326 7106 4378
rect 7130 4326 7140 4378
rect 7140 4326 7186 4378
rect 6890 4324 6946 4326
rect 6970 4324 7026 4326
rect 7050 4324 7106 4326
rect 7130 4324 7186 4326
rect 3923 3834 3979 3836
rect 4003 3834 4059 3836
rect 4083 3834 4139 3836
rect 4163 3834 4219 3836
rect 3923 3782 3969 3834
rect 3969 3782 3979 3834
rect 4003 3782 4033 3834
rect 4033 3782 4045 3834
rect 4045 3782 4059 3834
rect 4083 3782 4097 3834
rect 4097 3782 4109 3834
rect 4109 3782 4139 3834
rect 4163 3782 4173 3834
rect 4173 3782 4219 3834
rect 3923 3780 3979 3782
rect 4003 3780 4059 3782
rect 4083 3780 4139 3782
rect 4163 3780 4219 3782
rect 6890 3290 6946 3292
rect 6970 3290 7026 3292
rect 7050 3290 7106 3292
rect 7130 3290 7186 3292
rect 6890 3238 6936 3290
rect 6936 3238 6946 3290
rect 6970 3238 7000 3290
rect 7000 3238 7012 3290
rect 7012 3238 7026 3290
rect 7050 3238 7064 3290
rect 7064 3238 7076 3290
rect 7076 3238 7106 3290
rect 7130 3238 7140 3290
rect 7140 3238 7186 3290
rect 6890 3236 6946 3238
rect 6970 3236 7026 3238
rect 7050 3236 7106 3238
rect 7130 3236 7186 3238
rect 1582 2524 1584 2544
rect 1584 2524 1636 2544
rect 1636 2524 1638 2544
rect 1582 2488 1638 2524
rect 1490 1808 1546 1864
rect 1674 992 1730 1048
rect 2226 1400 2282 1456
rect 3923 2746 3979 2748
rect 4003 2746 4059 2748
rect 4083 2746 4139 2748
rect 4163 2746 4219 2748
rect 3923 2694 3969 2746
rect 3969 2694 3979 2746
rect 4003 2694 4033 2746
rect 4033 2694 4045 2746
rect 4045 2694 4059 2746
rect 4083 2694 4097 2746
rect 4097 2694 4109 2746
rect 4109 2694 4139 2746
rect 4163 2694 4173 2746
rect 4173 2694 4219 2746
rect 3923 2692 3979 2694
rect 4003 2692 4059 2694
rect 4083 2692 4139 2694
rect 4163 2692 4219 2694
rect 2318 1264 2374 1320
rect 3054 1536 3110 1592
rect 2962 992 3018 1048
rect 3606 1536 3662 1592
rect 3923 1658 3979 1660
rect 4003 1658 4059 1660
rect 4083 1658 4139 1660
rect 4163 1658 4219 1660
rect 3923 1606 3969 1658
rect 3969 1606 3979 1658
rect 4003 1606 4033 1658
rect 4033 1606 4045 1658
rect 4045 1606 4059 1658
rect 4083 1606 4097 1658
rect 4097 1606 4109 1658
rect 4109 1606 4139 1658
rect 4163 1606 4173 1658
rect 4173 1606 4219 1658
rect 3923 1604 3979 1606
rect 4003 1604 4059 1606
rect 4083 1604 4139 1606
rect 4163 1604 4219 1606
rect 4802 1264 4858 1320
rect 6274 2352 6330 2408
rect 6890 2202 6946 2204
rect 6970 2202 7026 2204
rect 7050 2202 7106 2204
rect 7130 2202 7186 2204
rect 6890 2150 6936 2202
rect 6936 2150 6946 2202
rect 6970 2150 7000 2202
rect 7000 2150 7012 2202
rect 7012 2150 7026 2202
rect 7050 2150 7064 2202
rect 7064 2150 7076 2202
rect 7076 2150 7106 2202
rect 7130 2150 7140 2202
rect 7140 2150 7186 2202
rect 6890 2148 6946 2150
rect 6970 2148 7026 2150
rect 7050 2148 7106 2150
rect 7130 2148 7186 2150
rect 6918 1944 6974 2000
rect 6890 1114 6946 1116
rect 6970 1114 7026 1116
rect 7050 1114 7106 1116
rect 7130 1114 7186 1116
rect 6890 1062 6936 1114
rect 6936 1062 6946 1114
rect 6970 1062 7000 1114
rect 7000 1062 7012 1114
rect 7012 1062 7026 1114
rect 7050 1062 7064 1114
rect 7064 1062 7076 1114
rect 7076 1062 7106 1114
rect 7130 1062 7140 1114
rect 7140 1062 7186 1114
rect 6890 1060 6946 1062
rect 6970 1060 7026 1062
rect 7050 1060 7106 1062
rect 7130 1060 7186 1062
rect 7562 2080 7618 2136
rect 6918 604 6974 640
rect 6918 584 6920 604
rect 6920 584 6972 604
rect 6972 584 6974 604
rect 9857 4922 9913 4924
rect 9937 4922 9993 4924
rect 10017 4922 10073 4924
rect 10097 4922 10153 4924
rect 9857 4870 9903 4922
rect 9903 4870 9913 4922
rect 9937 4870 9967 4922
rect 9967 4870 9979 4922
rect 9979 4870 9993 4922
rect 10017 4870 10031 4922
rect 10031 4870 10043 4922
rect 10043 4870 10073 4922
rect 10097 4870 10107 4922
rect 10107 4870 10153 4922
rect 9857 4868 9913 4870
rect 9937 4868 9993 4870
rect 10017 4868 10073 4870
rect 10097 4868 10153 4870
rect 8206 4120 8262 4176
rect 9857 3834 9913 3836
rect 9937 3834 9993 3836
rect 10017 3834 10073 3836
rect 10097 3834 10153 3836
rect 9857 3782 9903 3834
rect 9903 3782 9913 3834
rect 9937 3782 9967 3834
rect 9967 3782 9979 3834
rect 9979 3782 9993 3834
rect 10017 3782 10031 3834
rect 10031 3782 10043 3834
rect 10043 3782 10073 3834
rect 10097 3782 10107 3834
rect 10107 3782 10153 3834
rect 9857 3780 9913 3782
rect 9937 3780 9993 3782
rect 10017 3780 10073 3782
rect 10097 3780 10153 3782
rect 8206 3032 8262 3088
rect 12824 4378 12880 4380
rect 12904 4378 12960 4380
rect 12984 4378 13040 4380
rect 13064 4378 13120 4380
rect 12824 4326 12870 4378
rect 12870 4326 12880 4378
rect 12904 4326 12934 4378
rect 12934 4326 12946 4378
rect 12946 4326 12960 4378
rect 12984 4326 12998 4378
rect 12998 4326 13010 4378
rect 13010 4326 13040 4378
rect 13064 4326 13074 4378
rect 13074 4326 13120 4378
rect 12824 4324 12880 4326
rect 12904 4324 12960 4326
rect 12984 4324 13040 4326
rect 13064 4324 13120 4326
rect 12824 3290 12880 3292
rect 12904 3290 12960 3292
rect 12984 3290 13040 3292
rect 13064 3290 13120 3292
rect 12824 3238 12870 3290
rect 12870 3238 12880 3290
rect 12904 3238 12934 3290
rect 12934 3238 12946 3290
rect 12946 3238 12960 3290
rect 12984 3238 12998 3290
rect 12998 3238 13010 3290
rect 13010 3238 13040 3290
rect 13064 3238 13074 3290
rect 13074 3238 13120 3290
rect 12824 3236 12880 3238
rect 12904 3236 12960 3238
rect 12984 3236 13040 3238
rect 13064 3236 13120 3238
rect 8114 2252 8116 2272
rect 8116 2252 8168 2272
rect 8168 2252 8170 2272
rect 8114 2216 8170 2252
rect 7562 756 7564 776
rect 7564 756 7616 776
rect 7616 756 7618 776
rect 7562 720 7618 756
rect 7930 1672 7986 1728
rect 8206 1164 8208 1184
rect 8208 1164 8260 1184
rect 8260 1164 8262 1184
rect 8206 1128 8262 1164
rect 8482 1536 8538 1592
rect 8574 992 8630 1048
rect 9218 1672 9274 1728
rect 8942 1536 8998 1592
rect 8942 1128 8998 1184
rect 9857 2746 9913 2748
rect 9937 2746 9993 2748
rect 10017 2746 10073 2748
rect 10097 2746 10153 2748
rect 9857 2694 9903 2746
rect 9903 2694 9913 2746
rect 9937 2694 9967 2746
rect 9967 2694 9979 2746
rect 9979 2694 9993 2746
rect 10017 2694 10031 2746
rect 10031 2694 10043 2746
rect 10043 2694 10073 2746
rect 10097 2694 10107 2746
rect 10107 2694 10153 2746
rect 9857 2692 9913 2694
rect 9937 2692 9993 2694
rect 10017 2692 10073 2694
rect 10097 2692 10153 2694
rect 10230 1944 10286 2000
rect 10230 1672 10286 1728
rect 9857 1658 9913 1660
rect 9937 1658 9993 1660
rect 10017 1658 10073 1660
rect 10097 1658 10153 1660
rect 9857 1606 9903 1658
rect 9903 1606 9913 1658
rect 9937 1606 9967 1658
rect 9967 1606 9979 1658
rect 9979 1606 9993 1658
rect 10017 1606 10031 1658
rect 10031 1606 10043 1658
rect 10043 1606 10073 1658
rect 10097 1606 10107 1658
rect 10107 1606 10153 1658
rect 9857 1604 9913 1606
rect 9937 1604 9993 1606
rect 10017 1604 10073 1606
rect 10097 1604 10153 1606
rect 10322 992 10378 1048
rect 10598 584 10654 640
rect 11794 1944 11850 2000
rect 11702 1300 11704 1320
rect 11704 1300 11756 1320
rect 11756 1300 11758 1320
rect 11702 1264 11758 1300
rect 11334 720 11390 776
rect 12254 2488 12310 2544
rect 12254 2216 12310 2272
rect 12824 2202 12880 2204
rect 12904 2202 12960 2204
rect 12984 2202 13040 2204
rect 13064 2202 13120 2204
rect 12824 2150 12870 2202
rect 12870 2150 12880 2202
rect 12904 2150 12934 2202
rect 12934 2150 12946 2202
rect 12946 2150 12960 2202
rect 12984 2150 12998 2202
rect 12998 2150 13010 2202
rect 13010 2150 13040 2202
rect 13064 2150 13074 2202
rect 13074 2150 13120 2202
rect 12824 2148 12880 2150
rect 12904 2148 12960 2150
rect 12984 2148 13040 2150
rect 13064 2148 13120 2150
rect 12714 1264 12770 1320
rect 12824 1114 12880 1116
rect 12904 1114 12960 1116
rect 12984 1114 13040 1116
rect 13064 1114 13120 1116
rect 12824 1062 12870 1114
rect 12870 1062 12880 1114
rect 12904 1062 12934 1114
rect 12934 1062 12946 1114
rect 12946 1062 12960 1114
rect 12984 1062 12998 1114
rect 12998 1062 13010 1114
rect 13010 1062 13040 1114
rect 13064 1062 13074 1114
rect 13074 1062 13120 1114
rect 12824 1060 12880 1062
rect 12904 1060 12960 1062
rect 12984 1060 13040 1062
rect 13064 1060 13120 1062
rect 14370 2624 14426 2680
rect 14370 1400 14426 1456
rect 15791 4922 15847 4924
rect 15871 4922 15927 4924
rect 15951 4922 16007 4924
rect 16031 4922 16087 4924
rect 15791 4870 15837 4922
rect 15837 4870 15847 4922
rect 15871 4870 15901 4922
rect 15901 4870 15913 4922
rect 15913 4870 15927 4922
rect 15951 4870 15965 4922
rect 15965 4870 15977 4922
rect 15977 4870 16007 4922
rect 16031 4870 16041 4922
rect 16041 4870 16087 4922
rect 15791 4868 15847 4870
rect 15871 4868 15927 4870
rect 15951 4868 16007 4870
rect 16031 4868 16087 4870
rect 15791 3834 15847 3836
rect 15871 3834 15927 3836
rect 15951 3834 16007 3836
rect 16031 3834 16087 3836
rect 15791 3782 15837 3834
rect 15837 3782 15847 3834
rect 15871 3782 15901 3834
rect 15901 3782 15913 3834
rect 15913 3782 15927 3834
rect 15951 3782 15965 3834
rect 15965 3782 15977 3834
rect 15977 3782 16007 3834
rect 16031 3782 16041 3834
rect 16041 3782 16087 3834
rect 15791 3780 15847 3782
rect 15871 3780 15927 3782
rect 15951 3780 16007 3782
rect 16031 3780 16087 3782
rect 15791 2746 15847 2748
rect 15871 2746 15927 2748
rect 15951 2746 16007 2748
rect 16031 2746 16087 2748
rect 15791 2694 15837 2746
rect 15837 2694 15847 2746
rect 15871 2694 15901 2746
rect 15901 2694 15913 2746
rect 15913 2694 15927 2746
rect 15951 2694 15965 2746
rect 15965 2694 15977 2746
rect 15977 2694 16007 2746
rect 16031 2694 16041 2746
rect 16041 2694 16087 2746
rect 15791 2692 15847 2694
rect 15871 2692 15927 2694
rect 15951 2692 16007 2694
rect 16031 2692 16087 2694
rect 15791 1658 15847 1660
rect 15871 1658 15927 1660
rect 15951 1658 16007 1660
rect 16031 1658 16087 1660
rect 15791 1606 15837 1658
rect 15837 1606 15847 1658
rect 15871 1606 15901 1658
rect 15901 1606 15913 1658
rect 15913 1606 15927 1658
rect 15951 1606 15965 1658
rect 15965 1606 15977 1658
rect 15977 1606 16007 1658
rect 16031 1606 16041 1658
rect 16041 1606 16087 1658
rect 15791 1604 15847 1606
rect 15871 1604 15927 1606
rect 15951 1604 16007 1606
rect 16031 1604 16087 1606
rect 18758 4378 18814 4380
rect 18838 4378 18894 4380
rect 18918 4378 18974 4380
rect 18998 4378 19054 4380
rect 18758 4326 18804 4378
rect 18804 4326 18814 4378
rect 18838 4326 18868 4378
rect 18868 4326 18880 4378
rect 18880 4326 18894 4378
rect 18918 4326 18932 4378
rect 18932 4326 18944 4378
rect 18944 4326 18974 4378
rect 18998 4326 19008 4378
rect 19008 4326 19054 4378
rect 18758 4324 18814 4326
rect 18838 4324 18894 4326
rect 18918 4324 18974 4326
rect 18998 4324 19054 4326
rect 18758 3290 18814 3292
rect 18838 3290 18894 3292
rect 18918 3290 18974 3292
rect 18998 3290 19054 3292
rect 18758 3238 18804 3290
rect 18804 3238 18814 3290
rect 18838 3238 18868 3290
rect 18868 3238 18880 3290
rect 18880 3238 18894 3290
rect 18918 3238 18932 3290
rect 18932 3238 18944 3290
rect 18944 3238 18974 3290
rect 18998 3238 19008 3290
rect 19008 3238 19054 3290
rect 18758 3236 18814 3238
rect 18838 3236 18894 3238
rect 18918 3236 18974 3238
rect 18998 3236 19054 3238
rect 18142 2488 18198 2544
rect 19706 2388 19708 2408
rect 19708 2388 19760 2408
rect 19760 2388 19762 2408
rect 19706 2352 19762 2388
rect 18758 2202 18814 2204
rect 18838 2202 18894 2204
rect 18918 2202 18974 2204
rect 18998 2202 19054 2204
rect 18758 2150 18804 2202
rect 18804 2150 18814 2202
rect 18838 2150 18868 2202
rect 18868 2150 18880 2202
rect 18880 2150 18894 2202
rect 18918 2150 18932 2202
rect 18932 2150 18944 2202
rect 18944 2150 18974 2202
rect 18998 2150 19008 2202
rect 19008 2150 19054 2202
rect 18758 2148 18814 2150
rect 18838 2148 18894 2150
rect 18918 2148 18974 2150
rect 18998 2148 19054 2150
rect 18510 1400 18566 1456
rect 18758 1114 18814 1116
rect 18838 1114 18894 1116
rect 18918 1114 18974 1116
rect 18998 1114 19054 1116
rect 18758 1062 18804 1114
rect 18804 1062 18814 1114
rect 18838 1062 18868 1114
rect 18868 1062 18880 1114
rect 18880 1062 18894 1114
rect 18918 1062 18932 1114
rect 18932 1062 18944 1114
rect 18944 1062 18974 1114
rect 18998 1062 19008 1114
rect 19008 1062 19054 1114
rect 18758 1060 18814 1062
rect 18838 1060 18894 1062
rect 18918 1060 18974 1062
rect 18998 1060 19054 1062
rect 21725 6010 21781 6012
rect 21805 6010 21861 6012
rect 21885 6010 21941 6012
rect 21965 6010 22021 6012
rect 21725 5958 21771 6010
rect 21771 5958 21781 6010
rect 21805 5958 21835 6010
rect 21835 5958 21847 6010
rect 21847 5958 21861 6010
rect 21885 5958 21899 6010
rect 21899 5958 21911 6010
rect 21911 5958 21941 6010
rect 21965 5958 21975 6010
rect 21975 5958 22021 6010
rect 21725 5956 21781 5958
rect 21805 5956 21861 5958
rect 21885 5956 21941 5958
rect 21965 5956 22021 5958
rect 21725 4922 21781 4924
rect 21805 4922 21861 4924
rect 21885 4922 21941 4924
rect 21965 4922 22021 4924
rect 21725 4870 21771 4922
rect 21771 4870 21781 4922
rect 21805 4870 21835 4922
rect 21835 4870 21847 4922
rect 21847 4870 21861 4922
rect 21885 4870 21899 4922
rect 21899 4870 21911 4922
rect 21911 4870 21941 4922
rect 21965 4870 21975 4922
rect 21975 4870 22021 4922
rect 21725 4868 21781 4870
rect 21805 4868 21861 4870
rect 21885 4868 21941 4870
rect 21965 4868 22021 4870
rect 21725 3834 21781 3836
rect 21805 3834 21861 3836
rect 21885 3834 21941 3836
rect 21965 3834 22021 3836
rect 21725 3782 21771 3834
rect 21771 3782 21781 3834
rect 21805 3782 21835 3834
rect 21835 3782 21847 3834
rect 21847 3782 21861 3834
rect 21885 3782 21899 3834
rect 21899 3782 21911 3834
rect 21911 3782 21941 3834
rect 21965 3782 21975 3834
rect 21975 3782 22021 3834
rect 21725 3780 21781 3782
rect 21805 3780 21861 3782
rect 21885 3780 21941 3782
rect 21965 3780 22021 3782
rect 21725 2746 21781 2748
rect 21805 2746 21861 2748
rect 21885 2746 21941 2748
rect 21965 2746 22021 2748
rect 21725 2694 21771 2746
rect 21771 2694 21781 2746
rect 21805 2694 21835 2746
rect 21835 2694 21847 2746
rect 21847 2694 21861 2746
rect 21885 2694 21899 2746
rect 21899 2694 21911 2746
rect 21911 2694 21941 2746
rect 21965 2694 21975 2746
rect 21975 2694 22021 2746
rect 21725 2692 21781 2694
rect 21805 2692 21861 2694
rect 21885 2692 21941 2694
rect 21965 2692 22021 2694
rect 20258 1944 20314 2000
rect 20902 1808 20958 1864
rect 20166 1400 20222 1456
rect 21454 1128 21510 1184
rect 21725 1658 21781 1660
rect 21805 1658 21861 1660
rect 21885 1658 21941 1660
rect 21965 1658 22021 1660
rect 21725 1606 21771 1658
rect 21771 1606 21781 1658
rect 21805 1606 21835 1658
rect 21835 1606 21847 1658
rect 21847 1606 21861 1658
rect 21885 1606 21899 1658
rect 21899 1606 21911 1658
rect 21911 1606 21941 1658
rect 21965 1606 21975 1658
rect 21975 1606 22021 1658
rect 21725 1604 21781 1606
rect 21805 1604 21861 1606
rect 21885 1604 21941 1606
rect 21965 1604 22021 1606
rect 21822 1436 21824 1456
rect 21824 1436 21876 1456
rect 21876 1436 21878 1456
rect 21822 1400 21878 1436
rect 21730 1300 21732 1320
rect 21732 1300 21784 1320
rect 21784 1300 21786 1320
rect 21730 1264 21786 1300
rect 22374 992 22430 1048
rect 22650 1264 22706 1320
rect 22742 1128 22798 1184
rect 23846 992 23902 1048
rect 24692 6554 24748 6556
rect 24772 6554 24828 6556
rect 24852 6554 24908 6556
rect 24932 6554 24988 6556
rect 24692 6502 24738 6554
rect 24738 6502 24748 6554
rect 24772 6502 24802 6554
rect 24802 6502 24814 6554
rect 24814 6502 24828 6554
rect 24852 6502 24866 6554
rect 24866 6502 24878 6554
rect 24878 6502 24908 6554
rect 24932 6502 24942 6554
rect 24942 6502 24988 6554
rect 24692 6500 24748 6502
rect 24772 6500 24828 6502
rect 24852 6500 24908 6502
rect 24932 6500 24988 6502
rect 24692 5466 24748 5468
rect 24772 5466 24828 5468
rect 24852 5466 24908 5468
rect 24932 5466 24988 5468
rect 24692 5414 24738 5466
rect 24738 5414 24748 5466
rect 24772 5414 24802 5466
rect 24802 5414 24814 5466
rect 24814 5414 24828 5466
rect 24852 5414 24866 5466
rect 24866 5414 24878 5466
rect 24878 5414 24908 5466
rect 24932 5414 24942 5466
rect 24942 5414 24988 5466
rect 24692 5412 24748 5414
rect 24772 5412 24828 5414
rect 24852 5412 24908 5414
rect 24932 5412 24988 5414
rect 24030 1128 24086 1184
rect 24692 4378 24748 4380
rect 24772 4378 24828 4380
rect 24852 4378 24908 4380
rect 24932 4378 24988 4380
rect 24692 4326 24738 4378
rect 24738 4326 24748 4378
rect 24772 4326 24802 4378
rect 24802 4326 24814 4378
rect 24814 4326 24828 4378
rect 24852 4326 24866 4378
rect 24866 4326 24878 4378
rect 24878 4326 24908 4378
rect 24932 4326 24942 4378
rect 24942 4326 24988 4378
rect 24692 4324 24748 4326
rect 24772 4324 24828 4326
rect 24852 4324 24908 4326
rect 24932 4324 24988 4326
rect 24692 3290 24748 3292
rect 24772 3290 24828 3292
rect 24852 3290 24908 3292
rect 24932 3290 24988 3292
rect 24692 3238 24738 3290
rect 24738 3238 24748 3290
rect 24772 3238 24802 3290
rect 24802 3238 24814 3290
rect 24814 3238 24828 3290
rect 24852 3238 24866 3290
rect 24866 3238 24878 3290
rect 24878 3238 24908 3290
rect 24932 3238 24942 3290
rect 24942 3238 24988 3290
rect 24692 3236 24748 3238
rect 24772 3236 24828 3238
rect 24852 3236 24908 3238
rect 24932 3236 24988 3238
rect 24692 2202 24748 2204
rect 24772 2202 24828 2204
rect 24852 2202 24908 2204
rect 24932 2202 24988 2204
rect 24692 2150 24738 2202
rect 24738 2150 24748 2202
rect 24772 2150 24802 2202
rect 24802 2150 24814 2202
rect 24814 2150 24828 2202
rect 24852 2150 24866 2202
rect 24866 2150 24878 2202
rect 24878 2150 24908 2202
rect 24932 2150 24942 2202
rect 24942 2150 24988 2202
rect 24692 2148 24748 2150
rect 24772 2148 24828 2150
rect 24852 2148 24908 2150
rect 24932 2148 24988 2150
rect 24692 1114 24748 1116
rect 24772 1114 24828 1116
rect 24852 1114 24908 1116
rect 24932 1114 24988 1116
rect 24692 1062 24738 1114
rect 24738 1062 24748 1114
rect 24772 1062 24802 1114
rect 24802 1062 24814 1114
rect 24814 1062 24828 1114
rect 24852 1062 24866 1114
rect 24866 1062 24878 1114
rect 24878 1062 24908 1114
rect 24932 1062 24942 1114
rect 24942 1062 24988 1114
rect 24692 1060 24748 1062
rect 24772 1060 24828 1062
rect 24852 1060 24908 1062
rect 24932 1060 24988 1062
<< metal3 >>
rect 6880 6560 7196 6561
rect 6880 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7196 6560
rect 6880 6495 7196 6496
rect 12814 6560 13130 6561
rect 12814 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13130 6560
rect 12814 6495 13130 6496
rect 18748 6560 19064 6561
rect 18748 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19064 6560
rect 18748 6495 19064 6496
rect 24682 6560 24998 6561
rect 24682 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 24998 6560
rect 24682 6495 24998 6496
rect 3913 6016 4229 6017
rect 3913 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4229 6016
rect 3913 5951 4229 5952
rect 9847 6016 10163 6017
rect 9847 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10163 6016
rect 9847 5951 10163 5952
rect 15781 6016 16097 6017
rect 15781 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16097 6016
rect 15781 5951 16097 5952
rect 21715 6016 22031 6017
rect 21715 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22031 6016
rect 21715 5951 22031 5952
rect 6880 5472 7196 5473
rect 6880 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7196 5472
rect 6880 5407 7196 5408
rect 12814 5472 13130 5473
rect 12814 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13130 5472
rect 12814 5407 13130 5408
rect 18748 5472 19064 5473
rect 18748 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19064 5472
rect 18748 5407 19064 5408
rect 24682 5472 24998 5473
rect 24682 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 24998 5472
rect 24682 5407 24998 5408
rect 3913 4928 4229 4929
rect 3913 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4229 4928
rect 3913 4863 4229 4864
rect 9847 4928 10163 4929
rect 9847 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10163 4928
rect 9847 4863 10163 4864
rect 15781 4928 16097 4929
rect 15781 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16097 4928
rect 15781 4863 16097 4864
rect 21715 4928 22031 4929
rect 21715 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22031 4928
rect 21715 4863 22031 4864
rect 6880 4384 7196 4385
rect 6880 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7196 4384
rect 6880 4319 7196 4320
rect 12814 4384 13130 4385
rect 12814 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13130 4384
rect 12814 4319 13130 4320
rect 18748 4384 19064 4385
rect 18748 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19064 4384
rect 18748 4319 19064 4320
rect 24682 4384 24998 4385
rect 24682 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 24998 4384
rect 24682 4319 24998 4320
rect 8201 4178 8267 4181
rect 22134 4178 22140 4180
rect 8201 4176 22140 4178
rect 8201 4120 8206 4176
rect 8262 4120 22140 4176
rect 8201 4118 22140 4120
rect 8201 4115 8267 4118
rect 22134 4116 22140 4118
rect 22204 4116 22210 4180
rect 3913 3840 4229 3841
rect 3913 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4229 3840
rect 3913 3775 4229 3776
rect 9847 3840 10163 3841
rect 9847 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10163 3840
rect 9847 3775 10163 3776
rect 15781 3840 16097 3841
rect 15781 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16097 3840
rect 15781 3775 16097 3776
rect 21715 3840 22031 3841
rect 21715 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22031 3840
rect 21715 3775 22031 3776
rect 6880 3296 7196 3297
rect 6880 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7196 3296
rect 6880 3231 7196 3232
rect 12814 3296 13130 3297
rect 12814 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13130 3296
rect 12814 3231 13130 3232
rect 18748 3296 19064 3297
rect 18748 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19064 3296
rect 18748 3231 19064 3232
rect 24682 3296 24998 3297
rect 24682 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 24998 3296
rect 24682 3231 24998 3232
rect 8201 3090 8267 3093
rect 19190 3090 19196 3092
rect 8201 3088 19196 3090
rect 8201 3032 8206 3088
rect 8262 3032 19196 3088
rect 8201 3030 19196 3032
rect 8201 3027 8267 3030
rect 19190 3028 19196 3030
rect 19260 3028 19266 3092
rect 5390 2892 5396 2956
rect 5460 2954 5466 2956
rect 20662 2954 20668 2956
rect 5460 2894 20668 2954
rect 5460 2892 5466 2894
rect 20662 2892 20668 2894
rect 20732 2892 20738 2956
rect 3913 2752 4229 2753
rect 3913 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4229 2752
rect 3913 2687 4229 2688
rect 9847 2752 10163 2753
rect 9847 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10163 2752
rect 9847 2687 10163 2688
rect 15781 2752 16097 2753
rect 15781 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16097 2752
rect 15781 2687 16097 2688
rect 21715 2752 22031 2753
rect 21715 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22031 2752
rect 21715 2687 22031 2688
rect 14365 2682 14431 2685
rect 10366 2680 14431 2682
rect 10366 2624 14370 2680
rect 14426 2624 14431 2680
rect 10366 2622 14431 2624
rect 1577 2546 1643 2549
rect 10366 2546 10426 2622
rect 14365 2619 14431 2622
rect 1577 2544 10426 2546
rect 1577 2488 1582 2544
rect 1638 2488 10426 2544
rect 1577 2486 10426 2488
rect 12249 2546 12315 2549
rect 18137 2546 18203 2549
rect 12249 2544 18203 2546
rect 12249 2488 12254 2544
rect 12310 2488 18142 2544
rect 18198 2488 18203 2544
rect 12249 2486 18203 2488
rect 1577 2483 1643 2486
rect 12249 2483 12315 2486
rect 18137 2483 18203 2486
rect 6269 2410 6335 2413
rect 12198 2410 12204 2412
rect 6269 2408 12204 2410
rect 6269 2352 6274 2408
rect 6330 2352 12204 2408
rect 6269 2350 12204 2352
rect 6269 2347 6335 2350
rect 12198 2348 12204 2350
rect 12268 2348 12274 2412
rect 12566 2348 12572 2412
rect 12636 2410 12642 2412
rect 19701 2410 19767 2413
rect 12636 2408 19767 2410
rect 12636 2352 19706 2408
rect 19762 2352 19767 2408
rect 12636 2350 19767 2352
rect 12636 2348 12642 2350
rect 19701 2347 19767 2350
rect 8109 2274 8175 2277
rect 12249 2274 12315 2277
rect 8109 2272 12315 2274
rect 8109 2216 8114 2272
rect 8170 2216 12254 2272
rect 12310 2216 12315 2272
rect 8109 2214 12315 2216
rect 8109 2211 8175 2214
rect 12249 2211 12315 2214
rect 6880 2208 7196 2209
rect 6880 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7196 2208
rect 6880 2143 7196 2144
rect 12814 2208 13130 2209
rect 12814 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13130 2208
rect 12814 2143 13130 2144
rect 18748 2208 19064 2209
rect 18748 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19064 2208
rect 18748 2143 19064 2144
rect 24682 2208 24998 2209
rect 24682 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 24998 2208
rect 24682 2143 24998 2144
rect 7557 2138 7623 2141
rect 7557 2136 12450 2138
rect 7557 2080 7562 2136
rect 7618 2080 12450 2136
rect 7557 2078 12450 2080
rect 7557 2075 7623 2078
rect 6913 2002 6979 2005
rect 10225 2002 10291 2005
rect 6913 2000 10291 2002
rect 6913 1944 6918 2000
rect 6974 1944 10230 2000
rect 10286 1944 10291 2000
rect 6913 1942 10291 1944
rect 6913 1939 6979 1942
rect 10225 1939 10291 1942
rect 11094 1940 11100 2004
rect 11164 2002 11170 2004
rect 11789 2002 11855 2005
rect 11164 2000 11855 2002
rect 11164 1944 11794 2000
rect 11850 1944 11855 2000
rect 11164 1942 11855 1944
rect 12390 2002 12450 2078
rect 20253 2002 20319 2005
rect 12390 2000 20319 2002
rect 12390 1944 20258 2000
rect 20314 1944 20319 2000
rect 12390 1942 20319 1944
rect 11164 1940 11170 1942
rect 11789 1939 11855 1942
rect 20253 1939 20319 1942
rect 1485 1866 1551 1869
rect 20897 1866 20963 1869
rect 1485 1864 20963 1866
rect 1485 1808 1490 1864
rect 1546 1808 20902 1864
rect 20958 1808 20963 1864
rect 1485 1806 20963 1808
rect 1485 1803 1551 1806
rect 20897 1803 20963 1806
rect 7925 1730 7991 1733
rect 9213 1730 9279 1733
rect 7925 1728 9279 1730
rect 7925 1672 7930 1728
rect 7986 1672 9218 1728
rect 9274 1672 9279 1728
rect 7925 1670 9279 1672
rect 7925 1667 7991 1670
rect 9213 1667 9279 1670
rect 10225 1730 10291 1733
rect 10225 1728 15578 1730
rect 10225 1672 10230 1728
rect 10286 1672 15578 1728
rect 10225 1670 15578 1672
rect 10225 1667 10291 1670
rect 3913 1664 4229 1665
rect 3913 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4229 1664
rect 3913 1599 4229 1600
rect 9847 1664 10163 1665
rect 9847 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10163 1664
rect 9847 1599 10163 1600
rect 3049 1594 3115 1597
rect 3601 1594 3667 1597
rect 3049 1592 3667 1594
rect 3049 1536 3054 1592
rect 3110 1536 3606 1592
rect 3662 1536 3667 1592
rect 3049 1534 3667 1536
rect 3049 1531 3115 1534
rect 3601 1531 3667 1534
rect 8477 1594 8543 1597
rect 8937 1594 9003 1597
rect 8477 1592 9003 1594
rect 8477 1536 8482 1592
rect 8538 1536 8942 1592
rect 8998 1536 9003 1592
rect 8477 1534 9003 1536
rect 8477 1531 8543 1534
rect 8937 1531 9003 1534
rect 2221 1458 2287 1461
rect 14365 1458 14431 1461
rect 2221 1456 14431 1458
rect 2221 1400 2226 1456
rect 2282 1400 14370 1456
rect 14426 1400 14431 1456
rect 2221 1398 14431 1400
rect 15518 1458 15578 1670
rect 15781 1664 16097 1665
rect 15781 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16097 1664
rect 15781 1599 16097 1600
rect 21715 1664 22031 1665
rect 21715 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22031 1664
rect 21715 1599 22031 1600
rect 18505 1458 18571 1461
rect 15518 1456 18571 1458
rect 15518 1400 18510 1456
rect 18566 1400 18571 1456
rect 15518 1398 18571 1400
rect 2221 1395 2287 1398
rect 14365 1395 14431 1398
rect 18505 1395 18571 1398
rect 20161 1458 20227 1461
rect 21817 1458 21883 1461
rect 20161 1456 21883 1458
rect 20161 1400 20166 1456
rect 20222 1400 21822 1456
rect 21878 1400 21883 1456
rect 20161 1398 21883 1400
rect 20161 1395 20227 1398
rect 21817 1395 21883 1398
rect 2313 1322 2379 1325
rect 4797 1322 4863 1325
rect 5390 1322 5396 1324
rect 2313 1320 2790 1322
rect 2313 1264 2318 1320
rect 2374 1264 2790 1320
rect 2313 1262 2790 1264
rect 2313 1259 2379 1262
rect 2730 1186 2790 1262
rect 4797 1320 5396 1322
rect 4797 1264 4802 1320
rect 4858 1264 5396 1320
rect 4797 1262 5396 1264
rect 4797 1259 4863 1262
rect 5390 1260 5396 1262
rect 5460 1260 5466 1324
rect 11697 1322 11763 1325
rect 12709 1322 12775 1325
rect 5582 1320 11763 1322
rect 5582 1264 11702 1320
rect 11758 1264 11763 1320
rect 5582 1262 11763 1264
rect 5582 1186 5642 1262
rect 11697 1259 11763 1262
rect 12390 1320 12775 1322
rect 12390 1264 12714 1320
rect 12770 1264 12775 1320
rect 12390 1262 12775 1264
rect 2730 1126 5642 1186
rect 8201 1186 8267 1189
rect 8937 1186 9003 1189
rect 8201 1184 9003 1186
rect 8201 1128 8206 1184
rect 8262 1128 8942 1184
rect 8998 1128 9003 1184
rect 8201 1126 9003 1128
rect 8201 1123 8267 1126
rect 8937 1123 9003 1126
rect 6880 1120 7196 1121
rect 6880 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7196 1120
rect 6880 1055 7196 1056
rect 1669 1050 1735 1053
rect 2630 1050 2636 1052
rect 1669 1048 2636 1050
rect 1669 992 1674 1048
rect 1730 992 2636 1048
rect 1669 990 2636 992
rect 1669 987 1735 990
rect 2630 988 2636 990
rect 2700 988 2706 1052
rect 2957 1050 3023 1053
rect 8569 1050 8635 1053
rect 10317 1050 10383 1053
rect 2957 1048 6746 1050
rect 2957 992 2962 1048
rect 3018 992 6746 1048
rect 2957 990 6746 992
rect 2957 987 3023 990
rect 6686 914 6746 990
rect 8569 1048 10383 1050
rect 8569 992 8574 1048
rect 8630 992 10322 1048
rect 10378 992 10383 1048
rect 8569 990 10383 992
rect 8569 987 8635 990
rect 10317 987 10383 990
rect 12390 914 12450 1262
rect 12709 1259 12775 1262
rect 20662 1260 20668 1324
rect 20732 1322 20738 1324
rect 21725 1322 21791 1325
rect 20732 1320 21791 1322
rect 20732 1264 21730 1320
rect 21786 1264 21791 1320
rect 20732 1262 21791 1264
rect 20732 1260 20738 1262
rect 21725 1259 21791 1262
rect 22134 1260 22140 1324
rect 22204 1322 22210 1324
rect 22645 1322 22711 1325
rect 22204 1320 22711 1322
rect 22204 1264 22650 1320
rect 22706 1264 22711 1320
rect 22204 1262 22711 1264
rect 22204 1260 22210 1262
rect 22645 1259 22711 1262
rect 19190 1124 19196 1188
rect 19260 1186 19266 1188
rect 21449 1186 21515 1189
rect 19260 1184 21515 1186
rect 19260 1128 21454 1184
rect 21510 1128 21515 1184
rect 19260 1126 21515 1128
rect 19260 1124 19266 1126
rect 21449 1123 21515 1126
rect 22737 1186 22803 1189
rect 24025 1186 24091 1189
rect 22737 1184 24091 1186
rect 22737 1128 22742 1184
rect 22798 1128 24030 1184
rect 24086 1128 24091 1184
rect 22737 1126 24091 1128
rect 22737 1123 22803 1126
rect 24025 1123 24091 1126
rect 12814 1120 13130 1121
rect 12814 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13130 1120
rect 12814 1055 13130 1056
rect 18748 1120 19064 1121
rect 18748 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19064 1120
rect 18748 1055 19064 1056
rect 24682 1120 24998 1121
rect 24682 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 24998 1120
rect 24682 1055 24998 1056
rect 22369 1050 22435 1053
rect 23841 1050 23907 1053
rect 22369 1048 23907 1050
rect 22369 992 22374 1048
rect 22430 992 23846 1048
rect 23902 992 23907 1048
rect 22369 990 23907 992
rect 22369 987 22435 990
rect 23841 987 23907 990
rect 6686 854 12450 914
rect 7557 778 7623 781
rect 11329 778 11395 781
rect 7557 776 11395 778
rect 7557 720 7562 776
rect 7618 720 11334 776
rect 11390 720 11395 776
rect 7557 718 11395 720
rect 7557 715 7623 718
rect 11329 715 11395 718
rect 6913 642 6979 645
rect 10593 642 10659 645
rect 6913 640 10659 642
rect 6913 584 6918 640
rect 6974 584 10598 640
rect 10654 584 10659 640
rect 6913 582 10659 584
rect 6913 579 6979 582
rect 10593 579 10659 582
<< via3 >>
rect 6886 6556 6950 6560
rect 6886 6500 6890 6556
rect 6890 6500 6946 6556
rect 6946 6500 6950 6556
rect 6886 6496 6950 6500
rect 6966 6556 7030 6560
rect 6966 6500 6970 6556
rect 6970 6500 7026 6556
rect 7026 6500 7030 6556
rect 6966 6496 7030 6500
rect 7046 6556 7110 6560
rect 7046 6500 7050 6556
rect 7050 6500 7106 6556
rect 7106 6500 7110 6556
rect 7046 6496 7110 6500
rect 7126 6556 7190 6560
rect 7126 6500 7130 6556
rect 7130 6500 7186 6556
rect 7186 6500 7190 6556
rect 7126 6496 7190 6500
rect 12820 6556 12884 6560
rect 12820 6500 12824 6556
rect 12824 6500 12880 6556
rect 12880 6500 12884 6556
rect 12820 6496 12884 6500
rect 12900 6556 12964 6560
rect 12900 6500 12904 6556
rect 12904 6500 12960 6556
rect 12960 6500 12964 6556
rect 12900 6496 12964 6500
rect 12980 6556 13044 6560
rect 12980 6500 12984 6556
rect 12984 6500 13040 6556
rect 13040 6500 13044 6556
rect 12980 6496 13044 6500
rect 13060 6556 13124 6560
rect 13060 6500 13064 6556
rect 13064 6500 13120 6556
rect 13120 6500 13124 6556
rect 13060 6496 13124 6500
rect 18754 6556 18818 6560
rect 18754 6500 18758 6556
rect 18758 6500 18814 6556
rect 18814 6500 18818 6556
rect 18754 6496 18818 6500
rect 18834 6556 18898 6560
rect 18834 6500 18838 6556
rect 18838 6500 18894 6556
rect 18894 6500 18898 6556
rect 18834 6496 18898 6500
rect 18914 6556 18978 6560
rect 18914 6500 18918 6556
rect 18918 6500 18974 6556
rect 18974 6500 18978 6556
rect 18914 6496 18978 6500
rect 18994 6556 19058 6560
rect 18994 6500 18998 6556
rect 18998 6500 19054 6556
rect 19054 6500 19058 6556
rect 18994 6496 19058 6500
rect 24688 6556 24752 6560
rect 24688 6500 24692 6556
rect 24692 6500 24748 6556
rect 24748 6500 24752 6556
rect 24688 6496 24752 6500
rect 24768 6556 24832 6560
rect 24768 6500 24772 6556
rect 24772 6500 24828 6556
rect 24828 6500 24832 6556
rect 24768 6496 24832 6500
rect 24848 6556 24912 6560
rect 24848 6500 24852 6556
rect 24852 6500 24908 6556
rect 24908 6500 24912 6556
rect 24848 6496 24912 6500
rect 24928 6556 24992 6560
rect 24928 6500 24932 6556
rect 24932 6500 24988 6556
rect 24988 6500 24992 6556
rect 24928 6496 24992 6500
rect 3919 6012 3983 6016
rect 3919 5956 3923 6012
rect 3923 5956 3979 6012
rect 3979 5956 3983 6012
rect 3919 5952 3983 5956
rect 3999 6012 4063 6016
rect 3999 5956 4003 6012
rect 4003 5956 4059 6012
rect 4059 5956 4063 6012
rect 3999 5952 4063 5956
rect 4079 6012 4143 6016
rect 4079 5956 4083 6012
rect 4083 5956 4139 6012
rect 4139 5956 4143 6012
rect 4079 5952 4143 5956
rect 4159 6012 4223 6016
rect 4159 5956 4163 6012
rect 4163 5956 4219 6012
rect 4219 5956 4223 6012
rect 4159 5952 4223 5956
rect 9853 6012 9917 6016
rect 9853 5956 9857 6012
rect 9857 5956 9913 6012
rect 9913 5956 9917 6012
rect 9853 5952 9917 5956
rect 9933 6012 9997 6016
rect 9933 5956 9937 6012
rect 9937 5956 9993 6012
rect 9993 5956 9997 6012
rect 9933 5952 9997 5956
rect 10013 6012 10077 6016
rect 10013 5956 10017 6012
rect 10017 5956 10073 6012
rect 10073 5956 10077 6012
rect 10013 5952 10077 5956
rect 10093 6012 10157 6016
rect 10093 5956 10097 6012
rect 10097 5956 10153 6012
rect 10153 5956 10157 6012
rect 10093 5952 10157 5956
rect 15787 6012 15851 6016
rect 15787 5956 15791 6012
rect 15791 5956 15847 6012
rect 15847 5956 15851 6012
rect 15787 5952 15851 5956
rect 15867 6012 15931 6016
rect 15867 5956 15871 6012
rect 15871 5956 15927 6012
rect 15927 5956 15931 6012
rect 15867 5952 15931 5956
rect 15947 6012 16011 6016
rect 15947 5956 15951 6012
rect 15951 5956 16007 6012
rect 16007 5956 16011 6012
rect 15947 5952 16011 5956
rect 16027 6012 16091 6016
rect 16027 5956 16031 6012
rect 16031 5956 16087 6012
rect 16087 5956 16091 6012
rect 16027 5952 16091 5956
rect 21721 6012 21785 6016
rect 21721 5956 21725 6012
rect 21725 5956 21781 6012
rect 21781 5956 21785 6012
rect 21721 5952 21785 5956
rect 21801 6012 21865 6016
rect 21801 5956 21805 6012
rect 21805 5956 21861 6012
rect 21861 5956 21865 6012
rect 21801 5952 21865 5956
rect 21881 6012 21945 6016
rect 21881 5956 21885 6012
rect 21885 5956 21941 6012
rect 21941 5956 21945 6012
rect 21881 5952 21945 5956
rect 21961 6012 22025 6016
rect 21961 5956 21965 6012
rect 21965 5956 22021 6012
rect 22021 5956 22025 6012
rect 21961 5952 22025 5956
rect 6886 5468 6950 5472
rect 6886 5412 6890 5468
rect 6890 5412 6946 5468
rect 6946 5412 6950 5468
rect 6886 5408 6950 5412
rect 6966 5468 7030 5472
rect 6966 5412 6970 5468
rect 6970 5412 7026 5468
rect 7026 5412 7030 5468
rect 6966 5408 7030 5412
rect 7046 5468 7110 5472
rect 7046 5412 7050 5468
rect 7050 5412 7106 5468
rect 7106 5412 7110 5468
rect 7046 5408 7110 5412
rect 7126 5468 7190 5472
rect 7126 5412 7130 5468
rect 7130 5412 7186 5468
rect 7186 5412 7190 5468
rect 7126 5408 7190 5412
rect 12820 5468 12884 5472
rect 12820 5412 12824 5468
rect 12824 5412 12880 5468
rect 12880 5412 12884 5468
rect 12820 5408 12884 5412
rect 12900 5468 12964 5472
rect 12900 5412 12904 5468
rect 12904 5412 12960 5468
rect 12960 5412 12964 5468
rect 12900 5408 12964 5412
rect 12980 5468 13044 5472
rect 12980 5412 12984 5468
rect 12984 5412 13040 5468
rect 13040 5412 13044 5468
rect 12980 5408 13044 5412
rect 13060 5468 13124 5472
rect 13060 5412 13064 5468
rect 13064 5412 13120 5468
rect 13120 5412 13124 5468
rect 13060 5408 13124 5412
rect 18754 5468 18818 5472
rect 18754 5412 18758 5468
rect 18758 5412 18814 5468
rect 18814 5412 18818 5468
rect 18754 5408 18818 5412
rect 18834 5468 18898 5472
rect 18834 5412 18838 5468
rect 18838 5412 18894 5468
rect 18894 5412 18898 5468
rect 18834 5408 18898 5412
rect 18914 5468 18978 5472
rect 18914 5412 18918 5468
rect 18918 5412 18974 5468
rect 18974 5412 18978 5468
rect 18914 5408 18978 5412
rect 18994 5468 19058 5472
rect 18994 5412 18998 5468
rect 18998 5412 19054 5468
rect 19054 5412 19058 5468
rect 18994 5408 19058 5412
rect 24688 5468 24752 5472
rect 24688 5412 24692 5468
rect 24692 5412 24748 5468
rect 24748 5412 24752 5468
rect 24688 5408 24752 5412
rect 24768 5468 24832 5472
rect 24768 5412 24772 5468
rect 24772 5412 24828 5468
rect 24828 5412 24832 5468
rect 24768 5408 24832 5412
rect 24848 5468 24912 5472
rect 24848 5412 24852 5468
rect 24852 5412 24908 5468
rect 24908 5412 24912 5468
rect 24848 5408 24912 5412
rect 24928 5468 24992 5472
rect 24928 5412 24932 5468
rect 24932 5412 24988 5468
rect 24988 5412 24992 5468
rect 24928 5408 24992 5412
rect 3919 4924 3983 4928
rect 3919 4868 3923 4924
rect 3923 4868 3979 4924
rect 3979 4868 3983 4924
rect 3919 4864 3983 4868
rect 3999 4924 4063 4928
rect 3999 4868 4003 4924
rect 4003 4868 4059 4924
rect 4059 4868 4063 4924
rect 3999 4864 4063 4868
rect 4079 4924 4143 4928
rect 4079 4868 4083 4924
rect 4083 4868 4139 4924
rect 4139 4868 4143 4924
rect 4079 4864 4143 4868
rect 4159 4924 4223 4928
rect 4159 4868 4163 4924
rect 4163 4868 4219 4924
rect 4219 4868 4223 4924
rect 4159 4864 4223 4868
rect 9853 4924 9917 4928
rect 9853 4868 9857 4924
rect 9857 4868 9913 4924
rect 9913 4868 9917 4924
rect 9853 4864 9917 4868
rect 9933 4924 9997 4928
rect 9933 4868 9937 4924
rect 9937 4868 9993 4924
rect 9993 4868 9997 4924
rect 9933 4864 9997 4868
rect 10013 4924 10077 4928
rect 10013 4868 10017 4924
rect 10017 4868 10073 4924
rect 10073 4868 10077 4924
rect 10013 4864 10077 4868
rect 10093 4924 10157 4928
rect 10093 4868 10097 4924
rect 10097 4868 10153 4924
rect 10153 4868 10157 4924
rect 10093 4864 10157 4868
rect 15787 4924 15851 4928
rect 15787 4868 15791 4924
rect 15791 4868 15847 4924
rect 15847 4868 15851 4924
rect 15787 4864 15851 4868
rect 15867 4924 15931 4928
rect 15867 4868 15871 4924
rect 15871 4868 15927 4924
rect 15927 4868 15931 4924
rect 15867 4864 15931 4868
rect 15947 4924 16011 4928
rect 15947 4868 15951 4924
rect 15951 4868 16007 4924
rect 16007 4868 16011 4924
rect 15947 4864 16011 4868
rect 16027 4924 16091 4928
rect 16027 4868 16031 4924
rect 16031 4868 16087 4924
rect 16087 4868 16091 4924
rect 16027 4864 16091 4868
rect 21721 4924 21785 4928
rect 21721 4868 21725 4924
rect 21725 4868 21781 4924
rect 21781 4868 21785 4924
rect 21721 4864 21785 4868
rect 21801 4924 21865 4928
rect 21801 4868 21805 4924
rect 21805 4868 21861 4924
rect 21861 4868 21865 4924
rect 21801 4864 21865 4868
rect 21881 4924 21945 4928
rect 21881 4868 21885 4924
rect 21885 4868 21941 4924
rect 21941 4868 21945 4924
rect 21881 4864 21945 4868
rect 21961 4924 22025 4928
rect 21961 4868 21965 4924
rect 21965 4868 22021 4924
rect 22021 4868 22025 4924
rect 21961 4864 22025 4868
rect 6886 4380 6950 4384
rect 6886 4324 6890 4380
rect 6890 4324 6946 4380
rect 6946 4324 6950 4380
rect 6886 4320 6950 4324
rect 6966 4380 7030 4384
rect 6966 4324 6970 4380
rect 6970 4324 7026 4380
rect 7026 4324 7030 4380
rect 6966 4320 7030 4324
rect 7046 4380 7110 4384
rect 7046 4324 7050 4380
rect 7050 4324 7106 4380
rect 7106 4324 7110 4380
rect 7046 4320 7110 4324
rect 7126 4380 7190 4384
rect 7126 4324 7130 4380
rect 7130 4324 7186 4380
rect 7186 4324 7190 4380
rect 7126 4320 7190 4324
rect 12820 4380 12884 4384
rect 12820 4324 12824 4380
rect 12824 4324 12880 4380
rect 12880 4324 12884 4380
rect 12820 4320 12884 4324
rect 12900 4380 12964 4384
rect 12900 4324 12904 4380
rect 12904 4324 12960 4380
rect 12960 4324 12964 4380
rect 12900 4320 12964 4324
rect 12980 4380 13044 4384
rect 12980 4324 12984 4380
rect 12984 4324 13040 4380
rect 13040 4324 13044 4380
rect 12980 4320 13044 4324
rect 13060 4380 13124 4384
rect 13060 4324 13064 4380
rect 13064 4324 13120 4380
rect 13120 4324 13124 4380
rect 13060 4320 13124 4324
rect 18754 4380 18818 4384
rect 18754 4324 18758 4380
rect 18758 4324 18814 4380
rect 18814 4324 18818 4380
rect 18754 4320 18818 4324
rect 18834 4380 18898 4384
rect 18834 4324 18838 4380
rect 18838 4324 18894 4380
rect 18894 4324 18898 4380
rect 18834 4320 18898 4324
rect 18914 4380 18978 4384
rect 18914 4324 18918 4380
rect 18918 4324 18974 4380
rect 18974 4324 18978 4380
rect 18914 4320 18978 4324
rect 18994 4380 19058 4384
rect 18994 4324 18998 4380
rect 18998 4324 19054 4380
rect 19054 4324 19058 4380
rect 18994 4320 19058 4324
rect 24688 4380 24752 4384
rect 24688 4324 24692 4380
rect 24692 4324 24748 4380
rect 24748 4324 24752 4380
rect 24688 4320 24752 4324
rect 24768 4380 24832 4384
rect 24768 4324 24772 4380
rect 24772 4324 24828 4380
rect 24828 4324 24832 4380
rect 24768 4320 24832 4324
rect 24848 4380 24912 4384
rect 24848 4324 24852 4380
rect 24852 4324 24908 4380
rect 24908 4324 24912 4380
rect 24848 4320 24912 4324
rect 24928 4380 24992 4384
rect 24928 4324 24932 4380
rect 24932 4324 24988 4380
rect 24988 4324 24992 4380
rect 24928 4320 24992 4324
rect 22140 4116 22204 4180
rect 3919 3836 3983 3840
rect 3919 3780 3923 3836
rect 3923 3780 3979 3836
rect 3979 3780 3983 3836
rect 3919 3776 3983 3780
rect 3999 3836 4063 3840
rect 3999 3780 4003 3836
rect 4003 3780 4059 3836
rect 4059 3780 4063 3836
rect 3999 3776 4063 3780
rect 4079 3836 4143 3840
rect 4079 3780 4083 3836
rect 4083 3780 4139 3836
rect 4139 3780 4143 3836
rect 4079 3776 4143 3780
rect 4159 3836 4223 3840
rect 4159 3780 4163 3836
rect 4163 3780 4219 3836
rect 4219 3780 4223 3836
rect 4159 3776 4223 3780
rect 9853 3836 9917 3840
rect 9853 3780 9857 3836
rect 9857 3780 9913 3836
rect 9913 3780 9917 3836
rect 9853 3776 9917 3780
rect 9933 3836 9997 3840
rect 9933 3780 9937 3836
rect 9937 3780 9993 3836
rect 9993 3780 9997 3836
rect 9933 3776 9997 3780
rect 10013 3836 10077 3840
rect 10013 3780 10017 3836
rect 10017 3780 10073 3836
rect 10073 3780 10077 3836
rect 10013 3776 10077 3780
rect 10093 3836 10157 3840
rect 10093 3780 10097 3836
rect 10097 3780 10153 3836
rect 10153 3780 10157 3836
rect 10093 3776 10157 3780
rect 15787 3836 15851 3840
rect 15787 3780 15791 3836
rect 15791 3780 15847 3836
rect 15847 3780 15851 3836
rect 15787 3776 15851 3780
rect 15867 3836 15931 3840
rect 15867 3780 15871 3836
rect 15871 3780 15927 3836
rect 15927 3780 15931 3836
rect 15867 3776 15931 3780
rect 15947 3836 16011 3840
rect 15947 3780 15951 3836
rect 15951 3780 16007 3836
rect 16007 3780 16011 3836
rect 15947 3776 16011 3780
rect 16027 3836 16091 3840
rect 16027 3780 16031 3836
rect 16031 3780 16087 3836
rect 16087 3780 16091 3836
rect 16027 3776 16091 3780
rect 21721 3836 21785 3840
rect 21721 3780 21725 3836
rect 21725 3780 21781 3836
rect 21781 3780 21785 3836
rect 21721 3776 21785 3780
rect 21801 3836 21865 3840
rect 21801 3780 21805 3836
rect 21805 3780 21861 3836
rect 21861 3780 21865 3836
rect 21801 3776 21865 3780
rect 21881 3836 21945 3840
rect 21881 3780 21885 3836
rect 21885 3780 21941 3836
rect 21941 3780 21945 3836
rect 21881 3776 21945 3780
rect 21961 3836 22025 3840
rect 21961 3780 21965 3836
rect 21965 3780 22021 3836
rect 22021 3780 22025 3836
rect 21961 3776 22025 3780
rect 6886 3292 6950 3296
rect 6886 3236 6890 3292
rect 6890 3236 6946 3292
rect 6946 3236 6950 3292
rect 6886 3232 6950 3236
rect 6966 3292 7030 3296
rect 6966 3236 6970 3292
rect 6970 3236 7026 3292
rect 7026 3236 7030 3292
rect 6966 3232 7030 3236
rect 7046 3292 7110 3296
rect 7046 3236 7050 3292
rect 7050 3236 7106 3292
rect 7106 3236 7110 3292
rect 7046 3232 7110 3236
rect 7126 3292 7190 3296
rect 7126 3236 7130 3292
rect 7130 3236 7186 3292
rect 7186 3236 7190 3292
rect 7126 3232 7190 3236
rect 12820 3292 12884 3296
rect 12820 3236 12824 3292
rect 12824 3236 12880 3292
rect 12880 3236 12884 3292
rect 12820 3232 12884 3236
rect 12900 3292 12964 3296
rect 12900 3236 12904 3292
rect 12904 3236 12960 3292
rect 12960 3236 12964 3292
rect 12900 3232 12964 3236
rect 12980 3292 13044 3296
rect 12980 3236 12984 3292
rect 12984 3236 13040 3292
rect 13040 3236 13044 3292
rect 12980 3232 13044 3236
rect 13060 3292 13124 3296
rect 13060 3236 13064 3292
rect 13064 3236 13120 3292
rect 13120 3236 13124 3292
rect 13060 3232 13124 3236
rect 18754 3292 18818 3296
rect 18754 3236 18758 3292
rect 18758 3236 18814 3292
rect 18814 3236 18818 3292
rect 18754 3232 18818 3236
rect 18834 3292 18898 3296
rect 18834 3236 18838 3292
rect 18838 3236 18894 3292
rect 18894 3236 18898 3292
rect 18834 3232 18898 3236
rect 18914 3292 18978 3296
rect 18914 3236 18918 3292
rect 18918 3236 18974 3292
rect 18974 3236 18978 3292
rect 18914 3232 18978 3236
rect 18994 3292 19058 3296
rect 18994 3236 18998 3292
rect 18998 3236 19054 3292
rect 19054 3236 19058 3292
rect 18994 3232 19058 3236
rect 24688 3292 24752 3296
rect 24688 3236 24692 3292
rect 24692 3236 24748 3292
rect 24748 3236 24752 3292
rect 24688 3232 24752 3236
rect 24768 3292 24832 3296
rect 24768 3236 24772 3292
rect 24772 3236 24828 3292
rect 24828 3236 24832 3292
rect 24768 3232 24832 3236
rect 24848 3292 24912 3296
rect 24848 3236 24852 3292
rect 24852 3236 24908 3292
rect 24908 3236 24912 3292
rect 24848 3232 24912 3236
rect 24928 3292 24992 3296
rect 24928 3236 24932 3292
rect 24932 3236 24988 3292
rect 24988 3236 24992 3292
rect 24928 3232 24992 3236
rect 19196 3028 19260 3092
rect 5396 2892 5460 2956
rect 20668 2892 20732 2956
rect 3919 2748 3983 2752
rect 3919 2692 3923 2748
rect 3923 2692 3979 2748
rect 3979 2692 3983 2748
rect 3919 2688 3983 2692
rect 3999 2748 4063 2752
rect 3999 2692 4003 2748
rect 4003 2692 4059 2748
rect 4059 2692 4063 2748
rect 3999 2688 4063 2692
rect 4079 2748 4143 2752
rect 4079 2692 4083 2748
rect 4083 2692 4139 2748
rect 4139 2692 4143 2748
rect 4079 2688 4143 2692
rect 4159 2748 4223 2752
rect 4159 2692 4163 2748
rect 4163 2692 4219 2748
rect 4219 2692 4223 2748
rect 4159 2688 4223 2692
rect 9853 2748 9917 2752
rect 9853 2692 9857 2748
rect 9857 2692 9913 2748
rect 9913 2692 9917 2748
rect 9853 2688 9917 2692
rect 9933 2748 9997 2752
rect 9933 2692 9937 2748
rect 9937 2692 9993 2748
rect 9993 2692 9997 2748
rect 9933 2688 9997 2692
rect 10013 2748 10077 2752
rect 10013 2692 10017 2748
rect 10017 2692 10073 2748
rect 10073 2692 10077 2748
rect 10013 2688 10077 2692
rect 10093 2748 10157 2752
rect 10093 2692 10097 2748
rect 10097 2692 10153 2748
rect 10153 2692 10157 2748
rect 10093 2688 10157 2692
rect 15787 2748 15851 2752
rect 15787 2692 15791 2748
rect 15791 2692 15847 2748
rect 15847 2692 15851 2748
rect 15787 2688 15851 2692
rect 15867 2748 15931 2752
rect 15867 2692 15871 2748
rect 15871 2692 15927 2748
rect 15927 2692 15931 2748
rect 15867 2688 15931 2692
rect 15947 2748 16011 2752
rect 15947 2692 15951 2748
rect 15951 2692 16007 2748
rect 16007 2692 16011 2748
rect 15947 2688 16011 2692
rect 16027 2748 16091 2752
rect 16027 2692 16031 2748
rect 16031 2692 16087 2748
rect 16087 2692 16091 2748
rect 16027 2688 16091 2692
rect 21721 2748 21785 2752
rect 21721 2692 21725 2748
rect 21725 2692 21781 2748
rect 21781 2692 21785 2748
rect 21721 2688 21785 2692
rect 21801 2748 21865 2752
rect 21801 2692 21805 2748
rect 21805 2692 21861 2748
rect 21861 2692 21865 2748
rect 21801 2688 21865 2692
rect 21881 2748 21945 2752
rect 21881 2692 21885 2748
rect 21885 2692 21941 2748
rect 21941 2692 21945 2748
rect 21881 2688 21945 2692
rect 21961 2748 22025 2752
rect 21961 2692 21965 2748
rect 21965 2692 22021 2748
rect 22021 2692 22025 2748
rect 21961 2688 22025 2692
rect 12204 2348 12268 2412
rect 12572 2348 12636 2412
rect 6886 2204 6950 2208
rect 6886 2148 6890 2204
rect 6890 2148 6946 2204
rect 6946 2148 6950 2204
rect 6886 2144 6950 2148
rect 6966 2204 7030 2208
rect 6966 2148 6970 2204
rect 6970 2148 7026 2204
rect 7026 2148 7030 2204
rect 6966 2144 7030 2148
rect 7046 2204 7110 2208
rect 7046 2148 7050 2204
rect 7050 2148 7106 2204
rect 7106 2148 7110 2204
rect 7046 2144 7110 2148
rect 7126 2204 7190 2208
rect 7126 2148 7130 2204
rect 7130 2148 7186 2204
rect 7186 2148 7190 2204
rect 7126 2144 7190 2148
rect 12820 2204 12884 2208
rect 12820 2148 12824 2204
rect 12824 2148 12880 2204
rect 12880 2148 12884 2204
rect 12820 2144 12884 2148
rect 12900 2204 12964 2208
rect 12900 2148 12904 2204
rect 12904 2148 12960 2204
rect 12960 2148 12964 2204
rect 12900 2144 12964 2148
rect 12980 2204 13044 2208
rect 12980 2148 12984 2204
rect 12984 2148 13040 2204
rect 13040 2148 13044 2204
rect 12980 2144 13044 2148
rect 13060 2204 13124 2208
rect 13060 2148 13064 2204
rect 13064 2148 13120 2204
rect 13120 2148 13124 2204
rect 13060 2144 13124 2148
rect 18754 2204 18818 2208
rect 18754 2148 18758 2204
rect 18758 2148 18814 2204
rect 18814 2148 18818 2204
rect 18754 2144 18818 2148
rect 18834 2204 18898 2208
rect 18834 2148 18838 2204
rect 18838 2148 18894 2204
rect 18894 2148 18898 2204
rect 18834 2144 18898 2148
rect 18914 2204 18978 2208
rect 18914 2148 18918 2204
rect 18918 2148 18974 2204
rect 18974 2148 18978 2204
rect 18914 2144 18978 2148
rect 18994 2204 19058 2208
rect 18994 2148 18998 2204
rect 18998 2148 19054 2204
rect 19054 2148 19058 2204
rect 18994 2144 19058 2148
rect 24688 2204 24752 2208
rect 24688 2148 24692 2204
rect 24692 2148 24748 2204
rect 24748 2148 24752 2204
rect 24688 2144 24752 2148
rect 24768 2204 24832 2208
rect 24768 2148 24772 2204
rect 24772 2148 24828 2204
rect 24828 2148 24832 2204
rect 24768 2144 24832 2148
rect 24848 2204 24912 2208
rect 24848 2148 24852 2204
rect 24852 2148 24908 2204
rect 24908 2148 24912 2204
rect 24848 2144 24912 2148
rect 24928 2204 24992 2208
rect 24928 2148 24932 2204
rect 24932 2148 24988 2204
rect 24988 2148 24992 2204
rect 24928 2144 24992 2148
rect 11100 1940 11164 2004
rect 3919 1660 3983 1664
rect 3919 1604 3923 1660
rect 3923 1604 3979 1660
rect 3979 1604 3983 1660
rect 3919 1600 3983 1604
rect 3999 1660 4063 1664
rect 3999 1604 4003 1660
rect 4003 1604 4059 1660
rect 4059 1604 4063 1660
rect 3999 1600 4063 1604
rect 4079 1660 4143 1664
rect 4079 1604 4083 1660
rect 4083 1604 4139 1660
rect 4139 1604 4143 1660
rect 4079 1600 4143 1604
rect 4159 1660 4223 1664
rect 4159 1604 4163 1660
rect 4163 1604 4219 1660
rect 4219 1604 4223 1660
rect 4159 1600 4223 1604
rect 9853 1660 9917 1664
rect 9853 1604 9857 1660
rect 9857 1604 9913 1660
rect 9913 1604 9917 1660
rect 9853 1600 9917 1604
rect 9933 1660 9997 1664
rect 9933 1604 9937 1660
rect 9937 1604 9993 1660
rect 9993 1604 9997 1660
rect 9933 1600 9997 1604
rect 10013 1660 10077 1664
rect 10013 1604 10017 1660
rect 10017 1604 10073 1660
rect 10073 1604 10077 1660
rect 10013 1600 10077 1604
rect 10093 1660 10157 1664
rect 10093 1604 10097 1660
rect 10097 1604 10153 1660
rect 10153 1604 10157 1660
rect 10093 1600 10157 1604
rect 15787 1660 15851 1664
rect 15787 1604 15791 1660
rect 15791 1604 15847 1660
rect 15847 1604 15851 1660
rect 15787 1600 15851 1604
rect 15867 1660 15931 1664
rect 15867 1604 15871 1660
rect 15871 1604 15927 1660
rect 15927 1604 15931 1660
rect 15867 1600 15931 1604
rect 15947 1660 16011 1664
rect 15947 1604 15951 1660
rect 15951 1604 16007 1660
rect 16007 1604 16011 1660
rect 15947 1600 16011 1604
rect 16027 1660 16091 1664
rect 16027 1604 16031 1660
rect 16031 1604 16087 1660
rect 16087 1604 16091 1660
rect 16027 1600 16091 1604
rect 21721 1660 21785 1664
rect 21721 1604 21725 1660
rect 21725 1604 21781 1660
rect 21781 1604 21785 1660
rect 21721 1600 21785 1604
rect 21801 1660 21865 1664
rect 21801 1604 21805 1660
rect 21805 1604 21861 1660
rect 21861 1604 21865 1660
rect 21801 1600 21865 1604
rect 21881 1660 21945 1664
rect 21881 1604 21885 1660
rect 21885 1604 21941 1660
rect 21941 1604 21945 1660
rect 21881 1600 21945 1604
rect 21961 1660 22025 1664
rect 21961 1604 21965 1660
rect 21965 1604 22021 1660
rect 22021 1604 22025 1660
rect 21961 1600 22025 1604
rect 5396 1260 5460 1324
rect 6886 1116 6950 1120
rect 6886 1060 6890 1116
rect 6890 1060 6946 1116
rect 6946 1060 6950 1116
rect 6886 1056 6950 1060
rect 6966 1116 7030 1120
rect 6966 1060 6970 1116
rect 6970 1060 7026 1116
rect 7026 1060 7030 1116
rect 6966 1056 7030 1060
rect 7046 1116 7110 1120
rect 7046 1060 7050 1116
rect 7050 1060 7106 1116
rect 7106 1060 7110 1116
rect 7046 1056 7110 1060
rect 7126 1116 7190 1120
rect 7126 1060 7130 1116
rect 7130 1060 7186 1116
rect 7186 1060 7190 1116
rect 7126 1056 7190 1060
rect 2636 988 2700 1052
rect 20668 1260 20732 1324
rect 22140 1260 22204 1324
rect 19196 1124 19260 1188
rect 12820 1116 12884 1120
rect 12820 1060 12824 1116
rect 12824 1060 12880 1116
rect 12880 1060 12884 1116
rect 12820 1056 12884 1060
rect 12900 1116 12964 1120
rect 12900 1060 12904 1116
rect 12904 1060 12960 1116
rect 12960 1060 12964 1116
rect 12900 1056 12964 1060
rect 12980 1116 13044 1120
rect 12980 1060 12984 1116
rect 12984 1060 13040 1116
rect 13040 1060 13044 1116
rect 12980 1056 13044 1060
rect 13060 1116 13124 1120
rect 13060 1060 13064 1116
rect 13064 1060 13120 1116
rect 13120 1060 13124 1116
rect 13060 1056 13124 1060
rect 18754 1116 18818 1120
rect 18754 1060 18758 1116
rect 18758 1060 18814 1116
rect 18814 1060 18818 1116
rect 18754 1056 18818 1060
rect 18834 1116 18898 1120
rect 18834 1060 18838 1116
rect 18838 1060 18894 1116
rect 18894 1060 18898 1116
rect 18834 1056 18898 1060
rect 18914 1116 18978 1120
rect 18914 1060 18918 1116
rect 18918 1060 18974 1116
rect 18974 1060 18978 1116
rect 18914 1056 18978 1060
rect 18994 1116 19058 1120
rect 18994 1060 18998 1116
rect 18998 1060 19054 1116
rect 19054 1060 19058 1116
rect 18994 1056 19058 1060
rect 24688 1116 24752 1120
rect 24688 1060 24692 1116
rect 24692 1060 24748 1116
rect 24748 1060 24752 1116
rect 24688 1056 24752 1060
rect 24768 1116 24832 1120
rect 24768 1060 24772 1116
rect 24772 1060 24828 1116
rect 24828 1060 24832 1116
rect 24768 1056 24832 1060
rect 24848 1116 24912 1120
rect 24848 1060 24852 1116
rect 24852 1060 24908 1116
rect 24908 1060 24912 1116
rect 24848 1056 24912 1060
rect 24928 1116 24992 1120
rect 24928 1060 24932 1116
rect 24932 1060 24988 1116
rect 24988 1060 24992 1116
rect 24928 1056 24992 1060
<< metal4 >>
rect 3911 6016 4231 6576
rect 3911 5952 3919 6016
rect 3983 5952 3999 6016
rect 4063 5952 4079 6016
rect 4143 5952 4159 6016
rect 4223 5952 4231 6016
rect 3911 4928 4231 5952
rect 3911 4864 3919 4928
rect 3983 4864 3999 4928
rect 4063 4864 4079 4928
rect 4143 4864 4159 4928
rect 4223 4864 4231 4928
rect 3911 3840 4231 4864
rect 3911 3776 3919 3840
rect 3983 3776 3999 3840
rect 4063 3776 4079 3840
rect 4143 3776 4159 3840
rect 4223 3776 4231 3840
rect 3911 2752 4231 3776
rect 6878 6560 7198 6576
rect 6878 6496 6886 6560
rect 6950 6496 6966 6560
rect 7030 6496 7046 6560
rect 7110 6496 7126 6560
rect 7190 6496 7198 6560
rect 6878 5472 7198 6496
rect 6878 5408 6886 5472
rect 6950 5408 6966 5472
rect 7030 5408 7046 5472
rect 7110 5408 7126 5472
rect 7190 5408 7198 5472
rect 6878 4384 7198 5408
rect 6878 4320 6886 4384
rect 6950 4320 6966 4384
rect 7030 4320 7046 4384
rect 7110 4320 7126 4384
rect 7190 4320 7198 4384
rect 6878 3296 7198 4320
rect 6878 3232 6886 3296
rect 6950 3232 6966 3296
rect 7030 3232 7046 3296
rect 7110 3232 7126 3296
rect 7190 3232 7198 3296
rect 5395 2956 5461 2957
rect 5395 2892 5396 2956
rect 5460 2892 5461 2956
rect 5395 2891 5461 2892
rect 3911 2688 3919 2752
rect 3983 2688 3999 2752
rect 4063 2688 4079 2752
rect 4143 2688 4159 2752
rect 4223 2688 4231 2752
rect 3911 1664 4231 2688
rect 3911 1600 3919 1664
rect 3983 1600 3999 1664
rect 4063 1600 4079 1664
rect 4143 1600 4159 1664
rect 4223 1600 4231 1664
rect 3911 1040 4231 1600
rect 5398 1325 5458 2891
rect 6878 2208 7198 3232
rect 6878 2144 6886 2208
rect 6950 2144 6966 2208
rect 7030 2144 7046 2208
rect 7110 2144 7126 2208
rect 7190 2144 7198 2208
rect 5395 1324 5461 1325
rect 5395 1260 5396 1324
rect 5460 1260 5461 1324
rect 5395 1259 5461 1260
rect 6878 1120 7198 2144
rect 6878 1056 6886 1120
rect 6950 1056 6966 1120
rect 7030 1056 7046 1120
rect 7110 1056 7126 1120
rect 7190 1056 7198 1120
rect 6878 1040 7198 1056
rect 9845 6016 10165 6576
rect 9845 5952 9853 6016
rect 9917 5952 9933 6016
rect 9997 5952 10013 6016
rect 10077 5952 10093 6016
rect 10157 5952 10165 6016
rect 9845 4928 10165 5952
rect 9845 4864 9853 4928
rect 9917 4864 9933 4928
rect 9997 4864 10013 4928
rect 10077 4864 10093 4928
rect 10157 4864 10165 4928
rect 9845 3840 10165 4864
rect 9845 3776 9853 3840
rect 9917 3776 9933 3840
rect 9997 3776 10013 3840
rect 10077 3776 10093 3840
rect 10157 3776 10165 3840
rect 9845 2752 10165 3776
rect 9845 2688 9853 2752
rect 9917 2688 9933 2752
rect 9997 2688 10013 2752
rect 10077 2688 10093 2752
rect 10157 2688 10165 2752
rect 9845 1664 10165 2688
rect 12812 6560 13132 6576
rect 12812 6496 12820 6560
rect 12884 6496 12900 6560
rect 12964 6496 12980 6560
rect 13044 6496 13060 6560
rect 13124 6496 13132 6560
rect 12812 5472 13132 6496
rect 12812 5408 12820 5472
rect 12884 5408 12900 5472
rect 12964 5408 12980 5472
rect 13044 5408 13060 5472
rect 13124 5408 13132 5472
rect 12812 4384 13132 5408
rect 12812 4320 12820 4384
rect 12884 4320 12900 4384
rect 12964 4320 12980 4384
rect 13044 4320 13060 4384
rect 13124 4320 13132 4384
rect 12812 3296 13132 4320
rect 12812 3232 12820 3296
rect 12884 3232 12900 3296
rect 12964 3232 12980 3296
rect 13044 3232 13060 3296
rect 13124 3232 13132 3296
rect 12203 2412 12269 2413
rect 12203 2348 12204 2412
rect 12268 2410 12269 2412
rect 12571 2412 12637 2413
rect 12571 2410 12572 2412
rect 12268 2350 12572 2410
rect 12268 2348 12269 2350
rect 12203 2347 12269 2348
rect 12571 2348 12572 2350
rect 12636 2348 12637 2412
rect 12571 2347 12637 2348
rect 12812 2208 13132 3232
rect 12812 2144 12820 2208
rect 12884 2144 12900 2208
rect 12964 2144 12980 2208
rect 13044 2144 13060 2208
rect 13124 2144 13132 2208
rect 11099 2004 11165 2005
rect 11099 1940 11100 2004
rect 11164 1940 11165 2004
rect 11099 1939 11165 1940
rect 9845 1600 9853 1664
rect 9917 1600 9933 1664
rect 9997 1600 10013 1664
rect 10077 1600 10093 1664
rect 10157 1600 10165 1664
rect 9845 1040 10165 1600
rect 11102 1138 11162 1939
rect 12812 1120 13132 2144
rect 12812 1056 12820 1120
rect 12884 1056 12900 1120
rect 12964 1056 12980 1120
rect 13044 1056 13060 1120
rect 13124 1056 13132 1120
rect 12812 1040 13132 1056
rect 15779 6016 16099 6576
rect 15779 5952 15787 6016
rect 15851 5952 15867 6016
rect 15931 5952 15947 6016
rect 16011 5952 16027 6016
rect 16091 5952 16099 6016
rect 15779 4928 16099 5952
rect 15779 4864 15787 4928
rect 15851 4864 15867 4928
rect 15931 4864 15947 4928
rect 16011 4864 16027 4928
rect 16091 4864 16099 4928
rect 15779 3840 16099 4864
rect 15779 3776 15787 3840
rect 15851 3776 15867 3840
rect 15931 3776 15947 3840
rect 16011 3776 16027 3840
rect 16091 3776 16099 3840
rect 15779 2752 16099 3776
rect 15779 2688 15787 2752
rect 15851 2688 15867 2752
rect 15931 2688 15947 2752
rect 16011 2688 16027 2752
rect 16091 2688 16099 2752
rect 15779 1664 16099 2688
rect 15779 1600 15787 1664
rect 15851 1600 15867 1664
rect 15931 1600 15947 1664
rect 16011 1600 16027 1664
rect 16091 1600 16099 1664
rect 15779 1040 16099 1600
rect 18746 6560 19066 6576
rect 18746 6496 18754 6560
rect 18818 6496 18834 6560
rect 18898 6496 18914 6560
rect 18978 6496 18994 6560
rect 19058 6496 19066 6560
rect 18746 5472 19066 6496
rect 18746 5408 18754 5472
rect 18818 5408 18834 5472
rect 18898 5408 18914 5472
rect 18978 5408 18994 5472
rect 19058 5408 19066 5472
rect 18746 4384 19066 5408
rect 18746 4320 18754 4384
rect 18818 4320 18834 4384
rect 18898 4320 18914 4384
rect 18978 4320 18994 4384
rect 19058 4320 19066 4384
rect 18746 3296 19066 4320
rect 18746 3232 18754 3296
rect 18818 3232 18834 3296
rect 18898 3232 18914 3296
rect 18978 3232 18994 3296
rect 19058 3232 19066 3296
rect 18746 2208 19066 3232
rect 21713 6016 22033 6576
rect 21713 5952 21721 6016
rect 21785 5952 21801 6016
rect 21865 5952 21881 6016
rect 21945 5952 21961 6016
rect 22025 5952 22033 6016
rect 21713 4928 22033 5952
rect 21713 4864 21721 4928
rect 21785 4864 21801 4928
rect 21865 4864 21881 4928
rect 21945 4864 21961 4928
rect 22025 4864 22033 4928
rect 21713 3840 22033 4864
rect 24680 6560 25000 6576
rect 24680 6496 24688 6560
rect 24752 6496 24768 6560
rect 24832 6496 24848 6560
rect 24912 6496 24928 6560
rect 24992 6496 25000 6560
rect 24680 5472 25000 6496
rect 24680 5408 24688 5472
rect 24752 5408 24768 5472
rect 24832 5408 24848 5472
rect 24912 5408 24928 5472
rect 24992 5408 25000 5472
rect 24680 4384 25000 5408
rect 24680 4320 24688 4384
rect 24752 4320 24768 4384
rect 24832 4320 24848 4384
rect 24912 4320 24928 4384
rect 24992 4320 25000 4384
rect 22139 4180 22205 4181
rect 22139 4116 22140 4180
rect 22204 4116 22205 4180
rect 22139 4115 22205 4116
rect 21713 3776 21721 3840
rect 21785 3776 21801 3840
rect 21865 3776 21881 3840
rect 21945 3776 21961 3840
rect 22025 3776 22033 3840
rect 19195 3092 19261 3093
rect 19195 3028 19196 3092
rect 19260 3028 19261 3092
rect 19195 3027 19261 3028
rect 18746 2144 18754 2208
rect 18818 2144 18834 2208
rect 18898 2144 18914 2208
rect 18978 2144 18994 2208
rect 19058 2144 19066 2208
rect 18746 1120 19066 2144
rect 19198 1189 19258 3027
rect 20667 2956 20733 2957
rect 20667 2892 20668 2956
rect 20732 2892 20733 2956
rect 20667 2891 20733 2892
rect 20670 1325 20730 2891
rect 21713 2752 22033 3776
rect 21713 2688 21721 2752
rect 21785 2688 21801 2752
rect 21865 2688 21881 2752
rect 21945 2688 21961 2752
rect 22025 2688 22033 2752
rect 21713 1664 22033 2688
rect 21713 1600 21721 1664
rect 21785 1600 21801 1664
rect 21865 1600 21881 1664
rect 21945 1600 21961 1664
rect 22025 1600 22033 1664
rect 20667 1324 20733 1325
rect 20667 1260 20668 1324
rect 20732 1260 20733 1324
rect 20667 1259 20733 1260
rect 19195 1188 19261 1189
rect 19195 1124 19196 1188
rect 19260 1124 19261 1188
rect 19195 1123 19261 1124
rect 18746 1056 18754 1120
rect 18818 1056 18834 1120
rect 18898 1056 18914 1120
rect 18978 1056 18994 1120
rect 19058 1056 19066 1120
rect 18746 1040 19066 1056
rect 21713 1040 22033 1600
rect 22142 1325 22202 4115
rect 24680 3296 25000 4320
rect 24680 3232 24688 3296
rect 24752 3232 24768 3296
rect 24832 3232 24848 3296
rect 24912 3232 24928 3296
rect 24992 3232 25000 3296
rect 24680 2208 25000 3232
rect 24680 2144 24688 2208
rect 24752 2144 24768 2208
rect 24832 2144 24848 2208
rect 24912 2144 24928 2208
rect 24992 2144 25000 2208
rect 22139 1324 22205 1325
rect 22139 1260 22140 1324
rect 22204 1260 22205 1324
rect 22139 1259 22205 1260
rect 24680 1120 25000 2144
rect 24680 1056 24688 1120
rect 24752 1056 24768 1120
rect 24832 1056 24848 1120
rect 24912 1056 24928 1120
rect 24992 1056 25000 1120
rect 24680 1040 25000 1056
<< via4 >>
rect 2550 1052 2786 1138
rect 2550 988 2636 1052
rect 2636 988 2700 1052
rect 2700 988 2786 1052
rect 2550 902 2786 988
rect 11014 902 11250 1138
<< metal5 >>
rect 2508 1138 11292 1180
rect 2508 902 2550 1138
rect 2786 902 11014 1138
rect 11250 902 11292 1138
rect 2508 860 11292 902
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 12420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1688980957
transform 1 0 4048 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 17112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _36_
timestamp 1688980957
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _37_
timestamp 1688980957
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 12420 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 19780 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 24104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_10
timestamp 1688980957
transform 1 0 2024 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_138
timestamp 1688980957
transform 1 0 13800 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_231
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_241
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_254
timestamp 1688980957
transform 1 0 24472 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_42
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_96
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_102
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_106
timestamp 1688980957
transform 1 0 10856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_110
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_158
timestamp 1688980957
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_227
timestamp 1688980957
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_253
timestamp 1688980957
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_60
timestamp 1688980957
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_64
timestamp 1688980957
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_68
timestamp 1688980957
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_86
timestamp 1688980957
transform 1 0 9016 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_106
timestamp 1688980957
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_126
timestamp 1688980957
transform 1 0 12696 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_152
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_160
timestamp 1688980957
transform 1 0 15824 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_164
timestamp 1688980957
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_173
timestamp 1688980957
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_185
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_191
timestamp 1688980957
transform 1 0 18676 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_203
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_208
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_253
timestamp 1688980957
transform 1 0 24380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_71
timestamp 1688980957
transform 1 0 7636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_79
timestamp 1688980957
transform 1 0 8372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_96
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_104
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_124
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_150
timestamp 1688980957
transform 1 0 14904 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_158
timestamp 1688980957
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_162
timestamp 1688980957
transform 1 0 16008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_170
timestamp 1688980957
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_175
timestamp 1688980957
transform 1 0 17204 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_183
timestamp 1688980957
transform 1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_206
timestamp 1688980957
transform 1 0 20056 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_218
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_230
timestamp 1688980957
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_242
timestamp 1688980957
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_16
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_35
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_48
timestamp 1688980957
transform 1 0 5520 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_71
timestamp 1688980957
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_85
timestamp 1688980957
transform 1 0 8924 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_97
timestamp 1688980957
transform 1 0 10028 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_126
timestamp 1688980957
transform 1 0 12696 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_136
timestamp 1688980957
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_178
timestamp 1688980957
transform 1 0 17480 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_188
timestamp 1688980957
transform 1 0 18400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_206
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_228
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_240
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 24196 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 22908 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 23000 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 2392 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 3496 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 4600 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 1748 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 2944 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._00_
timestamp 1688980957
transform 1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._01_
timestamp 1688980957
transform 1 0 1472 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._02_
timestamp 1688980957
transform 1 0 6900 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._03_
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._04_
timestamp 1688980957
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._05_
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._06_
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._07_
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._08_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._09_
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._10_
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._11_
timestamp 1688980957
transform 1 0 14168 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._12_
timestamp 1688980957
transform 1 0 5428 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._13_
timestamp 1688980957
transform 1 0 5152 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._14_
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._15_
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._16_
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._17_
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._18_
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._19_
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._20_
timestamp 1688980957
transform 1 0 9752 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._21_
timestamp 1688980957
transform 1 0 9016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._22_
timestamp 1688980957
transform 1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._23_
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix._24_
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._25_
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._26_
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._27_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._28_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._29_
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._30_
timestamp 1688980957
transform 1 0 13524 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._31_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 17664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output59 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 15180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 17572 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 19228 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1688980957
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output70
timestamp 1688980957
transform 1 0 4416 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 10396 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 11776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 13248 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 20884 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 8740 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 23368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 6072 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 15732 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 18216 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 22724 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 24012 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 24288 0 -1 6528
box -38 -48 130 592
<< labels >>
flabel metal2 s 20350 0 20406 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 23110 0 23166 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 23386 0 23442 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 23662 0 23718 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 23938 0 23994 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 24214 0 24270 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 24490 0 24546 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 24766 0 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 25042 0 25098 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 25318 0 25374 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 25594 0 25650 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 20626 0 20682 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 20902 0 20958 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 21178 0 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 21454 0 21510 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 21730 0 21786 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 22006 0 22062 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 22282 0 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 22558 0 22614 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22834 0 22890 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 2134 7840 2190 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 14094 7840 14150 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 15290 7840 15346 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 16486 7840 16542 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 17682 7840 17738 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 18878 7840 18934 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 20074 7840 20130 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 21270 7840 21326 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 22466 7840 22522 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 23662 7840 23718 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 24858 7840 24914 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 3330 7840 3386 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 4526 7840 4582 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 5722 7840 5778 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 6918 7840 6974 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 8114 7840 8170 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 9310 7840 9366 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 10506 7840 10562 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 11702 7840 11758 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 12898 7840 12954 8000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 202 0 258 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 478 0 534 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 754 0 810 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 1030 0 1086 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 3790 0 3846 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 4066 0 4122 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 4342 0 4398 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 4618 0 4674 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 4894 0 4950 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 5170 0 5226 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 5446 0 5502 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 1582 0 1638 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 1858 0 1914 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 2134 0 2190 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 2410 0 2466 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 2686 0 2742 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 2962 0 3018 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 3238 0 3294 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 8482 0 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 8758 0 8814 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 9034 0 9090 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 9310 0 9366 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 9586 0 9642 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 9862 0 9918 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 5998 0 6054 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 6274 0 6330 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 6550 0 6606 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 6826 0 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 7102 0 7158 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 7654 0 7710 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 8206 0 8262 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 76 nsew signal tristate
flabel metal2 s 10414 0 10470 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 77 nsew signal tristate
flabel metal2 s 10690 0 10746 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 78 nsew signal tristate
flabel metal2 s 10966 0 11022 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 79 nsew signal tristate
flabel metal2 s 13450 0 13506 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 80 nsew signal tristate
flabel metal2 s 13726 0 13782 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 81 nsew signal tristate
flabel metal2 s 14002 0 14058 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 82 nsew signal tristate
flabel metal2 s 14278 0 14334 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 83 nsew signal tristate
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 84 nsew signal tristate
flabel metal2 s 14830 0 14886 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 85 nsew signal tristate
flabel metal2 s 15106 0 15162 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 86 nsew signal tristate
flabel metal2 s 15382 0 15438 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 87 nsew signal tristate
flabel metal2 s 11242 0 11298 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 88 nsew signal tristate
flabel metal2 s 11518 0 11574 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 89 nsew signal tristate
flabel metal2 s 11794 0 11850 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 90 nsew signal tristate
flabel metal2 s 12070 0 12126 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 91 nsew signal tristate
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 92 nsew signal tristate
flabel metal2 s 12622 0 12678 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 93 nsew signal tristate
flabel metal2 s 12898 0 12954 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 94 nsew signal tristate
flabel metal2 s 13174 0 13230 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 95 nsew signal tristate
flabel metal2 s 15658 0 15714 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 96 nsew signal tristate
flabel metal2 s 18418 0 18474 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 97 nsew signal tristate
flabel metal2 s 18694 0 18750 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 98 nsew signal tristate
flabel metal2 s 18970 0 19026 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 99 nsew signal tristate
flabel metal2 s 19246 0 19302 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 100 nsew signal tristate
flabel metal2 s 19522 0 19578 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 101 nsew signal tristate
flabel metal2 s 19798 0 19854 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 102 nsew signal tristate
flabel metal2 s 15934 0 15990 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 103 nsew signal tristate
flabel metal2 s 16210 0 16266 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 104 nsew signal tristate
flabel metal2 s 16486 0 16542 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 105 nsew signal tristate
flabel metal2 s 16762 0 16818 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 106 nsew signal tristate
flabel metal2 s 17038 0 17094 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 107 nsew signal tristate
flabel metal2 s 17314 0 17370 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 108 nsew signal tristate
flabel metal2 s 17590 0 17646 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 109 nsew signal tristate
flabel metal2 s 17866 0 17922 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 110 nsew signal tristate
flabel metal2 s 18142 0 18198 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 111 nsew signal tristate
flabel metal2 s 20074 0 20130 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 938 7840 994 8000 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6878 1040 7198 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12812 1040 13132 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18746 1040 19066 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24680 1040 25000 6576 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3911 1040 4231 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9845 1040 10165 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15779 1040 16099 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21713 1040 22033 6576 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 13052 6528 13052 6528 0 VGND
rlabel metal1 12972 5984 12972 5984 0 VPWR
rlabel metal2 20378 364 20378 364 0 FrameStrobe[0]
rlabel metal2 23138 483 23138 483 0 FrameStrobe[10]
rlabel metal2 23414 1044 23414 1044 0 FrameStrobe[11]
rlabel metal2 23690 483 23690 483 0 FrameStrobe[12]
rlabel metal2 23966 432 23966 432 0 FrameStrobe[13]
rlabel metal2 24242 228 24242 228 0 FrameStrobe[14]
rlabel metal1 24288 2958 24288 2958 0 FrameStrobe[15]
rlabel metal2 24695 68 24695 68 0 FrameStrobe[16]
rlabel metal1 24288 3094 24288 3094 0 FrameStrobe[17]
rlabel metal2 25346 772 25346 772 0 FrameStrobe[18]
rlabel metal2 25622 432 25622 432 0 FrameStrobe[19]
rlabel metal2 20601 68 20601 68 0 FrameStrobe[1]
rlabel metal2 20930 432 20930 432 0 FrameStrobe[2]
rlabel metal2 21305 68 21305 68 0 FrameStrobe[3]
rlabel metal2 21482 364 21482 364 0 FrameStrobe[4]
rlabel metal2 21705 68 21705 68 0 FrameStrobe[5]
rlabel metal2 22034 772 22034 772 0 FrameStrobe[6]
rlabel metal2 22363 68 22363 68 0 FrameStrobe[7]
rlabel metal2 22685 68 22685 68 0 FrameStrobe[8]
rlabel metal2 22862 1010 22862 1010 0 FrameStrobe[9]
rlabel metal1 2300 6426 2300 6426 0 FrameStrobe_O[0]
rlabel metal2 14221 7956 14221 7956 0 FrameStrobe_O[10]
rlabel metal2 15371 7956 15371 7956 0 FrameStrobe_O[11]
rlabel metal2 16705 7956 16705 7956 0 FrameStrobe_O[12]
rlabel metal2 17855 7956 17855 7956 0 FrameStrobe_O[13]
rlabel metal2 19189 7956 19189 7956 0 FrameStrobe_O[14]
rlabel metal2 20378 7191 20378 7191 0 FrameStrobe_O[15]
rlabel metal2 21574 7191 21574 7191 0 FrameStrobe_O[16]
rlabel metal2 22547 7956 22547 7956 0 FrameStrobe_O[17]
rlabel metal2 23690 7473 23690 7473 0 FrameStrobe_O[18]
rlabel metal1 24334 5882 24334 5882 0 FrameStrobe_O[19]
rlabel metal2 3595 7956 3595 7956 0 FrameStrobe_O[1]
rlabel metal2 4607 7956 4607 7956 0 FrameStrobe_O[2]
rlabel metal2 5941 7956 5941 7956 0 FrameStrobe_O[3]
rlabel metal2 7137 7956 7137 7956 0 FrameStrobe_O[4]
rlabel metal2 8287 7956 8287 7956 0 FrameStrobe_O[5]
rlabel metal2 9391 7956 9391 7956 0 FrameStrobe_O[6]
rlabel metal2 10587 7956 10587 7956 0 FrameStrobe_O[7]
rlabel metal2 12006 7191 12006 7191 0 FrameStrobe_O[8]
rlabel metal2 13202 7191 13202 7191 0 FrameStrobe_O[9]
rlabel metal2 8234 1530 8234 1530 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG0
rlabel metal1 1610 1326 1610 1326 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 7682 1292 7682 1292 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 7314 1326 7314 1326 0 Inst_N_term_RAM_IO_switch_matrix.S1BEG3
rlabel metal1 11730 2380 11730 2380 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG0
rlabel metal1 12466 1940 12466 1940 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG1
rlabel metal2 9522 1377 9522 1377 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 12282 2380 12282 2380 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG3
rlabel metal1 13294 2482 13294 2482 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 13478 2006 13478 2006 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG5
rlabel metal1 15686 1972 15686 1972 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG6
rlabel metal1 14766 2074 14766 2074 0 Inst_N_term_RAM_IO_switch_matrix.S2BEG7
rlabel metal1 5612 1326 5612 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb0
rlabel metal1 5290 1326 5290 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 4462 1326 4462 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb2
rlabel metal1 4002 1292 4002 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb3
rlabel metal2 2898 1904 2898 1904 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb4
rlabel metal1 4922 1292 4922 1292 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 6670 1326 6670 1326 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb6
rlabel metal1 9614 1930 9614 1930 0 Inst_N_term_RAM_IO_switch_matrix.S2BEGb7
rlabel metal1 10120 1734 10120 1734 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG0
rlabel metal2 16146 1258 16146 1258 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG1
rlabel metal1 18630 1326 18630 1326 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG10
rlabel metal3 15548 1564 15548 1564 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG11
rlabel metal1 18492 2482 18492 2482 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG12
rlabel metal1 19458 2380 19458 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG13
rlabel metal1 20562 2448 20562 2448 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG14
rlabel via2 21850 1445 21850 1445 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG15
rlabel metal1 10442 2380 10442 2380 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG2
rlabel metal2 16330 1258 16330 1258 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG3
rlabel metal1 15272 1938 15272 1938 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG4
rlabel metal1 16422 1530 16422 1530 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG5
rlabel metal1 17342 2448 17342 2448 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG6
rlabel metal1 17526 2074 17526 2074 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG7
rlabel metal1 17802 2074 17802 2074 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG8
rlabel metal1 21344 1530 21344 1530 0 Inst_N_term_RAM_IO_switch_matrix.S4BEG9
rlabel metal2 230 1214 230 1214 0 N1END[0]
rlabel metal2 506 1282 506 1282 0 N1END[1]
rlabel metal2 782 976 782 976 0 N1END[2]
rlabel metal2 1058 942 1058 942 0 N1END[3]
rlabel metal2 3542 296 3542 296 0 N2END[0]
rlabel metal2 3765 68 3765 68 0 N2END[1]
rlabel metal2 3995 68 3995 68 0 N2END[2]
rlabel metal2 4423 68 4423 68 0 N2END[3]
rlabel metal2 4646 1248 4646 1248 0 N2END[4]
rlabel metal2 4922 551 4922 551 0 N2END[5]
rlabel metal2 5145 68 5145 68 0 N2END[6]
rlabel metal2 5375 68 5375 68 0 N2END[7]
rlabel metal2 1334 1248 1334 1248 0 N2MID[0]
rlabel metal2 1709 68 1709 68 0 N2MID[1]
rlabel metal2 1886 670 1886 670 0 N2MID[2]
rlabel metal2 2162 1010 2162 1010 0 N2MID[3]
rlabel metal2 2339 68 2339 68 0 N2MID[4]
rlabel metal2 2714 670 2714 670 0 N2MID[5]
rlabel metal2 3089 68 3089 68 0 N2MID[6]
rlabel metal1 2714 1360 2714 1360 0 N2MID[7]
rlabel metal2 5750 636 5750 636 0 N4END[0]
rlabel metal2 8510 551 8510 551 0 N4END[10]
rlabel metal2 8786 619 8786 619 0 N4END[11]
rlabel metal2 9062 143 9062 143 0 N4END[12]
rlabel metal2 9338 1248 9338 1248 0 N4END[13]
rlabel metal2 9614 636 9614 636 0 N4END[14]
rlabel metal2 9890 143 9890 143 0 N4END[15]
rlabel metal2 6026 279 6026 279 0 N4END[1]
rlabel metal2 6302 976 6302 976 0 N4END[2]
rlabel metal2 6578 1010 6578 1010 0 N4END[3]
rlabel metal2 6854 364 6854 364 0 N4END[4]
rlabel metal2 7130 500 7130 500 0 N4END[5]
rlabel metal2 7406 1010 7406 1010 0 N4END[6]
rlabel metal2 7682 551 7682 551 0 N4END[7]
rlabel metal2 7958 398 7958 398 0 N4END[8]
rlabel metal2 8234 551 8234 551 0 N4END[9]
rlabel metal2 10113 68 10113 68 0 S1BEG[0]
rlabel metal2 10442 908 10442 908 0 S1BEG[1]
rlabel metal2 10718 670 10718 670 0 S1BEG[2]
rlabel metal2 10994 908 10994 908 0 S1BEG[3]
rlabel metal2 13478 636 13478 636 0 S2BEG[0]
rlabel metal2 13754 806 13754 806 0 S2BEG[1]
rlabel metal2 14030 636 14030 636 0 S2BEG[2]
rlabel metal2 14306 908 14306 908 0 S2BEG[3]
rlabel metal2 14681 68 14681 68 0 S2BEG[4]
rlabel metal2 14858 806 14858 806 0 S2BEG[5]
rlabel metal2 15134 296 15134 296 0 S2BEG[6]
rlabel metal2 15410 619 15410 619 0 S2BEG[7]
rlabel metal2 11171 68 11171 68 0 S2BEGb[0]
rlabel metal2 11546 211 11546 211 0 S2BEGb[1]
rlabel metal2 11822 908 11822 908 0 S2BEGb[2]
rlabel metal2 11999 68 11999 68 0 S2BEGb[3]
rlabel metal2 12374 636 12374 636 0 S2BEGb[4]
rlabel metal2 12650 636 12650 636 0 S2BEGb[5]
rlabel metal2 12926 398 12926 398 0 S2BEGb[6]
rlabel metal2 13202 636 13202 636 0 S2BEGb[7]
rlabel metal2 15686 908 15686 908 0 S4BEG[0]
rlabel metal2 18446 670 18446 670 0 S4BEG[10]
rlabel metal1 20654 1428 20654 1428 0 S4BEG[11]
rlabel metal2 18998 483 18998 483 0 S4BEG[12]
rlabel metal2 19274 687 19274 687 0 S4BEG[13]
rlabel metal2 19649 68 19649 68 0 S4BEG[14]
rlabel metal2 19826 806 19826 806 0 S4BEG[15]
rlabel metal2 15962 347 15962 347 0 S4BEG[1]
rlabel metal2 16238 738 16238 738 0 S4BEG[2]
rlabel metal2 16514 636 16514 636 0 S4BEG[3]
rlabel metal2 16790 908 16790 908 0 S4BEG[4]
rlabel metal2 17066 398 17066 398 0 S4BEG[5]
rlabel metal2 17342 347 17342 347 0 S4BEG[6]
rlabel metal2 17618 296 17618 296 0 S4BEG[7]
rlabel metal2 17894 959 17894 959 0 S4BEG[8]
rlabel metal2 18170 483 18170 483 0 S4BEG[9]
rlabel metal2 20102 1299 20102 1299 0 UserCLK
rlabel metal2 1157 7956 1157 7956 0 UserCLKo
rlabel metal1 21344 2074 21344 2074 0 net1
rlabel metal1 23414 2618 23414 2618 0 net10
rlabel metal1 20470 1224 20470 1224 0 net100
rlabel metal1 19458 2006 19458 2006 0 net101
rlabel metal1 20056 1938 20056 1938 0 net102
rlabel metal2 21114 2006 21114 2006 0 net103
rlabel metal1 20516 1326 20516 1326 0 net104
rlabel metal1 16698 1326 16698 1326 0 net105
rlabel metal2 16422 1122 16422 1122 0 net106
rlabel metal1 17388 1326 17388 1326 0 net107
rlabel metal1 16974 1904 16974 1904 0 net108
rlabel metal1 17940 1258 17940 1258 0 net109
rlabel metal2 22954 3604 22954 3604 0 net11
rlabel metal1 19504 1258 19504 1258 0 net110
rlabel metal1 18952 1938 18952 1938 0 net111
rlabel metal1 17940 2006 17940 2006 0 net112
rlabel metal1 18446 2006 18446 2006 0 net113
rlabel metal2 1518 4063 1518 4063 0 net114
rlabel metal1 14628 5202 14628 5202 0 net12
rlabel metal1 22586 1258 22586 1258 0 net13
rlabel metal1 22816 1190 22816 1190 0 net14
rlabel metal2 13294 1870 13294 1870 0 net15
rlabel metal2 17250 3978 17250 3978 0 net16
rlabel metal2 16698 2006 16698 2006 0 net17
rlabel metal2 15180 1530 15180 1530 0 net18
rlabel metal1 13432 5134 13432 5134 0 net19
rlabel metal1 17526 4182 17526 4182 0 net2
rlabel metal2 13662 4318 13662 4318 0 net20
rlabel metal2 3450 1700 3450 1700 0 net21
rlabel metal1 7084 1326 7084 1326 0 net22
rlabel metal1 1702 2006 1702 2006 0 net23
rlabel metal1 8602 1972 8602 1972 0 net24
rlabel metal2 2622 2006 2622 2006 0 net25
rlabel metal1 6900 1938 6900 1938 0 net26
rlabel metal1 4186 1326 4186 1326 0 net27
rlabel metal2 3082 1445 3082 1445 0 net28
rlabel metal1 3358 1428 3358 1428 0 net29
rlabel metal1 16146 5236 16146 5236 0 net3
rlabel metal1 3772 1326 3772 1326 0 net30
rlabel metal1 5382 1904 5382 1904 0 net31
rlabel metal1 5658 1870 5658 1870 0 net32
rlabel via2 1610 2533 1610 2533 0 net33
rlabel metal2 2254 1581 2254 1581 0 net34
rlabel metal1 2438 2312 2438 2312 0 net35
rlabel metal2 2346 1513 2346 1513 0 net36
rlabel metal3 2185 1020 2185 1020 0 net37
rlabel metal2 2070 1088 2070 1088 0 net38
rlabel metal2 12742 1853 12742 1853 0 net39
rlabel metal1 17342 5168 17342 5168 0 net4
rlabel metal1 2346 850 2346 850 0 net40
rlabel metal3 21229 1292 21229 1292 0 net41
rlabel metal1 15502 1190 15502 1190 0 net42
rlabel metal2 13570 1292 13570 1292 0 net43
rlabel metal2 8602 1326 8602 1326 0 net44
rlabel via1 9426 1938 9426 1938 0 net45
rlabel metal1 9062 1360 9062 1360 0 net46
rlabel metal1 9982 1972 9982 1972 0 net47
rlabel via2 19734 2397 19734 2397 0 net48
rlabel metal2 20286 2193 20286 2193 0 net49
rlabel metal1 19642 2550 19642 2550 0 net5
rlabel metal1 5750 1360 5750 1360 0 net50
rlabel metal1 6256 1326 6256 1326 0 net51
rlabel via2 8142 2261 8142 2261 0 net52
rlabel metal3 20355 1156 20355 1156 0 net53
rlabel metal2 7130 1632 7130 1632 0 net54
rlabel metal1 7682 2074 7682 2074 0 net55
rlabel metal2 7866 2312 7866 2312 0 net56
rlabel metal1 20746 2006 20746 2006 0 net57
rlabel metal2 5658 6256 5658 6256 0 net58
rlabel metal1 14582 6358 14582 6358 0 net59
rlabel metal1 23460 1938 23460 1938 0 net6
rlabel metal1 15548 6358 15548 6358 0 net60
rlabel metal1 17020 6358 17020 6358 0 net61
rlabel metal1 17940 6358 17940 6358 0 net62
rlabel metal1 19596 6358 19596 6358 0 net63
rlabel metal1 20194 6324 20194 6324 0 net64
rlabel metal1 21620 6290 21620 6290 0 net65
rlabel metal1 22724 6358 22724 6358 0 net66
rlabel metal1 23874 6392 23874 6392 0 net67
rlabel metal1 24012 5338 24012 5338 0 net68
rlabel metal1 3910 6188 3910 6188 0 net69
rlabel metal1 24150 2414 24150 2414 0 net7
rlabel metal1 12466 6324 12466 6324 0 net70
rlabel metal1 5750 6392 5750 6392 0 net71
rlabel metal1 7176 6358 7176 6358 0 net72
rlabel metal1 8372 6358 8372 6358 0 net73
rlabel metal1 9568 6358 9568 6358 0 net74
rlabel metal1 10764 6358 10764 6358 0 net75
rlabel metal1 12006 6290 12006 6290 0 net76
rlabel metal1 13202 6290 13202 6290 0 net77
rlabel metal1 9614 1292 9614 1292 0 net78
rlabel metal1 1472 1190 1472 1190 0 net79
rlabel metal1 23414 1394 23414 1394 0 net8
rlabel metal2 8970 1513 8970 1513 0 net80
rlabel metal1 10994 2040 10994 2040 0 net81
rlabel metal1 12558 1326 12558 1326 0 net82
rlabel metal1 14214 1360 14214 1360 0 net83
rlabel metal1 13570 850 13570 850 0 net84
rlabel metal1 14490 1904 14490 1904 0 net85
rlabel metal1 14858 1972 14858 1972 0 net86
rlabel metal1 15318 1292 15318 1292 0 net87
rlabel metal1 15686 1326 15686 1326 0 net88
rlabel metal1 15824 2414 15824 2414 0 net89
rlabel metal1 23092 2822 23092 2822 0 net9
rlabel metal2 10810 1122 10810 1122 0 net90
rlabel metal1 10212 1326 10212 1326 0 net91
rlabel metal2 4370 816 4370 816 0 net92
rlabel metal1 3910 1190 3910 1190 0 net93
rlabel metal1 12190 1258 12190 1258 0 net94
rlabel metal2 10074 2227 10074 2227 0 net95
rlabel metal1 11822 1292 11822 1292 0 net96
rlabel metal2 12512 1700 12512 1700 0 net97
rlabel metal1 15870 2040 15870 2040 0 net98
rlabel metal1 19182 1292 19182 1292 0 net99
rlabel metal2 20010 5508 20010 5508 0 strobe_inbuf_0.X
rlabel metal2 14582 5508 14582 5508 0 strobe_inbuf_1.X
rlabel metal2 14858 5508 14858 5508 0 strobe_inbuf_10.X
rlabel metal2 15962 5508 15962 5508 0 strobe_inbuf_11.X
rlabel metal2 17158 5508 17158 5508 0 strobe_inbuf_12.X
rlabel metal2 18446 5508 18446 5508 0 strobe_inbuf_13.X
rlabel metal1 23874 1904 23874 1904 0 strobe_inbuf_14.X
rlabel metal1 24104 1938 24104 1938 0 strobe_inbuf_15.X
rlabel metal2 22034 1887 22034 1887 0 strobe_inbuf_16.X
rlabel metal1 22862 1938 22862 1938 0 strobe_inbuf_17.X
rlabel metal2 24150 3332 24150 3332 0 strobe_inbuf_18.X
rlabel metal1 24242 4556 24242 4556 0 strobe_inbuf_19.X
rlabel metal2 12006 5508 12006 5508 0 strobe_inbuf_2.X
rlabel metal1 6348 5338 6348 5338 0 strobe_inbuf_3.X
rlabel metal2 7590 5508 7590 5508 0 strobe_inbuf_4.X
rlabel metal2 8786 5508 8786 5508 0 strobe_inbuf_5.X
rlabel metal2 9890 5508 9890 5508 0 strobe_inbuf_6.X
rlabel metal2 11086 5508 11086 5508 0 strobe_inbuf_7.X
rlabel metal2 12466 5508 12466 5508 0 strobe_inbuf_8.X
rlabel metal2 13478 5508 13478 5508 0 strobe_inbuf_9.X
rlabel metal1 20194 5882 20194 5882 0 strobe_outbuf_0.X
rlabel metal1 14536 5882 14536 5882 0 strobe_outbuf_1.X
rlabel metal1 14904 5542 14904 5542 0 strobe_outbuf_10.X
rlabel metal1 15732 5882 15732 5882 0 strobe_outbuf_11.X
rlabel metal1 17204 5882 17204 5882 0 strobe_outbuf_12.X
rlabel metal1 18308 5882 18308 5882 0 strobe_outbuf_13.X
rlabel metal2 20010 6052 20010 6052 0 strobe_outbuf_14.X
rlabel metal1 21022 6222 21022 6222 0 strobe_outbuf_15.X
rlabel metal1 21758 2074 21758 2074 0 strobe_outbuf_16.X
rlabel metal1 22954 2074 22954 2074 0 strobe_outbuf_17.X
rlabel metal1 23828 3706 23828 3706 0 strobe_outbuf_18.X
rlabel metal1 24196 4794 24196 4794 0 strobe_outbuf_19.X
rlabel metal1 12650 5848 12650 5848 0 strobe_outbuf_2.X
rlabel metal1 6348 5882 6348 5882 0 strobe_outbuf_3.X
rlabel metal1 7498 5882 7498 5882 0 strobe_outbuf_4.X
rlabel metal1 8694 5882 8694 5882 0 strobe_outbuf_5.X
rlabel metal2 9706 6086 9706 6086 0 strobe_outbuf_6.X
rlabel metal1 11040 5882 11040 5882 0 strobe_outbuf_7.X
rlabel metal1 12328 5882 12328 5882 0 strobe_outbuf_8.X
rlabel metal1 13432 5882 13432 5882 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 26000 8000
<< end >>
