magic
tech sky130A
magscale 1 2
timestamp 1732489020
<< viali >>
rect 2697 43401 2731 43435
rect 3065 43401 3099 43435
rect 3985 43401 4019 43435
rect 4537 43401 4571 43435
rect 5273 43401 5307 43435
rect 6009 43401 6043 43435
rect 6745 43401 6779 43435
rect 7481 43401 7515 43435
rect 8217 43401 8251 43435
rect 9137 43401 9171 43435
rect 9689 43401 9723 43435
rect 10425 43401 10459 43435
rect 11713 43401 11747 43435
rect 12633 43401 12667 43435
rect 13369 43401 13403 43435
rect 14289 43401 14323 43435
rect 1501 43265 1535 43299
rect 2145 43265 2179 43299
rect 2513 43265 2547 43299
rect 2973 43265 3007 43299
rect 3801 43265 3835 43299
rect 4353 43265 4387 43299
rect 5089 43265 5123 43299
rect 5825 43265 5859 43299
rect 6561 43265 6595 43299
rect 7297 43265 7331 43299
rect 8033 43265 8067 43299
rect 8953 43265 8987 43299
rect 9597 43265 9631 43299
rect 10241 43265 10275 43299
rect 11621 43265 11655 43299
rect 12081 43265 12115 43299
rect 12541 43265 12575 43299
rect 13185 43265 13219 43299
rect 13645 43265 13679 43299
rect 14105 43265 14139 43299
rect 2329 43129 2363 43163
rect 13829 43129 13863 43163
rect 1593 43061 1627 43095
rect 12265 43061 12299 43095
rect 2053 42857 2087 42891
rect 2789 42857 2823 42891
rect 3341 42857 3375 42891
rect 4169 42857 4203 42891
rect 5733 42857 5767 42891
rect 6469 42857 6503 42891
rect 7113 42857 7147 42891
rect 7849 42857 7883 42891
rect 8585 42857 8619 42891
rect 9321 42857 9355 42891
rect 10057 42857 10091 42891
rect 10793 42857 10827 42891
rect 12265 42857 12299 42891
rect 13001 42857 13035 42891
rect 14289 42857 14323 42891
rect 11529 42789 11563 42823
rect 12725 42789 12759 42823
rect 13829 42721 13863 42755
rect 2237 42653 2271 42687
rect 2973 42653 3007 42687
rect 3525 42653 3559 42687
rect 4353 42653 4387 42687
rect 5917 42653 5951 42687
rect 6653 42653 6687 42687
rect 7297 42653 7331 42687
rect 8033 42653 8067 42687
rect 8769 42653 8803 42687
rect 9505 42653 9539 42687
rect 10241 42653 10275 42687
rect 10977 42653 11011 42687
rect 11713 42653 11747 42687
rect 12449 42653 12483 42687
rect 12909 42653 12943 42687
rect 13185 42653 13219 42687
rect 14473 42653 14507 42687
rect 13553 42585 13587 42619
rect 2053 42313 2087 42347
rect 2881 42313 2915 42347
rect 5549 42313 5583 42347
rect 6377 42313 6411 42347
rect 7113 42313 7147 42347
rect 7941 42313 7975 42347
rect 8677 42313 8711 42347
rect 9321 42313 9355 42347
rect 10149 42313 10183 42347
rect 10793 42313 10827 42347
rect 11529 42313 11563 42347
rect 12265 42313 12299 42347
rect 12909 42313 12943 42347
rect 14013 42313 14047 42347
rect 14289 42313 14323 42347
rect 2237 42177 2271 42211
rect 3065 42177 3099 42211
rect 5733 42177 5767 42211
rect 6561 42177 6595 42211
rect 7297 42177 7331 42211
rect 8125 42177 8159 42211
rect 8861 42177 8895 42211
rect 9505 42177 9539 42211
rect 10333 42177 10367 42211
rect 10977 42177 11011 42211
rect 11713 42177 11747 42211
rect 12449 42177 12483 42211
rect 13093 42177 13127 42211
rect 13461 42177 13495 42211
rect 13921 42177 13955 42211
rect 14197 42177 14231 42211
rect 14473 42177 14507 42211
rect 13737 42041 13771 42075
rect 2881 41769 2915 41803
rect 14289 41769 14323 41803
rect 3065 41565 3099 41599
rect 14473 41565 14507 41599
rect 1409 41089 1443 41123
rect 1593 40885 1627 40919
rect 1409 40001 1443 40035
rect 13369 40001 13403 40035
rect 13921 40001 13955 40035
rect 1593 39797 1627 39831
rect 13645 39797 13679 39831
rect 14197 39797 14231 39831
rect 8953 39593 8987 39627
rect 9505 39593 9539 39627
rect 7389 39525 7423 39559
rect 8125 39525 8159 39559
rect 9229 39525 9263 39559
rect 13093 39525 13127 39559
rect 1409 39389 1443 39423
rect 7573 39389 7607 39423
rect 8309 39389 8343 39423
rect 8585 39389 8619 39423
rect 9137 39389 9171 39423
rect 9413 39389 9447 39423
rect 9689 39389 9723 39423
rect 12725 39389 12759 39423
rect 13001 39389 13035 39423
rect 13277 39389 13311 39423
rect 14197 39389 14231 39423
rect 13553 39321 13587 39355
rect 13921 39321 13955 39355
rect 1593 39253 1627 39287
rect 8401 39253 8435 39287
rect 12541 39253 12575 39287
rect 12817 39253 12851 39287
rect 14381 39253 14415 39287
rect 4997 39049 5031 39083
rect 11989 39049 12023 39083
rect 12817 39049 12851 39083
rect 13921 38981 13955 39015
rect 5181 38913 5215 38947
rect 12173 38913 12207 38947
rect 12449 38913 12483 38947
rect 12725 38913 12759 38947
rect 13001 38913 13035 38947
rect 13369 38913 13403 38947
rect 12265 38777 12299 38811
rect 12541 38709 12575 38743
rect 13645 38709 13679 38743
rect 14197 38709 14231 38743
rect 4813 38505 4847 38539
rect 12541 38505 12575 38539
rect 13001 38437 13035 38471
rect 1409 38301 1443 38335
rect 4997 38301 5031 38335
rect 12449 38301 12483 38335
rect 12725 38301 12759 38335
rect 13185 38301 13219 38335
rect 13553 38301 13587 38335
rect 13645 38301 13679 38335
rect 14197 38301 14231 38335
rect 1593 38165 1627 38199
rect 12265 38165 12299 38199
rect 13369 38165 13403 38199
rect 13829 38165 13863 38199
rect 14381 38165 14415 38199
rect 11529 37961 11563 37995
rect 11897 37961 11931 37995
rect 12357 37961 12391 37995
rect 12633 37961 12667 37995
rect 12909 37961 12943 37995
rect 13369 37893 13403 37927
rect 1409 37825 1443 37859
rect 11713 37825 11747 37859
rect 12081 37825 12115 37859
rect 12541 37825 12575 37859
rect 12817 37825 12851 37859
rect 13093 37825 13127 37859
rect 13921 37825 13955 37859
rect 1593 37621 1627 37655
rect 13645 37621 13679 37655
rect 14197 37621 14231 37655
rect 10793 37417 10827 37451
rect 11161 37417 11195 37451
rect 12357 37417 12391 37451
rect 12633 37417 12667 37451
rect 10977 37213 11011 37247
rect 11345 37213 11379 37247
rect 12541 37213 12575 37247
rect 12817 37213 12851 37247
rect 13093 37213 13127 37247
rect 13369 37213 13403 37247
rect 14197 37213 14231 37247
rect 13553 37145 13587 37179
rect 12909 37077 12943 37111
rect 13185 37077 13219 37111
rect 13645 37077 13679 37111
rect 14381 37077 14415 37111
rect 2145 36873 2179 36907
rect 9965 36873 9999 36907
rect 11621 36873 11655 36907
rect 11897 36873 11931 36907
rect 12173 36873 12207 36907
rect 1409 36737 1443 36771
rect 2329 36737 2363 36771
rect 10149 36737 10183 36771
rect 11805 36737 11839 36771
rect 12081 36737 12115 36771
rect 12333 36737 12367 36771
rect 12725 36737 12759 36771
rect 13001 36737 13035 36771
rect 13369 36737 13403 36771
rect 13553 36737 13587 36771
rect 14105 36737 14139 36771
rect 13185 36601 13219 36635
rect 1593 36533 1627 36567
rect 12541 36533 12575 36567
rect 12817 36533 12851 36567
rect 13829 36533 13863 36567
rect 14381 36533 14415 36567
rect 1593 36329 1627 36363
rect 12173 36329 12207 36363
rect 1409 36125 1443 36159
rect 12357 36125 12391 36159
rect 12633 36125 12667 36159
rect 13093 36125 13127 36159
rect 13369 36125 13403 36159
rect 14197 36125 14231 36159
rect 13553 36057 13587 36091
rect 12449 35989 12483 36023
rect 12909 35989 12943 36023
rect 13185 35989 13219 36023
rect 13829 35989 13863 36023
rect 14381 35989 14415 36023
rect 10241 35785 10275 35819
rect 10425 35649 10459 35683
rect 10701 35649 10735 35683
rect 11803 35649 11837 35683
rect 13001 35649 13035 35683
rect 13553 35649 13587 35683
rect 14105 35649 14139 35683
rect 11529 35581 11563 35615
rect 10517 35445 10551 35479
rect 12541 35445 12575 35479
rect 13277 35445 13311 35479
rect 13829 35445 13863 35479
rect 14381 35445 14415 35479
rect 1777 35241 1811 35275
rect 9505 35241 9539 35275
rect 11989 35241 12023 35275
rect 1593 35173 1627 35207
rect 9781 35173 9815 35207
rect 12265 35173 12299 35207
rect 12633 35173 12667 35207
rect 1409 35037 1443 35071
rect 1961 35037 1995 35071
rect 9689 35037 9723 35071
rect 9965 35037 9999 35071
rect 11897 35037 11931 35071
rect 12173 35037 12207 35071
rect 12449 35037 12483 35071
rect 12817 35037 12851 35071
rect 13093 35037 13127 35071
rect 13369 35037 13403 35071
rect 14289 35037 14323 35071
rect 13553 34969 13587 35003
rect 13921 34969 13955 35003
rect 11713 34901 11747 34935
rect 12909 34901 12943 34935
rect 13185 34901 13219 34935
rect 14105 34901 14139 34935
rect 1593 34697 1627 34731
rect 1777 34697 1811 34731
rect 8769 34697 8803 34731
rect 9781 34697 9815 34731
rect 10517 34697 10551 34731
rect 10977 34697 11011 34731
rect 11621 34697 11655 34731
rect 13001 34697 13035 34731
rect 13921 34629 13955 34663
rect 1409 34561 1443 34595
rect 1961 34561 1995 34595
rect 8953 34561 8987 34595
rect 9229 34561 9263 34595
rect 9505 34561 9539 34595
rect 9965 34561 9999 34595
rect 10701 34561 10735 34595
rect 11161 34561 11195 34595
rect 11805 34561 11839 34595
rect 12265 34561 12299 34595
rect 12541 34561 12575 34595
rect 12817 34561 12851 34595
rect 13185 34561 13219 34595
rect 13369 34561 13403 34595
rect 9045 34425 9079 34459
rect 9321 34425 9355 34459
rect 12081 34425 12115 34459
rect 12357 34425 12391 34459
rect 12633 34357 12667 34391
rect 13645 34357 13679 34391
rect 14197 34357 14231 34391
rect 1593 34153 1627 34187
rect 9229 34153 9263 34187
rect 10517 34153 10551 34187
rect 8953 34085 8987 34119
rect 10241 34085 10275 34119
rect 12633 34085 12667 34119
rect 13001 34085 13035 34119
rect 1777 33949 1811 33983
rect 9137 33949 9171 33983
rect 9413 33949 9447 33983
rect 10425 33949 10459 33983
rect 10701 33949 10735 33983
rect 10977 33949 11011 33983
rect 11621 33949 11655 33983
rect 11895 33949 11929 33983
rect 13185 33949 13219 33983
rect 13553 33949 13587 33983
rect 14197 33949 14231 33983
rect 13921 33881 13955 33915
rect 10793 33813 10827 33847
rect 14381 33813 14415 33847
rect 1593 33609 1627 33643
rect 8125 33609 8159 33643
rect 9597 33609 9631 33643
rect 9873 33609 9907 33643
rect 10425 33609 10459 33643
rect 13921 33541 13955 33575
rect 1409 33473 1443 33507
rect 8309 33473 8343 33507
rect 9781 33473 9815 33507
rect 10057 33473 10091 33507
rect 10609 33473 10643 33507
rect 11161 33473 11195 33507
rect 11803 33473 11837 33507
rect 13185 33473 13219 33507
rect 13369 33473 13403 33507
rect 11529 33405 11563 33439
rect 10977 33337 11011 33371
rect 12541 33269 12575 33303
rect 13001 33269 13035 33303
rect 13645 33269 13679 33303
rect 14197 33269 14231 33303
rect 10057 33065 10091 33099
rect 10885 33065 10919 33099
rect 11161 33065 11195 33099
rect 12265 33065 12299 33099
rect 11437 32997 11471 33031
rect 11713 32997 11747 33031
rect 11989 32997 12023 33031
rect 13185 32997 13219 33031
rect 1409 32861 1443 32895
rect 10241 32861 10275 32895
rect 11069 32861 11103 32895
rect 11345 32861 11379 32895
rect 11621 32861 11655 32895
rect 11897 32861 11931 32895
rect 12173 32861 12207 32895
rect 12449 32861 12483 32895
rect 12725 32861 12759 32895
rect 13001 32861 13035 32895
rect 13369 32861 13403 32895
rect 14105 32861 14139 32895
rect 13553 32793 13587 32827
rect 13921 32793 13955 32827
rect 1593 32725 1627 32759
rect 12541 32725 12575 32759
rect 12817 32725 12851 32759
rect 14289 32725 14323 32759
rect 8033 32385 8067 32419
rect 8291 32415 8325 32449
rect 9671 32415 9705 32449
rect 11345 32385 11379 32419
rect 11803 32385 11837 32419
rect 13185 32385 13219 32419
rect 13737 32385 13771 32419
rect 14197 32385 14231 32419
rect 9413 32317 9447 32351
rect 11529 32317 11563 32351
rect 9045 32181 9079 32215
rect 10425 32181 10459 32215
rect 11161 32181 11195 32215
rect 12541 32181 12575 32215
rect 13461 32181 13495 32215
rect 14013 32181 14047 32215
rect 14381 32181 14415 32215
rect 1593 31977 1627 32011
rect 12173 31977 12207 32011
rect 12633 31977 12667 32011
rect 7941 31909 7975 31943
rect 11345 31909 11379 31943
rect 11621 31909 11655 31943
rect 11897 31909 11931 31943
rect 6929 31841 6963 31875
rect 1409 31773 1443 31807
rect 7203 31773 7237 31807
rect 11529 31773 11563 31807
rect 11805 31773 11839 31807
rect 12081 31773 12115 31807
rect 12357 31773 12391 31807
rect 12817 31773 12851 31807
rect 13001 31773 13035 31807
rect 14381 31773 14415 31807
rect 13553 31705 13587 31739
rect 13277 31637 13311 31671
rect 13829 31637 13863 31671
rect 14197 31637 14231 31671
rect 10977 31433 11011 31467
rect 13369 31365 13403 31399
rect 13921 31365 13955 31399
rect 1409 31297 1443 31331
rect 7539 31297 7573 31331
rect 8935 31327 8969 31361
rect 11161 31297 11195 31331
rect 11771 31297 11805 31331
rect 13093 31297 13127 31331
rect 7297 31229 7331 31263
rect 8677 31229 8711 31263
rect 11529 31229 11563 31263
rect 1593 31093 1627 31127
rect 8309 31093 8343 31127
rect 9689 31093 9723 31127
rect 12541 31093 12575 31127
rect 12909 31093 12943 31127
rect 13645 31093 13679 31127
rect 14197 31093 14231 31127
rect 10333 30889 10367 30923
rect 10977 30889 11011 30923
rect 11529 30889 11563 30923
rect 11805 30889 11839 30923
rect 12081 30889 12115 30923
rect 9505 30821 9539 30855
rect 9689 30685 9723 30719
rect 10241 30685 10275 30719
rect 10517 30685 10551 30719
rect 10885 30685 10919 30719
rect 11161 30685 11195 30719
rect 11713 30685 11747 30719
rect 11989 30685 12023 30719
rect 12265 30685 12299 30719
rect 12449 30685 12483 30719
rect 14197 30685 14231 30719
rect 12817 30617 12851 30651
rect 13001 30617 13035 30651
rect 13369 30617 13403 30651
rect 13553 30617 13587 30651
rect 13921 30617 13955 30651
rect 10057 30549 10091 30583
rect 10701 30549 10735 30583
rect 14381 30549 14415 30583
rect 13461 30345 13495 30379
rect 1409 30209 1443 30243
rect 6377 30209 6411 30243
rect 6651 30209 6685 30243
rect 9137 30209 9171 30243
rect 10425 30209 10459 30243
rect 12817 30209 12851 30243
rect 14013 30209 14047 30243
rect 9229 30141 9263 30175
rect 9413 30141 9447 30175
rect 9873 30141 9907 30175
rect 10149 30141 10183 30175
rect 10287 30141 10321 30175
rect 11621 30141 11655 30175
rect 11805 30141 11839 30175
rect 12541 30141 12575 30175
rect 12679 30141 12713 30175
rect 1593 30073 1627 30107
rect 8953 30073 8987 30107
rect 12265 30073 12299 30107
rect 13829 30073 13863 30107
rect 7389 30005 7423 30039
rect 11069 30005 11103 30039
rect 14289 30005 14323 30039
rect 1593 29801 1627 29835
rect 10793 29801 10827 29835
rect 11345 29801 11379 29835
rect 13461 29801 13495 29835
rect 7573 29733 7607 29767
rect 8769 29733 8803 29767
rect 9597 29733 9631 29767
rect 12265 29733 12299 29767
rect 5549 29665 5583 29699
rect 7966 29665 8000 29699
rect 9137 29665 9171 29699
rect 10149 29665 10183 29699
rect 11805 29665 11839 29699
rect 12541 29665 12575 29699
rect 12817 29665 12851 29699
rect 1409 29597 1443 29631
rect 5823 29597 5857 29631
rect 6929 29597 6963 29631
rect 7113 29597 7147 29631
rect 7849 29597 7883 29631
rect 8125 29597 8159 29631
rect 8953 29597 8987 29631
rect 9873 29597 9907 29631
rect 10011 29597 10045 29631
rect 11069 29597 11103 29631
rect 11529 29597 11563 29631
rect 11621 29597 11655 29631
rect 12658 29597 12692 29631
rect 13737 29597 13771 29631
rect 14289 29597 14323 29631
rect 6561 29461 6595 29495
rect 10885 29461 10919 29495
rect 13553 29461 13587 29495
rect 14105 29461 14139 29495
rect 12081 29257 12115 29291
rect 12725 29257 12759 29291
rect 13001 29257 13035 29291
rect 8677 29189 8711 29223
rect 13369 29189 13403 29223
rect 13921 29189 13955 29223
rect 7874 29121 7908 29155
rect 8033 29121 8067 29155
rect 9011 29121 9045 29155
rect 11989 29121 12023 29155
rect 12265 29121 12299 29155
rect 12633 29121 12667 29155
rect 12909 29121 12943 29155
rect 13185 29121 13219 29155
rect 6837 29053 6871 29087
rect 7021 29053 7055 29087
rect 7481 29053 7515 29087
rect 7757 29053 7791 29087
rect 8769 29053 8803 29087
rect 11805 28985 11839 29019
rect 12449 28985 12483 29019
rect 9781 28917 9815 28951
rect 13645 28917 13679 28951
rect 14197 28917 14231 28951
rect 7665 28713 7699 28747
rect 13553 28713 13587 28747
rect 10425 28645 10459 28679
rect 12357 28645 12391 28679
rect 6653 28577 6687 28611
rect 9781 28577 9815 28611
rect 11713 28577 11747 28611
rect 12750 28577 12784 28611
rect 1409 28509 1443 28543
rect 6911 28509 6945 28543
rect 9965 28509 9999 28543
rect 10701 28509 10735 28543
rect 10818 28509 10852 28543
rect 10977 28509 11011 28543
rect 11897 28509 11931 28543
rect 12633 28509 12667 28543
rect 12909 28509 12943 28543
rect 13645 28509 13679 28543
rect 14197 28509 14231 28543
rect 1593 28373 1627 28407
rect 11621 28373 11655 28407
rect 13829 28373 13863 28407
rect 14381 28373 14415 28407
rect 10701 28169 10735 28203
rect 12725 28169 12759 28203
rect 13921 28101 13955 28135
rect 1501 28033 1535 28067
rect 8033 28033 8067 28067
rect 8307 28033 8341 28067
rect 9963 28033 9997 28067
rect 11971 28063 12005 28097
rect 13369 28033 13403 28067
rect 9689 27965 9723 27999
rect 11713 27965 11747 27999
rect 1593 27829 1627 27863
rect 9045 27829 9079 27863
rect 13645 27829 13679 27863
rect 14197 27829 14231 27863
rect 11345 27625 11379 27659
rect 11897 27625 11931 27659
rect 6101 27421 6135 27455
rect 6359 27391 6393 27425
rect 8953 27421 8987 27455
rect 9195 27421 9229 27455
rect 11529 27421 11563 27455
rect 11805 27421 11839 27455
rect 12081 27421 12115 27455
rect 12357 27421 12391 27455
rect 12817 27421 12851 27455
rect 13093 27421 13127 27455
rect 13369 27421 13403 27455
rect 13553 27421 13587 27455
rect 14197 27421 14231 27455
rect 13921 27353 13955 27387
rect 7113 27285 7147 27319
rect 9965 27285 9999 27319
rect 11621 27285 11655 27319
rect 12173 27285 12207 27319
rect 12633 27285 12667 27319
rect 12909 27285 12943 27319
rect 13185 27285 13219 27319
rect 14381 27285 14415 27319
rect 8493 27081 8527 27115
rect 10425 27081 10459 27115
rect 12081 27081 12115 27115
rect 12449 27013 12483 27047
rect 13001 27013 13035 27047
rect 1501 26945 1535 26979
rect 6837 26945 6871 26979
rect 9781 26945 9815 26979
rect 11989 26945 12023 26979
rect 12265 26945 12299 26979
rect 13553 26945 13587 26979
rect 14105 26945 14139 26979
rect 6653 26877 6687 26911
rect 7297 26877 7331 26911
rect 7573 26877 7607 26911
rect 7711 26877 7745 26911
rect 7849 26877 7883 26911
rect 8585 26877 8619 26911
rect 8769 26877 8803 26911
rect 9229 26877 9263 26911
rect 9505 26877 9539 26911
rect 9622 26877 9656 26911
rect 11805 26809 11839 26843
rect 1593 26741 1627 26775
rect 12541 26741 12575 26775
rect 13277 26741 13311 26775
rect 13829 26741 13863 26775
rect 14381 26741 14415 26775
rect 7481 26537 7515 26571
rect 10885 26469 10919 26503
rect 9873 26401 9907 26435
rect 11253 26401 11287 26435
rect 12633 26401 12667 26435
rect 6469 26333 6503 26367
rect 6711 26333 6745 26367
rect 10147 26333 10181 26367
rect 11511 26333 11545 26367
rect 12875 26333 12909 26367
rect 14197 26333 14231 26367
rect 1501 26265 1535 26299
rect 1685 26265 1719 26299
rect 12265 26197 12299 26231
rect 13645 26197 13679 26231
rect 14381 26197 14415 26231
rect 13369 25993 13403 26027
rect 14105 25925 14139 25959
rect 6635 25887 6669 25921
rect 8033 25857 8067 25891
rect 8307 25857 8341 25891
rect 10057 25857 10091 25891
rect 10315 25887 10349 25921
rect 11529 25857 11563 25891
rect 12725 25857 12759 25891
rect 13553 25857 13587 25891
rect 6377 25789 6411 25823
rect 11713 25789 11747 25823
rect 12449 25789 12483 25823
rect 12566 25789 12600 25823
rect 12173 25721 12207 25755
rect 7389 25653 7423 25687
rect 9045 25653 9079 25687
rect 11069 25653 11103 25687
rect 13829 25653 13863 25687
rect 14381 25653 14415 25687
rect 7481 25449 7515 25483
rect 5273 25381 5307 25415
rect 6285 25381 6319 25415
rect 12541 25381 12575 25415
rect 1685 25313 1719 25347
rect 6837 25313 6871 25347
rect 12081 25313 12115 25347
rect 12817 25313 12851 25347
rect 13093 25313 13127 25347
rect 1409 25245 1443 25279
rect 4261 25245 4295 25279
rect 4535 25245 4569 25279
rect 5641 25245 5675 25279
rect 5825 25245 5859 25279
rect 6561 25245 6595 25279
rect 6699 25245 6733 25279
rect 11897 25245 11931 25279
rect 12934 25245 12968 25279
rect 14197 25245 14231 25279
rect 13737 25109 13771 25143
rect 14381 25109 14415 25143
rect 1685 24837 1719 24871
rect 1501 24769 1535 24803
rect 6927 24769 6961 24803
rect 8033 24769 8067 24803
rect 9229 24769 9263 24803
rect 10207 24769 10241 24803
rect 12081 24769 12115 24803
rect 12447 24769 12481 24803
rect 13737 24769 13771 24803
rect 13921 24769 13955 24803
rect 6653 24701 6687 24735
rect 8217 24701 8251 24735
rect 8953 24701 8987 24735
rect 9091 24701 9125 24735
rect 9965 24701 9999 24735
rect 12173 24701 12207 24735
rect 7665 24633 7699 24667
rect 8677 24633 8711 24667
rect 13553 24633 13587 24667
rect 9873 24565 9907 24599
rect 10977 24565 11011 24599
rect 11897 24565 11931 24599
rect 13185 24565 13219 24599
rect 14197 24565 14231 24599
rect 11529 24361 11563 24395
rect 13093 24293 13127 24327
rect 7481 24225 7515 24259
rect 10333 24225 10367 24259
rect 10726 24225 10760 24259
rect 10885 24225 10919 24259
rect 11621 24225 11655 24259
rect 7723 24157 7757 24191
rect 9689 24157 9723 24191
rect 9873 24157 9907 24191
rect 10609 24157 10643 24191
rect 11863 24157 11897 24191
rect 13277 24157 13311 24191
rect 14197 24157 14231 24191
rect 13553 24089 13587 24123
rect 13921 24089 13955 24123
rect 8493 24021 8527 24055
rect 12633 24021 12667 24055
rect 14381 24021 14415 24055
rect 10149 23817 10183 23851
rect 14105 23749 14139 23783
rect 1685 23681 1719 23715
rect 7203 23681 7237 23715
rect 9379 23681 9413 23715
rect 11989 23681 12023 23715
rect 13185 23681 13219 23715
rect 1409 23613 1443 23647
rect 6929 23613 6963 23647
rect 9137 23613 9171 23647
rect 12173 23613 12207 23647
rect 12633 23613 12667 23647
rect 12909 23613 12943 23647
rect 13026 23613 13060 23647
rect 7941 23477 7975 23511
rect 13829 23477 13863 23511
rect 14381 23477 14415 23511
rect 13369 23273 13403 23307
rect 5273 23205 5307 23239
rect 6285 23205 6319 23239
rect 13093 23205 13127 23239
rect 14381 23205 14415 23239
rect 6561 23137 6595 23171
rect 6699 23137 6733 23171
rect 10885 23137 10919 23171
rect 4261 23069 4295 23103
rect 4535 23069 4569 23103
rect 5641 23069 5675 23103
rect 5825 23069 5859 23103
rect 6837 23069 6871 23103
rect 9505 23069 9539 23103
rect 9779 23059 9813 23093
rect 11159 23069 11193 23103
rect 13277 23069 13311 23103
rect 13553 23069 13587 23103
rect 13645 23069 13679 23103
rect 14197 23069 14231 23103
rect 1501 23001 1535 23035
rect 7481 23001 7515 23035
rect 1593 22933 1627 22967
rect 10517 22933 10551 22967
rect 11897 22933 11931 22967
rect 13829 22933 13863 22967
rect 13277 22729 13311 22763
rect 7665 22593 7699 22627
rect 8861 22593 8895 22627
rect 13185 22593 13219 22627
rect 13461 22593 13495 22627
rect 13737 22593 13771 22627
rect 13921 22593 13955 22627
rect 7849 22525 7883 22559
rect 8309 22525 8343 22559
rect 8585 22525 8619 22559
rect 8702 22525 8736 22559
rect 9505 22525 9539 22559
rect 13553 22457 13587 22491
rect 13001 22389 13035 22423
rect 14197 22389 14231 22423
rect 6469 22185 6503 22219
rect 11437 22185 11471 22219
rect 13645 22185 13679 22219
rect 14381 22185 14415 22219
rect 12449 22117 12483 22151
rect 5457 22049 5491 22083
rect 10425 22049 10459 22083
rect 12725 22049 12759 22083
rect 1685 21981 1719 22015
rect 3157 21981 3191 22015
rect 5731 21981 5765 22015
rect 6837 21981 6871 22015
rect 7111 21981 7145 22015
rect 10699 21981 10733 22015
rect 11805 21981 11839 22015
rect 11989 21981 12023 22015
rect 12863 21981 12897 22015
rect 13001 21981 13035 22015
rect 13921 21981 13955 22015
rect 14197 21981 14231 22015
rect 1501 21913 1535 21947
rect 3341 21845 3375 21879
rect 7849 21845 7883 21879
rect 13737 21845 13771 21879
rect 2697 21641 2731 21675
rect 3249 21641 3283 21675
rect 9321 21641 9355 21675
rect 10149 21641 10183 21675
rect 12725 21641 12759 21675
rect 13277 21641 13311 21675
rect 14381 21641 14415 21675
rect 1409 21573 1443 21607
rect 3433 21505 3467 21539
rect 7481 21505 7515 21539
rect 8401 21505 8435 21539
rect 8518 21505 8552 21539
rect 8677 21505 8711 21539
rect 10057 21505 10091 21539
rect 10333 21505 10367 21539
rect 11713 21505 11747 21539
rect 11971 21535 12005 21569
rect 13093 21505 13127 21539
rect 13553 21505 13587 21539
rect 14105 21505 14139 21539
rect 7665 21437 7699 21471
rect 8125 21437 8159 21471
rect 9873 21301 9907 21335
rect 13829 21301 13863 21335
rect 1593 21097 1627 21131
rect 5825 21097 5859 21131
rect 8493 21097 8527 21131
rect 9597 21097 9631 21131
rect 14381 21097 14415 21131
rect 10793 21029 10827 21063
rect 4445 20961 4479 20995
rect 5917 20961 5951 20995
rect 7481 20961 7515 20995
rect 10057 20961 10091 20995
rect 11345 20961 11379 20995
rect 1501 20893 1535 20927
rect 6159 20893 6193 20927
rect 7755 20893 7789 20927
rect 9505 20893 9539 20927
rect 9689 20893 9723 20927
rect 9781 20893 9815 20927
rect 9873 20893 9907 20927
rect 10149 20893 10183 20927
rect 10333 20893 10367 20927
rect 11069 20893 11103 20927
rect 11207 20893 11241 20927
rect 11989 20893 12023 20927
rect 12357 20893 12391 20927
rect 12449 20893 12483 20927
rect 12723 20893 12757 20927
rect 14197 20893 14231 20927
rect 4690 20825 4724 20859
rect 6929 20757 6963 20791
rect 10057 20757 10091 20791
rect 12173 20757 12207 20791
rect 13461 20757 13495 20791
rect 5549 20553 5583 20587
rect 8125 20553 8159 20587
rect 10609 20553 10643 20587
rect 11713 20553 11747 20587
rect 14289 20553 14323 20587
rect 1501 20417 1535 20451
rect 1685 20417 1719 20451
rect 5457 20417 5491 20451
rect 6009 20417 6043 20451
rect 6561 20417 6595 20451
rect 7113 20417 7147 20451
rect 7387 20417 7421 20451
rect 10517 20417 10551 20451
rect 11069 20417 11103 20451
rect 11897 20417 11931 20451
rect 12173 20417 12207 20451
rect 13277 20417 13311 20451
rect 13553 20417 13587 20451
rect 14473 20417 14507 20451
rect 6837 20349 6871 20383
rect 12357 20349 12391 20383
rect 12541 20349 12575 20383
rect 13394 20349 13428 20383
rect 10885 20281 10919 20315
rect 13001 20281 13035 20315
rect 6101 20213 6135 20247
rect 6653 20213 6687 20247
rect 6745 20213 6779 20247
rect 11989 20213 12023 20247
rect 14197 20213 14231 20247
rect 6377 20009 6411 20043
rect 6745 20009 6779 20043
rect 12725 20009 12759 20043
rect 14381 20009 14415 20043
rect 7113 19941 7147 19975
rect 9045 19873 9079 19907
rect 11713 19873 11747 19907
rect 6553 19805 6587 19839
rect 6653 19805 6687 19839
rect 6837 19805 6871 19839
rect 7297 19805 7331 19839
rect 9303 19775 9337 19809
rect 11987 19805 12021 19839
rect 13369 19805 13403 19839
rect 14197 19805 14231 19839
rect 1501 19737 1535 19771
rect 1685 19737 1719 19771
rect 13737 19737 13771 19771
rect 10057 19669 10091 19703
rect 11345 19465 11379 19499
rect 14013 19465 14047 19499
rect 14381 19465 14415 19499
rect 5641 19329 5675 19363
rect 5833 19319 5867 19353
rect 6101 19329 6135 19363
rect 7279 19359 7313 19393
rect 8861 19329 8895 19363
rect 9505 19329 9539 19363
rect 9689 19329 9723 19363
rect 11621 19329 11655 19363
rect 11879 19359 11913 19393
rect 13093 19329 13127 19363
rect 13737 19329 13771 19363
rect 14197 19329 14231 19363
rect 7021 19261 7055 19295
rect 10149 19261 10183 19295
rect 10425 19261 10459 19295
rect 10542 19261 10576 19295
rect 10701 19261 10735 19295
rect 5917 19193 5951 19227
rect 5733 19125 5767 19159
rect 8033 19125 8067 19159
rect 8677 19125 8711 19159
rect 12633 19125 12667 19159
rect 13369 19125 13403 19159
rect 1593 18921 1627 18955
rect 10977 18921 11011 18955
rect 12173 18921 12207 18955
rect 5365 18853 5399 18887
rect 9045 18853 9079 18887
rect 13737 18853 13771 18887
rect 6009 18785 6043 18819
rect 7481 18785 7515 18819
rect 9505 18785 9539 18819
rect 9965 18785 9999 18819
rect 12357 18785 12391 18819
rect 1409 18717 1443 18751
rect 4353 18717 4387 18751
rect 4611 18687 4645 18721
rect 5733 18717 5767 18751
rect 5825 18717 5859 18751
rect 6101 18717 6135 18751
rect 6359 18717 6393 18751
rect 7755 18717 7789 18751
rect 8953 18717 8987 18751
rect 9137 18717 9171 18751
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 10239 18717 10273 18751
rect 11529 18717 11563 18751
rect 12599 18717 12633 18751
rect 13921 18717 13955 18751
rect 14289 18717 14323 18751
rect 11897 18649 11931 18683
rect 6009 18581 6043 18615
rect 7113 18581 7147 18615
rect 8493 18581 8527 18615
rect 9505 18581 9539 18615
rect 11345 18581 11379 18615
rect 13369 18581 13403 18615
rect 14105 18581 14139 18615
rect 5549 18377 5583 18411
rect 5825 18377 5859 18411
rect 10333 18377 10367 18411
rect 11345 18377 11379 18411
rect 13645 18377 13679 18411
rect 14105 18309 14139 18343
rect 14473 18309 14507 18343
rect 1501 18241 1535 18275
rect 4169 18241 4203 18275
rect 4436 18241 4470 18275
rect 5733 18241 5767 18275
rect 6193 18241 6227 18275
rect 6561 18241 6595 18275
rect 8769 18241 8803 18275
rect 9045 18241 9079 18275
rect 9689 18241 9723 18275
rect 10241 18241 10275 18275
rect 11069 18241 11103 18275
rect 11161 18241 11195 18275
rect 11803 18241 11837 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 7849 18173 7883 18207
rect 8033 18173 8067 18207
rect 8493 18173 8527 18207
rect 8907 18173 8941 18207
rect 11529 18173 11563 18207
rect 1685 18105 1719 18139
rect 6009 18105 6043 18139
rect 6377 18037 6411 18071
rect 10885 18037 10919 18071
rect 12541 18037 12575 18071
rect 13001 18037 13035 18071
rect 10241 17833 10275 17867
rect 10701 17833 10735 17867
rect 12541 17833 12575 17867
rect 13277 17833 13311 17867
rect 14381 17833 14415 17867
rect 7205 17765 7239 17799
rect 13829 17765 13863 17799
rect 10793 17697 10827 17731
rect 10425 17629 10459 17663
rect 10517 17629 10551 17663
rect 11067 17629 11101 17663
rect 12357 17629 12391 17663
rect 12633 17629 12667 17663
rect 13001 17629 13035 17663
rect 14197 17629 14231 17663
rect 5089 17561 5123 17595
rect 5917 17561 5951 17595
rect 6193 17561 6227 17595
rect 6285 17561 6319 17595
rect 6653 17561 6687 17595
rect 13553 17561 13587 17595
rect 5181 17493 5215 17527
rect 7021 17493 7055 17527
rect 11805 17493 11839 17527
rect 12817 17493 12851 17527
rect 1593 17289 1627 17323
rect 13369 17289 13403 17323
rect 14197 17289 14231 17323
rect 1501 17153 1535 17187
rect 4905 17153 4939 17187
rect 5179 17153 5213 17187
rect 6469 17153 6503 17187
rect 6743 17153 6777 17187
rect 9413 17153 9447 17187
rect 12449 17153 12483 17187
rect 12725 17153 12759 17187
rect 13553 17153 13587 17187
rect 13921 17153 13955 17187
rect 9597 17085 9631 17119
rect 10333 17085 10367 17119
rect 10471 17085 10505 17119
rect 10609 17085 10643 17119
rect 11529 17085 11563 17119
rect 11713 17085 11747 17119
rect 12173 17085 12207 17119
rect 12587 17085 12621 17119
rect 5917 17017 5951 17051
rect 10057 17017 10091 17051
rect 7481 16949 7515 16983
rect 11253 16949 11287 16983
rect 13645 16949 13679 16983
rect 6561 16745 6595 16779
rect 10425 16745 10459 16779
rect 11805 16745 11839 16779
rect 14381 16745 14415 16779
rect 1685 16677 1719 16711
rect 8125 16677 8159 16711
rect 13921 16677 13955 16711
rect 5549 16609 5583 16643
rect 7113 16609 7147 16643
rect 12265 16609 12299 16643
rect 12725 16609 12759 16643
rect 13118 16609 13152 16643
rect 13277 16609 13311 16643
rect 5791 16541 5825 16575
rect 7355 16541 7389 16575
rect 9413 16541 9447 16575
rect 9687 16541 9721 16575
rect 11989 16541 12023 16575
rect 12081 16541 12115 16575
rect 13001 16541 13035 16575
rect 14289 16541 14323 16575
rect 1501 16473 1535 16507
rect 10425 16201 10459 16235
rect 12357 16201 12391 16235
rect 14473 16201 14507 16235
rect 1685 16133 1719 16167
rect 9321 16133 9355 16167
rect 1501 16065 1535 16099
rect 7481 16065 7515 16099
rect 8401 16065 8435 16099
rect 8539 16065 8573 16099
rect 8677 16065 8711 16099
rect 9687 16065 9721 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 12817 16065 12851 16099
rect 13829 16065 13863 16099
rect 7665 15997 7699 16031
rect 9413 15997 9447 16031
rect 13277 15997 13311 16031
rect 13553 15997 13587 16031
rect 13670 15997 13704 16031
rect 8125 15929 8159 15963
rect 13277 15657 13311 15691
rect 14381 15657 14415 15691
rect 12173 15589 12207 15623
rect 12265 15521 12299 15555
rect 1409 15453 1443 15487
rect 1683 15453 1717 15487
rect 5549 15453 5583 15487
rect 5823 15453 5857 15487
rect 9505 15453 9539 15487
rect 9747 15453 9781 15487
rect 12507 15453 12541 15487
rect 13737 15453 13771 15487
rect 11989 15385 12023 15419
rect 14289 15385 14323 15419
rect 2421 15317 2455 15351
rect 6561 15317 6595 15351
rect 10517 15317 10551 15351
rect 13829 15317 13863 15351
rect 13829 15113 13863 15147
rect 11345 15045 11379 15079
rect 14289 15045 14323 15079
rect 1683 14977 1717 15011
rect 7849 14977 7883 15011
rect 7987 14977 8021 15011
rect 8125 14977 8159 15011
rect 10425 14977 10459 15011
rect 10701 14977 10735 15011
rect 12541 14977 12575 15011
rect 13059 14977 13093 15011
rect 1409 14909 1443 14943
rect 6929 14909 6963 14943
rect 7113 14909 7147 14943
rect 7573 14909 7607 14943
rect 9505 14909 9539 14943
rect 9689 14909 9723 14943
rect 10542 14909 10576 14943
rect 12817 14909 12851 14943
rect 10149 14841 10183 14875
rect 2421 14773 2455 14807
rect 8769 14773 8803 14807
rect 12725 14773 12759 14807
rect 14381 14773 14415 14807
rect 1593 14569 1627 14603
rect 7481 14569 7515 14603
rect 9965 14569 9999 14603
rect 13185 14569 13219 14603
rect 14473 14501 14507 14535
rect 13921 14433 13955 14467
rect 2237 14365 2271 14399
rect 2513 14365 2547 14399
rect 6469 14365 6503 14399
rect 6727 14335 6761 14369
rect 8953 14365 8987 14399
rect 9195 14365 9229 14399
rect 10425 14365 10459 14399
rect 10699 14365 10733 14399
rect 11805 14365 11839 14399
rect 12047 14365 12081 14399
rect 13369 14365 13403 14399
rect 13737 14365 13771 14399
rect 1501 14297 1535 14331
rect 14289 14297 14323 14331
rect 2053 14229 2087 14263
rect 2329 14229 2363 14263
rect 11437 14229 11471 14263
rect 12817 14229 12851 14263
rect 7389 14025 7423 14059
rect 9873 14025 9907 14059
rect 2421 13957 2455 13991
rect 13369 13957 13403 13991
rect 1869 13889 1903 13923
rect 6377 13889 6411 13923
rect 6651 13889 6685 13923
rect 9070 13889 9104 13923
rect 9229 13889 9263 13923
rect 10331 13889 10365 13923
rect 12725 13889 12759 13923
rect 8033 13821 8067 13855
rect 8217 13821 8251 13855
rect 8677 13821 8711 13855
rect 8953 13821 8987 13855
rect 10057 13821 10091 13855
rect 11529 13821 11563 13855
rect 11713 13821 11747 13855
rect 12173 13821 12207 13855
rect 12449 13821 12483 13855
rect 12566 13821 12600 13855
rect 13645 13821 13679 13855
rect 13921 13821 13955 13855
rect 1961 13685 1995 13719
rect 2513 13685 2547 13719
rect 11069 13685 11103 13719
rect 5733 13481 5767 13515
rect 13921 13481 13955 13515
rect 14105 13481 14139 13515
rect 4721 13345 4755 13379
rect 12725 13345 12759 13379
rect 13001 13345 13035 13379
rect 13118 13345 13152 13379
rect 1409 13277 1443 13311
rect 1683 13277 1717 13311
rect 4963 13277 4997 13311
rect 6101 13277 6135 13311
rect 6359 13247 6393 13281
rect 7481 13277 7515 13311
rect 7723 13277 7757 13311
rect 9689 13277 9723 13311
rect 9963 13277 9997 13311
rect 12081 13277 12115 13311
rect 12265 13277 12299 13311
rect 13277 13277 13311 13311
rect 14289 13277 14323 13311
rect 2421 13141 2455 13175
rect 7113 13141 7147 13175
rect 8493 13141 8527 13175
rect 10701 13141 10735 13175
rect 9413 12937 9447 12971
rect 11989 12937 12023 12971
rect 12265 12937 12299 12971
rect 13369 12937 13403 12971
rect 13921 12937 13955 12971
rect 14473 12937 14507 12971
rect 1667 12831 1701 12865
rect 8493 12801 8527 12835
rect 8610 12801 8644 12835
rect 8769 12801 8803 12835
rect 9779 12801 9813 12835
rect 11805 12801 11839 12835
rect 12081 12801 12115 12835
rect 12615 12831 12649 12865
rect 13737 12801 13771 12835
rect 14013 12801 14047 12835
rect 14289 12801 14323 12835
rect 1409 12733 1443 12767
rect 7573 12733 7607 12767
rect 7757 12733 7791 12767
rect 8217 12733 8251 12767
rect 9505 12733 9539 12767
rect 12357 12733 12391 12767
rect 2421 12597 2455 12631
rect 10517 12597 10551 12631
rect 14197 12597 14231 12631
rect 2329 12393 2363 12427
rect 13461 12393 13495 12427
rect 13921 12325 13955 12359
rect 7573 12257 7607 12291
rect 7966 12257 8000 12291
rect 11621 12257 11655 12291
rect 12265 12257 12299 12291
rect 2237 12189 2271 12223
rect 2513 12189 2547 12223
rect 6929 12189 6963 12223
rect 7113 12189 7147 12223
rect 7849 12189 7883 12223
rect 8125 12189 8159 12223
rect 11805 12189 11839 12223
rect 12541 12189 12575 12223
rect 12658 12189 12692 12223
rect 12817 12189 12851 12223
rect 13737 12189 13771 12223
rect 14289 12189 14323 12223
rect 1501 12121 1535 12155
rect 10057 12121 10091 12155
rect 10149 12121 10183 12155
rect 10517 12121 10551 12155
rect 1593 12053 1627 12087
rect 2053 12053 2087 12087
rect 8769 12053 8803 12087
rect 9781 12053 9815 12087
rect 10885 12053 10919 12087
rect 11069 12053 11103 12087
rect 14473 12053 14507 12087
rect 7757 11849 7791 11883
rect 14381 11849 14415 11883
rect 1501 11713 1535 11747
rect 6745 11713 6779 11747
rect 7019 11713 7053 11747
rect 8861 11713 8895 11747
rect 9103 11713 9137 11747
rect 12265 11713 12299 11747
rect 12725 11713 12759 11747
rect 13461 11713 13495 11747
rect 12541 11645 12575 11679
rect 13578 11645 13612 11679
rect 13737 11645 13771 11679
rect 13185 11577 13219 11611
rect 1593 11509 1627 11543
rect 9873 11509 9907 11543
rect 12449 11509 12483 11543
rect 6653 11305 6687 11339
rect 11989 11305 12023 11339
rect 13369 11305 13403 11339
rect 13921 11305 13955 11339
rect 14473 11237 14507 11271
rect 5641 11169 5675 11203
rect 5883 11101 5917 11135
rect 10977 11101 11011 11135
rect 11251 11101 11285 11135
rect 12357 11101 12391 11135
rect 12599 11101 12633 11135
rect 13737 11101 13771 11135
rect 14289 11101 14323 11135
rect 1961 10761 1995 10795
rect 13829 10761 13863 10795
rect 14473 10761 14507 10795
rect 1501 10625 1535 10659
rect 2145 10625 2179 10659
rect 4503 10625 4537 10659
rect 5917 10625 5951 10659
rect 6803 10625 6837 10659
rect 10299 10625 10333 10659
rect 11897 10625 11931 10659
rect 13059 10625 13093 10659
rect 14289 10625 14323 10659
rect 4261 10557 4295 10591
rect 6561 10557 6595 10591
rect 8217 10557 8251 10591
rect 10057 10557 10091 10591
rect 12173 10557 12207 10591
rect 12817 10557 12851 10591
rect 1593 10421 1627 10455
rect 5273 10421 5307 10455
rect 5733 10421 5767 10455
rect 7573 10421 7607 10455
rect 11069 10421 11103 10455
rect 13093 10217 13127 10251
rect 13645 10217 13679 10251
rect 13921 10217 13955 10251
rect 14381 10217 14415 10251
rect 6561 10149 6595 10183
rect 7573 10149 7607 10183
rect 5549 10081 5583 10115
rect 7113 10081 7147 10115
rect 7849 10081 7883 10115
rect 7987 10081 8021 10115
rect 9137 10081 9171 10115
rect 9321 10081 9355 10115
rect 12081 10081 12115 10115
rect 1409 10013 1443 10047
rect 1683 10013 1717 10047
rect 4997 10013 5031 10047
rect 5181 10013 5215 10047
rect 5273 10013 5307 10047
rect 5823 10013 5857 10047
rect 6929 10013 6963 10047
rect 8125 10013 8159 10047
rect 9595 10013 9629 10047
rect 10701 10013 10735 10047
rect 10975 10013 11009 10047
rect 12355 10013 12389 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 14289 9945 14323 9979
rect 2421 9877 2455 9911
rect 5181 9877 5215 9911
rect 5365 9877 5399 9911
rect 8769 9877 8803 9911
rect 10333 9877 10367 9911
rect 11713 9877 11747 9911
rect 1685 9673 1719 9707
rect 2053 9673 2087 9707
rect 5917 9673 5951 9707
rect 14473 9605 14507 9639
rect 1593 9537 1627 9571
rect 1869 9537 1903 9571
rect 2329 9537 2363 9571
rect 5089 9537 5123 9571
rect 5181 9537 5215 9571
rect 6101 9537 6135 9571
rect 8309 9537 8343 9571
rect 9689 9537 9723 9571
rect 10701 9537 10735 9571
rect 11345 9537 11379 9571
rect 11805 9537 11839 9571
rect 12081 9537 12115 9571
rect 12383 9537 12417 9571
rect 12633 9537 12667 9571
rect 13553 9537 13587 9571
rect 13829 9537 13863 9571
rect 5365 9469 5399 9503
rect 7113 9469 7147 9503
rect 7297 9469 7331 9503
rect 7757 9469 7791 9503
rect 8033 9469 8067 9503
rect 8171 9469 8205 9503
rect 9505 9469 9539 9503
rect 10425 9469 10459 9503
rect 10542 9469 10576 9503
rect 12771 9469 12805 9503
rect 13670 9469 13704 9503
rect 10149 9401 10183 9435
rect 11989 9401 12023 9435
rect 13277 9401 13311 9435
rect 2145 9333 2179 9367
rect 5273 9333 5307 9367
rect 8953 9333 8987 9367
rect 12265 9333 12299 9367
rect 12541 9333 12575 9367
rect 9597 9061 9631 9095
rect 11529 9061 11563 9095
rect 1409 8993 1443 9027
rect 9873 8993 9907 9027
rect 10149 8993 10183 9027
rect 10885 8993 10919 9027
rect 11805 8993 11839 9027
rect 1667 8895 1701 8929
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9990 8925 10024 8959
rect 11069 8925 11103 8959
rect 11943 8925 11977 8959
rect 12081 8925 12115 8959
rect 12817 8925 12851 8959
rect 13093 8925 13127 8959
rect 13369 8925 13403 8959
rect 14289 8925 14323 8959
rect 10793 8857 10827 8891
rect 12725 8857 12759 8891
rect 2421 8789 2455 8823
rect 13001 8789 13035 8823
rect 14473 8789 14507 8823
rect 6653 8585 6687 8619
rect 13369 8585 13403 8619
rect 14105 8585 14139 8619
rect 1685 8517 1719 8551
rect 2329 8449 2363 8483
rect 4905 8449 4939 8483
rect 5163 8479 5197 8513
rect 6377 8449 6411 8483
rect 6745 8449 6779 8483
rect 7021 8449 7055 8483
rect 7205 8449 7239 8483
rect 9413 8449 9447 8483
rect 10450 8449 10484 8483
rect 10609 8449 10643 8483
rect 11253 8449 11287 8483
rect 11529 8449 11563 8483
rect 12449 8449 12483 8483
rect 12566 8449 12600 8483
rect 13921 8449 13955 8483
rect 14289 8449 14323 8483
rect 6653 8381 6687 8415
rect 7113 8381 7147 8415
rect 8585 8381 8619 8415
rect 9597 8381 9631 8415
rect 10333 8381 10367 8415
rect 11713 8381 11747 8415
rect 12173 8381 12207 8415
rect 12725 8381 12759 8415
rect 1869 8313 1903 8347
rect 5917 8313 5951 8347
rect 6469 8313 6503 8347
rect 6837 8313 6871 8347
rect 10063 8313 10097 8347
rect 2145 8245 2179 8279
rect 8493 8245 8527 8279
rect 14381 8245 14415 8279
rect 1593 8041 1627 8075
rect 6377 8041 6411 8075
rect 12357 8041 12391 8075
rect 6653 7973 6687 8007
rect 14473 7973 14507 8007
rect 7113 7905 7147 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 7966 7905 8000 7939
rect 9597 7905 9631 7939
rect 10057 7905 10091 7939
rect 10333 7905 10367 7939
rect 10609 7905 10643 7939
rect 11345 7905 11379 7939
rect 13921 7905 13955 7939
rect 1501 7837 1535 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 8125 7837 8159 7871
rect 9413 7837 9447 7871
rect 10450 7837 10484 7871
rect 11619 7837 11653 7871
rect 14289 7837 14323 7871
rect 12817 7769 12851 7803
rect 13737 7769 13771 7803
rect 8769 7701 8803 7735
rect 11253 7701 11287 7735
rect 12909 7701 12943 7735
rect 1961 7497 1995 7531
rect 7573 7497 7607 7531
rect 9781 7497 9815 7531
rect 14473 7497 14507 7531
rect 1501 7429 1535 7463
rect 2145 7361 2179 7395
rect 6561 7361 6595 7395
rect 6835 7361 6869 7395
rect 8999 7361 9033 7395
rect 10057 7361 10091 7395
rect 10331 7361 10365 7395
rect 11989 7361 12023 7395
rect 12633 7361 12667 7395
rect 12817 7361 12851 7395
rect 13553 7361 13587 7395
rect 13691 7361 13725 7395
rect 7941 7293 7975 7327
rect 8125 7293 8159 7327
rect 8585 7293 8619 7327
rect 8861 7293 8895 7327
rect 9137 7293 9171 7327
rect 11713 7293 11747 7327
rect 13829 7293 13863 7327
rect 11069 7225 11103 7259
rect 13277 7225 13311 7259
rect 1593 7157 1627 7191
rect 2421 6953 2455 6987
rect 14381 6953 14415 6987
rect 9965 6817 9999 6851
rect 10425 6817 10459 6851
rect 10818 6817 10852 6851
rect 10977 6817 11011 6851
rect 1409 6749 1443 6783
rect 1683 6749 1717 6783
rect 9781 6749 9815 6783
rect 10701 6749 10735 6783
rect 12817 6749 12851 6783
rect 12909 6749 12943 6783
rect 13277 6749 13311 6783
rect 14289 6749 14323 6783
rect 12541 6681 12575 6715
rect 11621 6613 11655 6647
rect 13645 6613 13679 6647
rect 13829 6613 13863 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 12357 6409 12391 6443
rect 13645 6409 13679 6443
rect 1501 6341 1535 6375
rect 12725 6341 12759 6375
rect 13461 6341 13495 6375
rect 2237 6273 2271 6307
rect 2513 6273 2547 6307
rect 7631 6273 7665 6307
rect 8953 6273 8987 6307
rect 9689 6273 9723 6307
rect 12633 6273 12667 6307
rect 13093 6273 13127 6307
rect 14289 6273 14323 6307
rect 7389 6205 7423 6239
rect 8769 6205 8803 6239
rect 9806 6205 9840 6239
rect 9965 6205 9999 6239
rect 9413 6137 9447 6171
rect 14473 6137 14507 6171
rect 2053 6069 2087 6103
rect 8401 6069 8435 6103
rect 10609 6069 10643 6103
rect 2421 5865 2455 5899
rect 8401 5865 8435 5899
rect 13553 5865 13587 5899
rect 14381 5865 14415 5899
rect 13921 5797 13955 5831
rect 7389 5729 7423 5763
rect 9781 5729 9815 5763
rect 9965 5729 9999 5763
rect 10425 5729 10459 5763
rect 10701 5729 10735 5763
rect 10977 5729 11011 5763
rect 11897 5729 11931 5763
rect 12357 5729 12391 5763
rect 12633 5729 12667 5763
rect 12750 5729 12784 5763
rect 1409 5661 1443 5695
rect 1667 5631 1701 5665
rect 7631 5661 7665 5695
rect 10839 5661 10873 5695
rect 11713 5661 11747 5695
rect 12909 5661 12943 5695
rect 13737 5661 13771 5695
rect 14289 5593 14323 5627
rect 11621 5525 11655 5559
rect 9045 5321 9079 5355
rect 12173 5321 12207 5355
rect 13277 5321 13311 5355
rect 1685 5253 1719 5287
rect 2237 5253 2271 5287
rect 2145 5185 2179 5219
rect 8033 5185 8067 5219
rect 8291 5215 8325 5249
rect 11989 5185 12023 5219
rect 12507 5185 12541 5219
rect 13645 5185 13679 5219
rect 13921 5185 13955 5219
rect 12253 5117 12287 5151
rect 1777 4981 1811 5015
rect 1593 4777 1627 4811
rect 10885 4777 10919 4811
rect 12265 4777 12299 4811
rect 13645 4777 13679 4811
rect 14381 4777 14415 4811
rect 9873 4641 9907 4675
rect 11253 4641 11287 4675
rect 12633 4641 12667 4675
rect 1501 4573 1535 4607
rect 10115 4573 10149 4607
rect 11495 4573 11529 4607
rect 12891 4543 12925 4577
rect 14289 4573 14323 4607
rect 1409 4097 1443 4131
rect 8767 4097 8801 4131
rect 11863 4097 11897 4131
rect 13259 4127 13293 4161
rect 8493 4029 8527 4063
rect 11621 4029 11655 4063
rect 13001 4029 13035 4063
rect 9505 3961 9539 3995
rect 1593 3893 1627 3927
rect 12633 3893 12667 3927
rect 14013 3893 14047 3927
rect 13093 3689 13127 3723
rect 14381 3689 14415 3723
rect 12081 3553 12115 3587
rect 12323 3485 12357 3519
rect 14289 3485 14323 3519
rect 4445 2601 4479 2635
rect 4353 2329 4387 2363
rect 4077 2057 4111 2091
rect 5089 2057 5123 2091
rect 5825 2057 5859 2091
rect 6561 2057 6595 2091
rect 7205 2057 7239 2091
rect 7941 2057 7975 2091
rect 8677 2057 8711 2091
rect 10885 2057 10919 2091
rect 12357 2057 12391 2091
rect 13093 2057 13127 2091
rect 14197 2057 14231 2091
rect 14105 1989 14139 2023
rect 2145 1921 2179 1955
rect 4261 1921 4295 1955
rect 4997 1921 5031 1955
rect 5733 1921 5767 1955
rect 6469 1921 6503 1955
rect 7113 1921 7147 1955
rect 7849 1921 7883 1955
rect 8585 1921 8619 1955
rect 9321 1921 9355 1955
rect 10057 1921 10091 1955
rect 10793 1921 10827 1955
rect 11621 1921 11655 1955
rect 12265 1921 12299 1955
rect 13001 1921 13035 1955
rect 13737 1921 13771 1955
rect 13921 1921 13955 1955
rect 2973 1853 3007 1887
rect 10241 1785 10275 1819
rect 9413 1717 9447 1751
rect 11713 1717 11747 1751
rect 4353 1513 4387 1547
rect 5089 1513 5123 1547
rect 5825 1513 5859 1547
rect 6561 1513 6595 1547
rect 7297 1513 7331 1547
rect 8033 1513 8067 1547
rect 8953 1513 8987 1547
rect 9505 1513 9539 1547
rect 10241 1513 10275 1547
rect 10977 1513 11011 1547
rect 11713 1513 11747 1547
rect 12449 1513 12483 1547
rect 13185 1513 13219 1547
rect 13461 1513 13495 1547
rect 13737 1513 13771 1547
rect 1409 1309 1443 1343
rect 2697 1309 2731 1343
rect 3801 1309 3835 1343
rect 4537 1309 4571 1343
rect 5273 1309 5307 1343
rect 6009 1309 6043 1343
rect 6745 1309 6779 1343
rect 7481 1309 7515 1343
rect 8217 1309 8251 1343
rect 9137 1309 9171 1343
rect 9689 1309 9723 1343
rect 10425 1309 10459 1343
rect 11161 1309 11195 1343
rect 11897 1309 11931 1343
rect 12633 1309 12667 1343
rect 13093 1309 13127 1343
rect 13369 1309 13403 1343
rect 13645 1309 13679 1343
rect 13921 1309 13955 1343
rect 2237 1241 2271 1275
rect 3433 1241 3467 1275
rect 4077 1241 4111 1275
rect 14197 1241 14231 1275
rect 14381 1241 14415 1275
rect 12909 1173 12943 1207
<< metal1 >>
rect 1104 43546 14971 43568
rect 1104 43494 4376 43546
rect 4428 43494 4440 43546
rect 4492 43494 4504 43546
rect 4556 43494 4568 43546
rect 4620 43494 4632 43546
rect 4684 43494 7803 43546
rect 7855 43494 7867 43546
rect 7919 43494 7931 43546
rect 7983 43494 7995 43546
rect 8047 43494 8059 43546
rect 8111 43494 11230 43546
rect 11282 43494 11294 43546
rect 11346 43494 11358 43546
rect 11410 43494 11422 43546
rect 11474 43494 11486 43546
rect 11538 43494 14657 43546
rect 14709 43494 14721 43546
rect 14773 43494 14785 43546
rect 14837 43494 14849 43546
rect 14901 43494 14913 43546
rect 14965 43494 14971 43546
rect 1104 43472 14971 43494
rect 566 43392 572 43444
rect 624 43432 630 43444
rect 2685 43435 2743 43441
rect 2685 43432 2697 43435
rect 624 43404 2697 43432
rect 624 43392 630 43404
rect 2685 43401 2697 43404
rect 2731 43401 2743 43435
rect 2685 43395 2743 43401
rect 2774 43392 2780 43444
rect 2832 43432 2838 43444
rect 3053 43435 3111 43441
rect 3053 43432 3065 43435
rect 2832 43404 3065 43432
rect 2832 43392 2838 43404
rect 3053 43401 3065 43404
rect 3099 43401 3111 43435
rect 3053 43395 3111 43401
rect 3510 43392 3516 43444
rect 3568 43432 3574 43444
rect 3973 43435 4031 43441
rect 3973 43432 3985 43435
rect 3568 43404 3985 43432
rect 3568 43392 3574 43404
rect 3973 43401 3985 43404
rect 4019 43401 4031 43435
rect 3973 43395 4031 43401
rect 4246 43392 4252 43444
rect 4304 43432 4310 43444
rect 4525 43435 4583 43441
rect 4525 43432 4537 43435
rect 4304 43404 4537 43432
rect 4304 43392 4310 43404
rect 4525 43401 4537 43404
rect 4571 43401 4583 43435
rect 4525 43395 4583 43401
rect 4982 43392 4988 43444
rect 5040 43432 5046 43444
rect 5261 43435 5319 43441
rect 5261 43432 5273 43435
rect 5040 43404 5273 43432
rect 5040 43392 5046 43404
rect 5261 43401 5273 43404
rect 5307 43401 5319 43435
rect 5261 43395 5319 43401
rect 5718 43392 5724 43444
rect 5776 43432 5782 43444
rect 5997 43435 6055 43441
rect 5997 43432 6009 43435
rect 5776 43404 6009 43432
rect 5776 43392 5782 43404
rect 5997 43401 6009 43404
rect 6043 43401 6055 43435
rect 5997 43395 6055 43401
rect 6454 43392 6460 43444
rect 6512 43432 6518 43444
rect 6733 43435 6791 43441
rect 6733 43432 6745 43435
rect 6512 43404 6745 43432
rect 6512 43392 6518 43404
rect 6733 43401 6745 43404
rect 6779 43401 6791 43435
rect 6733 43395 6791 43401
rect 7190 43392 7196 43444
rect 7248 43432 7254 43444
rect 7469 43435 7527 43441
rect 7469 43432 7481 43435
rect 7248 43404 7481 43432
rect 7248 43392 7254 43404
rect 7469 43401 7481 43404
rect 7515 43401 7527 43435
rect 7469 43395 7527 43401
rect 8202 43392 8208 43444
rect 8260 43392 8266 43444
rect 8662 43392 8668 43444
rect 8720 43432 8726 43444
rect 9125 43435 9183 43441
rect 9125 43432 9137 43435
rect 8720 43404 9137 43432
rect 8720 43392 8726 43404
rect 9125 43401 9137 43404
rect 9171 43401 9183 43435
rect 9125 43395 9183 43401
rect 9398 43392 9404 43444
rect 9456 43432 9462 43444
rect 9677 43435 9735 43441
rect 9677 43432 9689 43435
rect 9456 43404 9689 43432
rect 9456 43392 9462 43404
rect 9677 43401 9689 43404
rect 9723 43401 9735 43435
rect 9677 43395 9735 43401
rect 10134 43392 10140 43444
rect 10192 43432 10198 43444
rect 10413 43435 10471 43441
rect 10413 43432 10425 43435
rect 10192 43404 10425 43432
rect 10192 43392 10198 43404
rect 10413 43401 10425 43404
rect 10459 43401 10471 43435
rect 10413 43395 10471 43401
rect 10870 43392 10876 43444
rect 10928 43432 10934 43444
rect 11701 43435 11759 43441
rect 11701 43432 11713 43435
rect 10928 43404 11713 43432
rect 10928 43392 10934 43404
rect 11701 43401 11713 43404
rect 11747 43401 11759 43435
rect 11701 43395 11759 43401
rect 12342 43392 12348 43444
rect 12400 43432 12406 43444
rect 12621 43435 12679 43441
rect 12621 43432 12633 43435
rect 12400 43404 12633 43432
rect 12400 43392 12406 43404
rect 12621 43401 12633 43404
rect 12667 43401 12679 43435
rect 12621 43395 12679 43401
rect 13078 43392 13084 43444
rect 13136 43432 13142 43444
rect 13357 43435 13415 43441
rect 13357 43432 13369 43435
rect 13136 43404 13369 43432
rect 13136 43392 13142 43404
rect 13357 43401 13369 43404
rect 13403 43401 13415 43435
rect 13357 43395 13415 43401
rect 13814 43392 13820 43444
rect 13872 43432 13878 43444
rect 14277 43435 14335 43441
rect 14277 43432 14289 43435
rect 13872 43404 14289 43432
rect 13872 43392 13878 43404
rect 14277 43401 14289 43404
rect 14323 43401 14335 43435
rect 14277 43395 14335 43401
rect 1489 43299 1547 43305
rect 1489 43265 1501 43299
rect 1535 43296 1547 43299
rect 1762 43296 1768 43308
rect 1535 43268 1768 43296
rect 1535 43265 1547 43268
rect 1489 43259 1547 43265
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 2130 43256 2136 43308
rect 2188 43256 2194 43308
rect 2498 43256 2504 43308
rect 2556 43256 2562 43308
rect 2961 43299 3019 43305
rect 2961 43265 2973 43299
rect 3007 43296 3019 43299
rect 3050 43296 3056 43308
rect 3007 43268 3056 43296
rect 3007 43265 3019 43268
rect 2961 43259 3019 43265
rect 3050 43256 3056 43268
rect 3108 43256 3114 43308
rect 3786 43256 3792 43308
rect 3844 43256 3850 43308
rect 4338 43256 4344 43308
rect 4396 43256 4402 43308
rect 5074 43256 5080 43308
rect 5132 43256 5138 43308
rect 5810 43256 5816 43308
rect 5868 43256 5874 43308
rect 6546 43256 6552 43308
rect 6604 43256 6610 43308
rect 7282 43256 7288 43308
rect 7340 43256 7346 43308
rect 8018 43256 8024 43308
rect 8076 43256 8082 43308
rect 8938 43256 8944 43308
rect 8996 43256 9002 43308
rect 9306 43256 9312 43308
rect 9364 43296 9370 43308
rect 9585 43299 9643 43305
rect 9585 43296 9597 43299
rect 9364 43268 9597 43296
rect 9364 43256 9370 43268
rect 9585 43265 9597 43268
rect 9631 43265 9643 43299
rect 9585 43259 9643 43265
rect 10226 43256 10232 43308
rect 10284 43256 10290 43308
rect 11606 43256 11612 43308
rect 11664 43256 11670 43308
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 12526 43256 12532 43308
rect 12584 43256 12590 43308
rect 13173 43299 13231 43305
rect 13173 43265 13185 43299
rect 13219 43296 13231 43299
rect 13262 43296 13268 43308
rect 13219 43268 13268 43296
rect 13219 43265 13231 43268
rect 13173 43259 13231 43265
rect 13262 43256 13268 43268
rect 13320 43256 13326 43308
rect 13630 43256 13636 43308
rect 13688 43256 13694 43308
rect 14090 43256 14096 43308
rect 14148 43256 14154 43308
rect 14550 43188 14556 43240
rect 14608 43188 14614 43240
rect 2038 43120 2044 43172
rect 2096 43160 2102 43172
rect 2317 43163 2375 43169
rect 2317 43160 2329 43163
rect 2096 43132 2329 43160
rect 2096 43120 2102 43132
rect 2317 43129 2329 43132
rect 2363 43129 2375 43163
rect 2317 43123 2375 43129
rect 13817 43163 13875 43169
rect 13817 43129 13829 43163
rect 13863 43160 13875 43163
rect 14568 43160 14596 43188
rect 13863 43132 14596 43160
rect 13863 43129 13875 43132
rect 13817 43123 13875 43129
rect 1394 43052 1400 43104
rect 1452 43092 1458 43104
rect 1581 43095 1639 43101
rect 1581 43092 1593 43095
rect 1452 43064 1593 43092
rect 1452 43052 1458 43064
rect 1581 43061 1593 43064
rect 1627 43061 1639 43095
rect 1581 43055 1639 43061
rect 11698 43052 11704 43104
rect 11756 43092 11762 43104
rect 12253 43095 12311 43101
rect 12253 43092 12265 43095
rect 11756 43064 12265 43092
rect 11756 43052 11762 43064
rect 12253 43061 12265 43064
rect 12299 43061 12311 43095
rect 12253 43055 12311 43061
rect 1104 43002 14812 43024
rect 1104 42950 2663 43002
rect 2715 42950 2727 43002
rect 2779 42950 2791 43002
rect 2843 42950 2855 43002
rect 2907 42950 2919 43002
rect 2971 42950 6090 43002
rect 6142 42950 6154 43002
rect 6206 42950 6218 43002
rect 6270 42950 6282 43002
rect 6334 42950 6346 43002
rect 6398 42950 9517 43002
rect 9569 42950 9581 43002
rect 9633 42950 9645 43002
rect 9697 42950 9709 43002
rect 9761 42950 9773 43002
rect 9825 42950 12944 43002
rect 12996 42950 13008 43002
rect 13060 42950 13072 43002
rect 13124 42950 13136 43002
rect 13188 42950 13200 43002
rect 13252 42950 14812 43002
rect 1104 42928 14812 42950
rect 2041 42891 2099 42897
rect 2041 42857 2053 42891
rect 2087 42888 2099 42891
rect 2130 42888 2136 42900
rect 2087 42860 2136 42888
rect 2087 42857 2099 42860
rect 2041 42851 2099 42857
rect 2130 42848 2136 42860
rect 2188 42848 2194 42900
rect 2777 42891 2835 42897
rect 2777 42857 2789 42891
rect 2823 42888 2835 42891
rect 3050 42888 3056 42900
rect 2823 42860 3056 42888
rect 2823 42857 2835 42860
rect 2777 42851 2835 42857
rect 3050 42848 3056 42860
rect 3108 42848 3114 42900
rect 3329 42891 3387 42897
rect 3329 42857 3341 42891
rect 3375 42888 3387 42891
rect 3786 42888 3792 42900
rect 3375 42860 3792 42888
rect 3375 42857 3387 42860
rect 3329 42851 3387 42857
rect 3786 42848 3792 42860
rect 3844 42848 3850 42900
rect 4157 42891 4215 42897
rect 4157 42857 4169 42891
rect 4203 42888 4215 42891
rect 4338 42888 4344 42900
rect 4203 42860 4344 42888
rect 4203 42857 4215 42860
rect 4157 42851 4215 42857
rect 4338 42848 4344 42860
rect 4396 42848 4402 42900
rect 5721 42891 5779 42897
rect 5721 42857 5733 42891
rect 5767 42888 5779 42891
rect 5810 42888 5816 42900
rect 5767 42860 5816 42888
rect 5767 42857 5779 42860
rect 5721 42851 5779 42857
rect 5810 42848 5816 42860
rect 5868 42848 5874 42900
rect 6457 42891 6515 42897
rect 6457 42857 6469 42891
rect 6503 42888 6515 42891
rect 6546 42888 6552 42900
rect 6503 42860 6552 42888
rect 6503 42857 6515 42860
rect 6457 42851 6515 42857
rect 6546 42848 6552 42860
rect 6604 42848 6610 42900
rect 7101 42891 7159 42897
rect 7101 42857 7113 42891
rect 7147 42888 7159 42891
rect 7282 42888 7288 42900
rect 7147 42860 7288 42888
rect 7147 42857 7159 42860
rect 7101 42851 7159 42857
rect 7282 42848 7288 42860
rect 7340 42848 7346 42900
rect 7837 42891 7895 42897
rect 7837 42857 7849 42891
rect 7883 42888 7895 42891
rect 8018 42888 8024 42900
rect 7883 42860 8024 42888
rect 7883 42857 7895 42860
rect 7837 42851 7895 42857
rect 8018 42848 8024 42860
rect 8076 42848 8082 42900
rect 8573 42891 8631 42897
rect 8573 42857 8585 42891
rect 8619 42888 8631 42891
rect 8938 42888 8944 42900
rect 8619 42860 8944 42888
rect 8619 42857 8631 42860
rect 8573 42851 8631 42857
rect 8938 42848 8944 42860
rect 8996 42848 9002 42900
rect 9306 42848 9312 42900
rect 9364 42848 9370 42900
rect 10045 42891 10103 42897
rect 10045 42857 10057 42891
rect 10091 42888 10103 42891
rect 10226 42888 10232 42900
rect 10091 42860 10232 42888
rect 10091 42857 10103 42860
rect 10045 42851 10103 42857
rect 10226 42848 10232 42860
rect 10284 42848 10290 42900
rect 10781 42891 10839 42897
rect 10781 42857 10793 42891
rect 10827 42888 10839 42891
rect 11606 42888 11612 42900
rect 10827 42860 11612 42888
rect 10827 42857 10839 42860
rect 10781 42851 10839 42857
rect 11606 42848 11612 42860
rect 11664 42848 11670 42900
rect 12066 42848 12072 42900
rect 12124 42848 12130 42900
rect 12253 42891 12311 42897
rect 12253 42857 12265 42891
rect 12299 42888 12311 42891
rect 12526 42888 12532 42900
rect 12299 42860 12532 42888
rect 12299 42857 12311 42860
rect 12253 42851 12311 42857
rect 12526 42848 12532 42860
rect 12584 42848 12590 42900
rect 12989 42891 13047 42897
rect 12989 42857 13001 42891
rect 13035 42888 13047 42891
rect 13262 42888 13268 42900
rect 13035 42860 13268 42888
rect 13035 42857 13047 42860
rect 12989 42851 13047 42857
rect 13262 42848 13268 42860
rect 13320 42848 13326 42900
rect 13630 42848 13636 42900
rect 13688 42848 13694 42900
rect 14090 42848 14096 42900
rect 14148 42888 14154 42900
rect 14277 42891 14335 42897
rect 14277 42888 14289 42891
rect 14148 42860 14289 42888
rect 14148 42848 14154 42860
rect 14277 42857 14289 42860
rect 14323 42857 14335 42891
rect 14277 42851 14335 42857
rect 11517 42823 11575 42829
rect 11517 42789 11529 42823
rect 11563 42820 11575 42823
rect 12084 42820 12112 42848
rect 11563 42792 12112 42820
rect 12713 42823 12771 42829
rect 11563 42789 11575 42792
rect 11517 42783 11575 42789
rect 12713 42789 12725 42823
rect 12759 42820 12771 42823
rect 13648 42820 13676 42848
rect 12759 42792 13676 42820
rect 12759 42789 12771 42792
rect 12713 42783 12771 42789
rect 13817 42755 13875 42761
rect 13817 42721 13829 42755
rect 13863 42752 13875 42755
rect 15286 42752 15292 42764
rect 13863 42724 15292 42752
rect 13863 42721 13875 42724
rect 13817 42715 13875 42721
rect 15286 42712 15292 42724
rect 15344 42712 15350 42764
rect 2222 42644 2228 42696
rect 2280 42644 2286 42696
rect 2958 42644 2964 42696
rect 3016 42644 3022 42696
rect 3510 42644 3516 42696
rect 3568 42644 3574 42696
rect 4341 42687 4399 42693
rect 4341 42653 4353 42687
rect 4387 42653 4399 42687
rect 4341 42647 4399 42653
rect 1210 42576 1216 42628
rect 1268 42616 1274 42628
rect 4356 42616 4384 42647
rect 5902 42644 5908 42696
rect 5960 42644 5966 42696
rect 6638 42644 6644 42696
rect 6696 42644 6702 42696
rect 7282 42644 7288 42696
rect 7340 42644 7346 42696
rect 8021 42687 8079 42693
rect 8021 42653 8033 42687
rect 8067 42684 8079 42687
rect 8202 42684 8208 42696
rect 8067 42656 8208 42684
rect 8067 42653 8079 42656
rect 8021 42647 8079 42653
rect 8202 42644 8208 42656
rect 8260 42644 8266 42696
rect 8754 42644 8760 42696
rect 8812 42644 8818 42696
rect 9490 42644 9496 42696
rect 9548 42644 9554 42696
rect 10226 42644 10232 42696
rect 10284 42644 10290 42696
rect 10962 42644 10968 42696
rect 11020 42644 11026 42696
rect 11698 42644 11704 42696
rect 11756 42644 11762 42696
rect 12434 42644 12440 42696
rect 12492 42644 12498 42696
rect 12897 42687 12955 42693
rect 12897 42653 12909 42687
rect 12943 42653 12955 42687
rect 12897 42647 12955 42653
rect 1268 42588 4384 42616
rect 1268 42576 1274 42588
rect 12912 42548 12940 42647
rect 13170 42644 13176 42696
rect 13228 42644 13234 42696
rect 14090 42644 14096 42696
rect 14148 42684 14154 42696
rect 14461 42687 14519 42693
rect 14461 42684 14473 42687
rect 14148 42656 14473 42684
rect 14148 42644 14154 42656
rect 14461 42653 14473 42656
rect 14507 42653 14519 42687
rect 14461 42647 14519 42653
rect 13538 42576 13544 42628
rect 13596 42576 13602 42628
rect 14274 42548 14280 42560
rect 12912 42520 14280 42548
rect 14274 42508 14280 42520
rect 14332 42508 14338 42560
rect 1104 42458 14971 42480
rect 1104 42406 4376 42458
rect 4428 42406 4440 42458
rect 4492 42406 4504 42458
rect 4556 42406 4568 42458
rect 4620 42406 4632 42458
rect 4684 42406 7803 42458
rect 7855 42406 7867 42458
rect 7919 42406 7931 42458
rect 7983 42406 7995 42458
rect 8047 42406 8059 42458
rect 8111 42406 11230 42458
rect 11282 42406 11294 42458
rect 11346 42406 11358 42458
rect 11410 42406 11422 42458
rect 11474 42406 11486 42458
rect 11538 42406 14657 42458
rect 14709 42406 14721 42458
rect 14773 42406 14785 42458
rect 14837 42406 14849 42458
rect 14901 42406 14913 42458
rect 14965 42406 14971 42458
rect 1104 42384 14971 42406
rect 2041 42347 2099 42353
rect 2041 42313 2053 42347
rect 2087 42344 2099 42347
rect 2222 42344 2228 42356
rect 2087 42316 2228 42344
rect 2087 42313 2099 42316
rect 2041 42307 2099 42313
rect 2222 42304 2228 42316
rect 2280 42304 2286 42356
rect 2869 42347 2927 42353
rect 2869 42313 2881 42347
rect 2915 42344 2927 42347
rect 2958 42344 2964 42356
rect 2915 42316 2964 42344
rect 2915 42313 2927 42316
rect 2869 42307 2927 42313
rect 2958 42304 2964 42316
rect 3016 42304 3022 42356
rect 5537 42347 5595 42353
rect 5537 42313 5549 42347
rect 5583 42344 5595 42347
rect 5902 42344 5908 42356
rect 5583 42316 5908 42344
rect 5583 42313 5595 42316
rect 5537 42307 5595 42313
rect 5902 42304 5908 42316
rect 5960 42304 5966 42356
rect 6365 42347 6423 42353
rect 6365 42313 6377 42347
rect 6411 42344 6423 42347
rect 6638 42344 6644 42356
rect 6411 42316 6644 42344
rect 6411 42313 6423 42316
rect 6365 42307 6423 42313
rect 6638 42304 6644 42316
rect 6696 42304 6702 42356
rect 7101 42347 7159 42353
rect 7101 42313 7113 42347
rect 7147 42344 7159 42347
rect 7282 42344 7288 42356
rect 7147 42316 7288 42344
rect 7147 42313 7159 42316
rect 7101 42307 7159 42313
rect 7282 42304 7288 42316
rect 7340 42304 7346 42356
rect 7929 42347 7987 42353
rect 7929 42313 7941 42347
rect 7975 42344 7987 42347
rect 8202 42344 8208 42356
rect 7975 42316 8208 42344
rect 7975 42313 7987 42316
rect 7929 42307 7987 42313
rect 8202 42304 8208 42316
rect 8260 42304 8266 42356
rect 8665 42347 8723 42353
rect 8665 42313 8677 42347
rect 8711 42344 8723 42347
rect 8754 42344 8760 42356
rect 8711 42316 8760 42344
rect 8711 42313 8723 42316
rect 8665 42307 8723 42313
rect 8754 42304 8760 42316
rect 8812 42304 8818 42356
rect 9309 42347 9367 42353
rect 9309 42313 9321 42347
rect 9355 42344 9367 42347
rect 9490 42344 9496 42356
rect 9355 42316 9496 42344
rect 9355 42313 9367 42316
rect 9309 42307 9367 42313
rect 9490 42304 9496 42316
rect 9548 42304 9554 42356
rect 10137 42347 10195 42353
rect 10137 42313 10149 42347
rect 10183 42344 10195 42347
rect 10226 42344 10232 42356
rect 10183 42316 10232 42344
rect 10183 42313 10195 42316
rect 10137 42307 10195 42313
rect 10226 42304 10232 42316
rect 10284 42304 10290 42356
rect 10781 42347 10839 42353
rect 10781 42313 10793 42347
rect 10827 42344 10839 42347
rect 10962 42344 10968 42356
rect 10827 42316 10968 42344
rect 10827 42313 10839 42316
rect 10781 42307 10839 42313
rect 10962 42304 10968 42316
rect 11020 42304 11026 42356
rect 11517 42347 11575 42353
rect 11517 42313 11529 42347
rect 11563 42344 11575 42347
rect 11698 42344 11704 42356
rect 11563 42316 11704 42344
rect 11563 42313 11575 42316
rect 11517 42307 11575 42313
rect 11698 42304 11704 42316
rect 11756 42304 11762 42356
rect 12253 42347 12311 42353
rect 12253 42313 12265 42347
rect 12299 42344 12311 42347
rect 12434 42344 12440 42356
rect 12299 42316 12440 42344
rect 12299 42313 12311 42316
rect 12253 42307 12311 42313
rect 12434 42304 12440 42316
rect 12492 42304 12498 42356
rect 12897 42347 12955 42353
rect 12897 42313 12909 42347
rect 12943 42344 12955 42347
rect 13170 42344 13176 42356
rect 12943 42316 13176 42344
rect 12943 42313 12955 42316
rect 12897 42307 12955 42313
rect 13170 42304 13176 42316
rect 13228 42304 13234 42356
rect 13538 42304 13544 42356
rect 13596 42344 13602 42356
rect 14001 42347 14059 42353
rect 14001 42344 14013 42347
rect 13596 42316 14013 42344
rect 13596 42304 13602 42316
rect 14001 42313 14013 42316
rect 14047 42313 14059 42347
rect 14001 42307 14059 42313
rect 14274 42304 14280 42356
rect 14332 42304 14338 42356
rect 2406 42236 2412 42288
rect 2464 42276 2470 42288
rect 2464 42248 9536 42276
rect 2464 42236 2470 42248
rect 2222 42168 2228 42220
rect 2280 42168 2286 42220
rect 3050 42168 3056 42220
rect 3108 42168 3114 42220
rect 5718 42168 5724 42220
rect 5776 42168 5782 42220
rect 6546 42168 6552 42220
rect 6604 42168 6610 42220
rect 7282 42168 7288 42220
rect 7340 42168 7346 42220
rect 8110 42168 8116 42220
rect 8168 42168 8174 42220
rect 9508 42217 9536 42248
rect 14090 42236 14096 42288
rect 14148 42236 14154 42288
rect 8849 42211 8907 42217
rect 8849 42177 8861 42211
rect 8895 42177 8907 42211
rect 8849 42171 8907 42177
rect 9493 42211 9551 42217
rect 9493 42177 9505 42211
rect 9539 42177 9551 42211
rect 9493 42171 9551 42177
rect 10321 42211 10379 42217
rect 10321 42177 10333 42211
rect 10367 42177 10379 42211
rect 10321 42171 10379 42177
rect 3602 42100 3608 42152
rect 3660 42140 3666 42152
rect 8864 42140 8892 42171
rect 3660 42112 8892 42140
rect 3660 42100 3666 42112
rect 3234 42032 3240 42084
rect 3292 42072 3298 42084
rect 10336 42072 10364 42171
rect 10962 42168 10968 42220
rect 11020 42168 11026 42220
rect 11698 42168 11704 42220
rect 11756 42168 11762 42220
rect 12434 42168 12440 42220
rect 12492 42168 12498 42220
rect 13081 42211 13139 42217
rect 13081 42177 13093 42211
rect 13127 42177 13139 42211
rect 13081 42171 13139 42177
rect 13449 42211 13507 42217
rect 13449 42177 13461 42211
rect 13495 42208 13507 42211
rect 13909 42211 13967 42217
rect 13909 42208 13921 42211
rect 13495 42180 13921 42208
rect 13495 42177 13507 42180
rect 13449 42171 13507 42177
rect 13909 42177 13921 42180
rect 13955 42208 13967 42211
rect 13998 42208 14004 42220
rect 13955 42180 14004 42208
rect 13955 42177 13967 42180
rect 13909 42171 13967 42177
rect 3292 42044 10364 42072
rect 3292 42032 3298 42044
rect 13096 42004 13124 42171
rect 13998 42168 14004 42180
rect 14056 42168 14062 42220
rect 13725 42075 13783 42081
rect 13725 42041 13737 42075
rect 13771 42072 13783 42075
rect 14108 42072 14136 42236
rect 14182 42168 14188 42220
rect 14240 42168 14246 42220
rect 14461 42211 14519 42217
rect 14461 42177 14473 42211
rect 14507 42208 14519 42211
rect 15746 42208 15752 42220
rect 14507 42180 15752 42208
rect 14507 42177 14519 42180
rect 14461 42171 14519 42177
rect 15746 42168 15752 42180
rect 15804 42168 15810 42220
rect 13771 42044 14136 42072
rect 13771 42041 13783 42044
rect 13725 42035 13783 42041
rect 15102 42004 15108 42016
rect 13096 41976 15108 42004
rect 15102 41964 15108 41976
rect 15160 41964 15166 42016
rect 1104 41914 14812 41936
rect 1104 41862 2663 41914
rect 2715 41862 2727 41914
rect 2779 41862 2791 41914
rect 2843 41862 2855 41914
rect 2907 41862 2919 41914
rect 2971 41862 6090 41914
rect 6142 41862 6154 41914
rect 6206 41862 6218 41914
rect 6270 41862 6282 41914
rect 6334 41862 6346 41914
rect 6398 41862 9517 41914
rect 9569 41862 9581 41914
rect 9633 41862 9645 41914
rect 9697 41862 9709 41914
rect 9761 41862 9773 41914
rect 9825 41862 12944 41914
rect 12996 41862 13008 41914
rect 13060 41862 13072 41914
rect 13124 41862 13136 41914
rect 13188 41862 13200 41914
rect 13252 41862 14812 41914
rect 1104 41840 14812 41862
rect 2869 41803 2927 41809
rect 2869 41769 2881 41803
rect 2915 41800 2927 41803
rect 3050 41800 3056 41812
rect 2915 41772 3056 41800
rect 2915 41769 2927 41772
rect 2869 41763 2927 41769
rect 3050 41760 3056 41772
rect 3108 41760 3114 41812
rect 14182 41760 14188 41812
rect 14240 41800 14246 41812
rect 14277 41803 14335 41809
rect 14277 41800 14289 41803
rect 14240 41772 14289 41800
rect 14240 41760 14246 41772
rect 14277 41769 14289 41772
rect 14323 41769 14335 41803
rect 14277 41763 14335 41769
rect 13998 41624 14004 41676
rect 14056 41664 14062 41676
rect 15010 41664 15016 41676
rect 14056 41636 15016 41664
rect 14056 41624 14062 41636
rect 15010 41624 15016 41636
rect 15068 41624 15074 41676
rect 3053 41599 3111 41605
rect 3053 41565 3065 41599
rect 3099 41596 3111 41599
rect 6914 41596 6920 41608
rect 3099 41568 6920 41596
rect 3099 41565 3111 41568
rect 3053 41559 3111 41565
rect 6914 41556 6920 41568
rect 6972 41556 6978 41608
rect 14461 41599 14519 41605
rect 14461 41565 14473 41599
rect 14507 41596 14519 41599
rect 15470 41596 15476 41608
rect 14507 41568 15476 41596
rect 14507 41565 14519 41568
rect 14461 41559 14519 41565
rect 15470 41556 15476 41568
rect 15528 41556 15534 41608
rect 1104 41370 14971 41392
rect 1104 41318 4376 41370
rect 4428 41318 4440 41370
rect 4492 41318 4504 41370
rect 4556 41318 4568 41370
rect 4620 41318 4632 41370
rect 4684 41318 7803 41370
rect 7855 41318 7867 41370
rect 7919 41318 7931 41370
rect 7983 41318 7995 41370
rect 8047 41318 8059 41370
rect 8111 41318 11230 41370
rect 11282 41318 11294 41370
rect 11346 41318 11358 41370
rect 11410 41318 11422 41370
rect 11474 41318 11486 41370
rect 11538 41318 14657 41370
rect 14709 41318 14721 41370
rect 14773 41318 14785 41370
rect 14837 41318 14849 41370
rect 14901 41318 14913 41370
rect 14965 41318 14971 41370
rect 1104 41296 14971 41318
rect 750 41080 756 41132
rect 808 41120 814 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 808 41092 1409 41120
rect 808 41080 814 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 8202 40916 8208 40928
rect 1627 40888 8208 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 8202 40876 8208 40888
rect 8260 40876 8266 40928
rect 1104 40826 14812 40848
rect 1104 40774 2663 40826
rect 2715 40774 2727 40826
rect 2779 40774 2791 40826
rect 2843 40774 2855 40826
rect 2907 40774 2919 40826
rect 2971 40774 6090 40826
rect 6142 40774 6154 40826
rect 6206 40774 6218 40826
rect 6270 40774 6282 40826
rect 6334 40774 6346 40826
rect 6398 40774 9517 40826
rect 9569 40774 9581 40826
rect 9633 40774 9645 40826
rect 9697 40774 9709 40826
rect 9761 40774 9773 40826
rect 9825 40774 12944 40826
rect 12996 40774 13008 40826
rect 13060 40774 13072 40826
rect 13124 40774 13136 40826
rect 13188 40774 13200 40826
rect 13252 40774 14812 40826
rect 1104 40752 14812 40774
rect 1104 40282 14971 40304
rect 1104 40230 4376 40282
rect 4428 40230 4440 40282
rect 4492 40230 4504 40282
rect 4556 40230 4568 40282
rect 4620 40230 4632 40282
rect 4684 40230 7803 40282
rect 7855 40230 7867 40282
rect 7919 40230 7931 40282
rect 7983 40230 7995 40282
rect 8047 40230 8059 40282
rect 8111 40230 11230 40282
rect 11282 40230 11294 40282
rect 11346 40230 11358 40282
rect 11410 40230 11422 40282
rect 11474 40230 11486 40282
rect 11538 40230 14657 40282
rect 14709 40230 14721 40282
rect 14773 40230 14785 40282
rect 14837 40230 14849 40282
rect 14901 40230 14913 40282
rect 14965 40230 14971 40282
rect 1104 40208 14971 40230
rect 1394 39992 1400 40044
rect 1452 39992 1458 40044
rect 13354 39992 13360 40044
rect 13412 39992 13418 40044
rect 13909 40035 13967 40041
rect 13909 40001 13921 40035
rect 13955 40001 13967 40035
rect 13909 39995 13967 40001
rect 10962 39924 10968 39976
rect 11020 39964 11026 39976
rect 13924 39964 13952 39995
rect 11020 39936 13952 39964
rect 11020 39924 11026 39936
rect 1581 39831 1639 39837
rect 1581 39797 1593 39831
rect 1627 39828 1639 39831
rect 7374 39828 7380 39840
rect 1627 39800 7380 39828
rect 1627 39797 1639 39800
rect 1581 39791 1639 39797
rect 7374 39788 7380 39800
rect 7432 39788 7438 39840
rect 13633 39831 13691 39837
rect 13633 39797 13645 39831
rect 13679 39828 13691 39831
rect 13998 39828 14004 39840
rect 13679 39800 14004 39828
rect 13679 39797 13691 39800
rect 13633 39791 13691 39797
rect 13998 39788 14004 39800
rect 14056 39788 14062 39840
rect 14182 39788 14188 39840
rect 14240 39788 14246 39840
rect 1104 39738 14812 39760
rect 1104 39686 2663 39738
rect 2715 39686 2727 39738
rect 2779 39686 2791 39738
rect 2843 39686 2855 39738
rect 2907 39686 2919 39738
rect 2971 39686 6090 39738
rect 6142 39686 6154 39738
rect 6206 39686 6218 39738
rect 6270 39686 6282 39738
rect 6334 39686 6346 39738
rect 6398 39686 9517 39738
rect 9569 39686 9581 39738
rect 9633 39686 9645 39738
rect 9697 39686 9709 39738
rect 9761 39686 9773 39738
rect 9825 39686 12944 39738
rect 12996 39686 13008 39738
rect 13060 39686 13072 39738
rect 13124 39686 13136 39738
rect 13188 39686 13200 39738
rect 13252 39686 14812 39738
rect 1104 39664 14812 39686
rect 8941 39627 8999 39633
rect 8941 39593 8953 39627
rect 8987 39624 8999 39627
rect 9493 39627 9551 39633
rect 8987 39596 9444 39624
rect 8987 39593 8999 39596
rect 8941 39587 8999 39593
rect 7377 39559 7435 39565
rect 7377 39525 7389 39559
rect 7423 39525 7435 39559
rect 7377 39519 7435 39525
rect 8113 39559 8171 39565
rect 8113 39525 8125 39559
rect 8159 39556 8171 39559
rect 9217 39559 9275 39565
rect 8159 39528 9168 39556
rect 8159 39525 8171 39528
rect 8113 39519 8171 39525
rect 7392 39488 7420 39519
rect 7392 39460 8340 39488
rect 750 39380 756 39432
rect 808 39420 814 39432
rect 8312 39429 8340 39460
rect 1397 39423 1455 39429
rect 1397 39420 1409 39423
rect 808 39392 1409 39420
rect 808 39380 814 39392
rect 1397 39389 1409 39392
rect 1443 39389 1455 39423
rect 7561 39423 7619 39429
rect 7561 39420 7573 39423
rect 1397 39383 1455 39389
rect 7392 39392 7573 39420
rect 7392 39364 7420 39392
rect 7561 39389 7573 39392
rect 7607 39389 7619 39423
rect 7561 39383 7619 39389
rect 8297 39423 8355 39429
rect 8297 39389 8309 39423
rect 8343 39389 8355 39423
rect 8297 39383 8355 39389
rect 8386 39380 8392 39432
rect 8444 39420 8450 39432
rect 9140 39429 9168 39528
rect 9217 39525 9229 39559
rect 9263 39525 9275 39559
rect 9416 39556 9444 39596
rect 9493 39593 9505 39627
rect 9539 39624 9551 39627
rect 10962 39624 10968 39636
rect 9539 39596 10968 39624
rect 9539 39593 9551 39596
rect 9493 39587 9551 39593
rect 10962 39584 10968 39596
rect 11020 39584 11026 39636
rect 13354 39624 13360 39636
rect 12406 39596 13360 39624
rect 12406 39556 12434 39596
rect 13354 39584 13360 39596
rect 13412 39584 13418 39636
rect 9416 39528 12434 39556
rect 13081 39559 13139 39565
rect 9217 39519 9275 39525
rect 13081 39525 13093 39559
rect 13127 39525 13139 39559
rect 13081 39519 13139 39525
rect 9232 39488 9260 39519
rect 9232 39460 9720 39488
rect 9692 39429 9720 39460
rect 8573 39423 8631 39429
rect 8573 39420 8585 39423
rect 8444 39392 8585 39420
rect 8444 39380 8450 39392
rect 8573 39389 8585 39392
rect 8619 39389 8631 39423
rect 8573 39383 8631 39389
rect 9125 39423 9183 39429
rect 9125 39389 9137 39423
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9401 39423 9459 39429
rect 9401 39389 9413 39423
rect 9447 39389 9459 39423
rect 9401 39383 9459 39389
rect 9677 39423 9735 39429
rect 9677 39389 9689 39423
rect 9723 39389 9735 39423
rect 9677 39383 9735 39389
rect 7374 39312 7380 39364
rect 7432 39312 7438 39364
rect 9416 39352 9444 39383
rect 12710 39380 12716 39432
rect 12768 39380 12774 39432
rect 12989 39423 13047 39429
rect 12989 39389 13001 39423
rect 13035 39420 13047 39423
rect 13096 39420 13124 39519
rect 13035 39392 13124 39420
rect 13265 39423 13323 39429
rect 13035 39389 13047 39392
rect 12989 39383 13047 39389
rect 13265 39389 13277 39423
rect 13311 39420 13323 39423
rect 13354 39420 13360 39432
rect 13311 39392 13360 39420
rect 13311 39389 13323 39392
rect 13265 39383 13323 39389
rect 13354 39380 13360 39392
rect 13412 39380 13418 39432
rect 14185 39423 14243 39429
rect 14185 39389 14197 39423
rect 14231 39389 14243 39423
rect 14185 39383 14243 39389
rect 13541 39355 13599 39361
rect 13541 39352 13553 39355
rect 8404 39324 9444 39352
rect 12544 39324 13553 39352
rect 1581 39287 1639 39293
rect 1581 39253 1593 39287
rect 1627 39284 1639 39287
rect 7558 39284 7564 39296
rect 1627 39256 7564 39284
rect 1627 39253 1639 39256
rect 1581 39247 1639 39253
rect 7558 39244 7564 39256
rect 7616 39244 7622 39296
rect 8404 39293 8432 39324
rect 12544 39293 12572 39324
rect 13541 39321 13553 39324
rect 13587 39321 13599 39355
rect 13541 39315 13599 39321
rect 13906 39312 13912 39364
rect 13964 39312 13970 39364
rect 8389 39287 8447 39293
rect 8389 39253 8401 39287
rect 8435 39253 8447 39287
rect 8389 39247 8447 39253
rect 12529 39287 12587 39293
rect 12529 39253 12541 39287
rect 12575 39253 12587 39287
rect 12529 39247 12587 39253
rect 12805 39287 12863 39293
rect 12805 39253 12817 39287
rect 12851 39284 12863 39287
rect 14200 39284 14228 39383
rect 12851 39256 14228 39284
rect 12851 39253 12863 39256
rect 12805 39247 12863 39253
rect 14366 39244 14372 39296
rect 14424 39244 14430 39296
rect 1104 39194 14971 39216
rect 1104 39142 4376 39194
rect 4428 39142 4440 39194
rect 4492 39142 4504 39194
rect 4556 39142 4568 39194
rect 4620 39142 4632 39194
rect 4684 39142 7803 39194
rect 7855 39142 7867 39194
rect 7919 39142 7931 39194
rect 7983 39142 7995 39194
rect 8047 39142 8059 39194
rect 8111 39142 11230 39194
rect 11282 39142 11294 39194
rect 11346 39142 11358 39194
rect 11410 39142 11422 39194
rect 11474 39142 11486 39194
rect 11538 39142 14657 39194
rect 14709 39142 14721 39194
rect 14773 39142 14785 39194
rect 14837 39142 14849 39194
rect 14901 39142 14913 39194
rect 14965 39142 14971 39194
rect 1104 39120 14971 39142
rect 4985 39083 5043 39089
rect 4985 39049 4997 39083
rect 5031 39080 5043 39083
rect 5074 39080 5080 39092
rect 5031 39052 5080 39080
rect 5031 39049 5043 39052
rect 4985 39043 5043 39049
rect 5074 39040 5080 39052
rect 5132 39040 5138 39092
rect 11977 39083 12035 39089
rect 11977 39049 11989 39083
rect 12023 39080 12035 39083
rect 12710 39080 12716 39092
rect 12023 39052 12716 39080
rect 12023 39049 12035 39052
rect 11977 39043 12035 39049
rect 12710 39040 12716 39052
rect 12768 39040 12774 39092
rect 12805 39083 12863 39089
rect 12805 39049 12817 39083
rect 12851 39049 12863 39083
rect 12805 39043 12863 39049
rect 7558 38972 7564 39024
rect 7616 39012 7622 39024
rect 12820 39012 12848 39043
rect 13909 39015 13967 39021
rect 13909 39012 13921 39015
rect 7616 38984 12572 39012
rect 12820 38984 13921 39012
rect 7616 38972 7622 38984
rect 5166 38904 5172 38956
rect 5224 38904 5230 38956
rect 12161 38947 12219 38953
rect 12161 38913 12173 38947
rect 12207 38944 12219 38947
rect 12437 38947 12495 38953
rect 12207 38916 12296 38944
rect 12207 38913 12219 38916
rect 12161 38907 12219 38913
rect 12268 38817 12296 38916
rect 12437 38913 12449 38947
rect 12483 38944 12495 38947
rect 12544 38944 12572 38984
rect 13909 38981 13921 38984
rect 13955 38981 13967 39015
rect 13909 38975 13967 38981
rect 12483 38916 12572 38944
rect 12483 38913 12495 38916
rect 12437 38907 12495 38913
rect 12253 38811 12311 38817
rect 12253 38777 12265 38811
rect 12299 38777 12311 38811
rect 12544 38808 12572 38916
rect 12618 38904 12624 38956
rect 12676 38944 12682 38956
rect 12713 38947 12771 38953
rect 12713 38944 12725 38947
rect 12676 38916 12725 38944
rect 12676 38904 12682 38916
rect 12713 38913 12725 38916
rect 12759 38913 12771 38947
rect 12713 38907 12771 38913
rect 12802 38904 12808 38956
rect 12860 38944 12866 38956
rect 12989 38947 13047 38953
rect 12989 38944 13001 38947
rect 12860 38916 13001 38944
rect 12860 38904 12866 38916
rect 12989 38913 13001 38916
rect 13035 38913 13047 38947
rect 12989 38907 13047 38913
rect 13357 38947 13415 38953
rect 13357 38913 13369 38947
rect 13403 38944 13415 38947
rect 13446 38944 13452 38956
rect 13403 38916 13452 38944
rect 13403 38913 13415 38916
rect 13357 38907 13415 38913
rect 13446 38904 13452 38916
rect 13504 38904 13510 38956
rect 12544 38780 14504 38808
rect 12253 38771 12311 38777
rect 14476 38752 14504 38780
rect 12529 38743 12587 38749
rect 12529 38709 12541 38743
rect 12575 38740 12587 38743
rect 13262 38740 13268 38752
rect 12575 38712 13268 38740
rect 12575 38709 12587 38712
rect 12529 38703 12587 38709
rect 13262 38700 13268 38712
rect 13320 38700 13326 38752
rect 13630 38700 13636 38752
rect 13688 38700 13694 38752
rect 14182 38700 14188 38752
rect 14240 38700 14246 38752
rect 14458 38700 14464 38752
rect 14516 38700 14522 38752
rect 1104 38650 14812 38672
rect 1104 38598 2663 38650
rect 2715 38598 2727 38650
rect 2779 38598 2791 38650
rect 2843 38598 2855 38650
rect 2907 38598 2919 38650
rect 2971 38598 6090 38650
rect 6142 38598 6154 38650
rect 6206 38598 6218 38650
rect 6270 38598 6282 38650
rect 6334 38598 6346 38650
rect 6398 38598 9517 38650
rect 9569 38598 9581 38650
rect 9633 38598 9645 38650
rect 9697 38598 9709 38650
rect 9761 38598 9773 38650
rect 9825 38598 12944 38650
rect 12996 38598 13008 38650
rect 13060 38598 13072 38650
rect 13124 38598 13136 38650
rect 13188 38598 13200 38650
rect 13252 38598 14812 38650
rect 1104 38576 14812 38598
rect 4801 38539 4859 38545
rect 4801 38505 4813 38539
rect 4847 38536 4859 38539
rect 5166 38536 5172 38548
rect 4847 38508 5172 38536
rect 4847 38505 4859 38508
rect 4801 38499 4859 38505
rect 5166 38496 5172 38508
rect 5224 38496 5230 38548
rect 12529 38539 12587 38545
rect 12529 38505 12541 38539
rect 12575 38536 12587 38539
rect 13354 38536 13360 38548
rect 12575 38508 13360 38536
rect 12575 38505 12587 38508
rect 12529 38499 12587 38505
rect 13354 38496 13360 38508
rect 13412 38496 13418 38548
rect 12434 38428 12440 38480
rect 12492 38468 12498 38480
rect 12710 38468 12716 38480
rect 12492 38440 12716 38468
rect 12492 38428 12498 38440
rect 12710 38428 12716 38440
rect 12768 38428 12774 38480
rect 12989 38471 13047 38477
rect 12989 38437 13001 38471
rect 13035 38437 13047 38471
rect 12989 38431 13047 38437
rect 13004 38400 13032 38431
rect 13004 38372 14228 38400
rect 750 38292 756 38344
rect 808 38332 814 38344
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 808 38304 1409 38332
rect 808 38292 814 38304
rect 1397 38301 1409 38304
rect 1443 38301 1455 38335
rect 1397 38295 1455 38301
rect 2130 38292 2136 38344
rect 2188 38332 2194 38344
rect 4985 38335 5043 38341
rect 4985 38332 4997 38335
rect 2188 38304 4997 38332
rect 2188 38292 2194 38304
rect 4985 38301 4997 38304
rect 5031 38301 5043 38335
rect 4985 38295 5043 38301
rect 11606 38292 11612 38344
rect 11664 38332 11670 38344
rect 12437 38335 12495 38341
rect 12437 38332 12449 38335
rect 11664 38304 12449 38332
rect 11664 38292 11670 38304
rect 12437 38301 12449 38304
rect 12483 38301 12495 38335
rect 12437 38295 12495 38301
rect 12713 38335 12771 38341
rect 12713 38301 12725 38335
rect 12759 38301 12771 38335
rect 12713 38295 12771 38301
rect 9398 38264 9404 38276
rect 1596 38236 9404 38264
rect 1596 38205 1624 38236
rect 9398 38224 9404 38236
rect 9456 38264 9462 38276
rect 12728 38264 12756 38295
rect 13170 38292 13176 38344
rect 13228 38292 13234 38344
rect 13262 38292 13268 38344
rect 13320 38292 13326 38344
rect 13354 38292 13360 38344
rect 13412 38332 13418 38344
rect 14200 38341 14228 38372
rect 13541 38335 13599 38341
rect 13541 38332 13553 38335
rect 13412 38304 13553 38332
rect 13412 38292 13418 38304
rect 13541 38301 13553 38304
rect 13587 38301 13599 38335
rect 13541 38295 13599 38301
rect 13633 38335 13691 38341
rect 13633 38301 13645 38335
rect 13679 38301 13691 38335
rect 13633 38295 13691 38301
rect 14185 38335 14243 38341
rect 14185 38301 14197 38335
rect 14231 38301 14243 38335
rect 14185 38295 14243 38301
rect 9456 38236 12756 38264
rect 13280 38264 13308 38292
rect 13648 38264 13676 38295
rect 13280 38236 13676 38264
rect 9456 38224 9462 38236
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38165 1639 38199
rect 1581 38159 1639 38165
rect 12253 38199 12311 38205
rect 12253 38165 12265 38199
rect 12299 38196 12311 38199
rect 12618 38196 12624 38208
rect 12299 38168 12624 38196
rect 12299 38165 12311 38168
rect 12253 38159 12311 38165
rect 12618 38156 12624 38168
rect 12676 38156 12682 38208
rect 13262 38156 13268 38208
rect 13320 38196 13326 38208
rect 13357 38199 13415 38205
rect 13357 38196 13369 38199
rect 13320 38168 13369 38196
rect 13320 38156 13326 38168
rect 13357 38165 13369 38168
rect 13403 38165 13415 38199
rect 13357 38159 13415 38165
rect 13814 38156 13820 38208
rect 13872 38156 13878 38208
rect 14366 38156 14372 38208
rect 14424 38156 14430 38208
rect 1104 38106 14971 38128
rect 1104 38054 4376 38106
rect 4428 38054 4440 38106
rect 4492 38054 4504 38106
rect 4556 38054 4568 38106
rect 4620 38054 4632 38106
rect 4684 38054 7803 38106
rect 7855 38054 7867 38106
rect 7919 38054 7931 38106
rect 7983 38054 7995 38106
rect 8047 38054 8059 38106
rect 8111 38054 11230 38106
rect 11282 38054 11294 38106
rect 11346 38054 11358 38106
rect 11410 38054 11422 38106
rect 11474 38054 11486 38106
rect 11538 38054 14657 38106
rect 14709 38054 14721 38106
rect 14773 38054 14785 38106
rect 14837 38054 14849 38106
rect 14901 38054 14913 38106
rect 14965 38054 14971 38106
rect 1104 38032 14971 38054
rect 11517 37995 11575 38001
rect 11517 37961 11529 37995
rect 11563 37992 11575 37995
rect 11790 37992 11796 38004
rect 11563 37964 11796 37992
rect 11563 37961 11575 37964
rect 11517 37955 11575 37961
rect 11790 37952 11796 37964
rect 11848 37952 11854 38004
rect 11885 37995 11943 38001
rect 11885 37961 11897 37995
rect 11931 37961 11943 37995
rect 11885 37955 11943 37961
rect 12345 37995 12403 38001
rect 12345 37961 12357 37995
rect 12391 37992 12403 37995
rect 12526 37992 12532 38004
rect 12391 37964 12532 37992
rect 12391 37961 12403 37964
rect 12345 37955 12403 37961
rect 11900 37924 11928 37955
rect 12526 37952 12532 37964
rect 12584 37952 12590 38004
rect 12621 37995 12679 38001
rect 12621 37961 12633 37995
rect 12667 37992 12679 37995
rect 12897 37995 12955 38001
rect 12667 37964 12848 37992
rect 12667 37961 12679 37964
rect 12621 37955 12679 37961
rect 12434 37924 12440 37936
rect 11900 37896 12440 37924
rect 12434 37884 12440 37896
rect 12492 37884 12498 37936
rect 12820 37924 12848 37964
rect 12897 37961 12909 37995
rect 12943 37992 12955 37995
rect 13170 37992 13176 38004
rect 12943 37964 13176 37992
rect 12943 37961 12955 37964
rect 12897 37955 12955 37961
rect 13170 37952 13176 37964
rect 13228 37952 13234 38004
rect 13357 37927 13415 37933
rect 13357 37924 13369 37927
rect 12820 37896 13369 37924
rect 13357 37893 13369 37896
rect 13403 37893 13415 37927
rect 13357 37887 13415 37893
rect 750 37816 756 37868
rect 808 37856 814 37868
rect 1397 37859 1455 37865
rect 1397 37856 1409 37859
rect 808 37828 1409 37856
rect 808 37816 814 37828
rect 1397 37825 1409 37828
rect 1443 37825 1455 37859
rect 1397 37819 1455 37825
rect 10778 37816 10784 37868
rect 10836 37856 10842 37868
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 10836 37828 11713 37856
rect 10836 37816 10842 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 12066 37816 12072 37868
rect 12124 37816 12130 37868
rect 12526 37816 12532 37868
rect 12584 37816 12590 37868
rect 12805 37859 12863 37865
rect 12805 37825 12817 37859
rect 12851 37825 12863 37859
rect 12805 37819 12863 37825
rect 12820 37788 12848 37819
rect 13078 37816 13084 37868
rect 13136 37816 13142 37868
rect 13262 37816 13268 37868
rect 13320 37816 13326 37868
rect 13909 37859 13967 37865
rect 13909 37825 13921 37859
rect 13955 37825 13967 37859
rect 13909 37819 13967 37825
rect 13280 37788 13308 37816
rect 12820 37760 13308 37788
rect 12342 37680 12348 37732
rect 12400 37720 12406 37732
rect 13924 37720 13952 37819
rect 12400 37692 13952 37720
rect 12400 37680 12406 37692
rect 1581 37655 1639 37661
rect 1581 37621 1593 37655
rect 1627 37652 1639 37655
rect 5718 37652 5724 37664
rect 1627 37624 5724 37652
rect 1627 37621 1639 37624
rect 1581 37615 1639 37621
rect 5718 37612 5724 37624
rect 5776 37652 5782 37664
rect 6546 37652 6552 37664
rect 5776 37624 6552 37652
rect 5776 37612 5782 37624
rect 6546 37612 6552 37624
rect 6604 37612 6610 37664
rect 12618 37612 12624 37664
rect 12676 37652 12682 37664
rect 13538 37652 13544 37664
rect 12676 37624 13544 37652
rect 12676 37612 12682 37624
rect 13538 37612 13544 37624
rect 13596 37612 13602 37664
rect 13630 37612 13636 37664
rect 13688 37612 13694 37664
rect 14182 37612 14188 37664
rect 14240 37612 14246 37664
rect 1104 37562 14812 37584
rect 1104 37510 2663 37562
rect 2715 37510 2727 37562
rect 2779 37510 2791 37562
rect 2843 37510 2855 37562
rect 2907 37510 2919 37562
rect 2971 37510 6090 37562
rect 6142 37510 6154 37562
rect 6206 37510 6218 37562
rect 6270 37510 6282 37562
rect 6334 37510 6346 37562
rect 6398 37510 9517 37562
rect 9569 37510 9581 37562
rect 9633 37510 9645 37562
rect 9697 37510 9709 37562
rect 9761 37510 9773 37562
rect 9825 37510 12944 37562
rect 12996 37510 13008 37562
rect 13060 37510 13072 37562
rect 13124 37510 13136 37562
rect 13188 37510 13200 37562
rect 13252 37510 14812 37562
rect 1104 37488 14812 37510
rect 10778 37408 10784 37460
rect 10836 37408 10842 37460
rect 11149 37451 11207 37457
rect 11149 37417 11161 37451
rect 11195 37448 11207 37451
rect 12066 37448 12072 37460
rect 11195 37420 12072 37448
rect 11195 37417 11207 37420
rect 11149 37411 11207 37417
rect 12066 37408 12072 37420
rect 12124 37408 12130 37460
rect 12342 37408 12348 37460
rect 12400 37408 12406 37460
rect 12621 37451 12679 37457
rect 12621 37417 12633 37451
rect 12667 37417 12679 37451
rect 12621 37411 12679 37417
rect 12636 37324 12664 37411
rect 12618 37272 12624 37324
rect 12676 37272 12682 37324
rect 10962 37204 10968 37256
rect 11020 37204 11026 37256
rect 11333 37247 11391 37253
rect 11333 37213 11345 37247
rect 11379 37213 11391 37247
rect 11333 37207 11391 37213
rect 6546 37136 6552 37188
rect 6604 37176 6610 37188
rect 11348 37176 11376 37207
rect 11882 37204 11888 37256
rect 11940 37244 11946 37256
rect 12529 37247 12587 37253
rect 12529 37244 12541 37247
rect 11940 37216 12541 37244
rect 11940 37204 11946 37216
rect 12529 37213 12541 37216
rect 12575 37213 12587 37247
rect 12529 37207 12587 37213
rect 12802 37204 12808 37256
rect 12860 37204 12866 37256
rect 12894 37204 12900 37256
rect 12952 37244 12958 37256
rect 13081 37247 13139 37253
rect 13081 37244 13093 37247
rect 12952 37216 13093 37244
rect 12952 37204 12958 37216
rect 13081 37213 13093 37216
rect 13127 37213 13139 37247
rect 13081 37207 13139 37213
rect 13262 37204 13268 37256
rect 13320 37244 13326 37256
rect 13357 37247 13415 37253
rect 13357 37244 13369 37247
rect 13320 37216 13369 37244
rect 13320 37204 13326 37216
rect 13357 37213 13369 37216
rect 13403 37213 13415 37247
rect 14185 37247 14243 37253
rect 14185 37244 14197 37247
rect 13357 37207 13415 37213
rect 13464 37216 14197 37244
rect 6604 37148 11376 37176
rect 6604 37136 6610 37148
rect 12158 37136 12164 37188
rect 12216 37176 12222 37188
rect 13464 37176 13492 37216
rect 14185 37213 14197 37216
rect 14231 37213 14243 37247
rect 14185 37207 14243 37213
rect 12216 37148 13492 37176
rect 12216 37136 12222 37148
rect 13538 37136 13544 37188
rect 13596 37136 13602 37188
rect 12710 37068 12716 37120
rect 12768 37108 12774 37120
rect 12897 37111 12955 37117
rect 12897 37108 12909 37111
rect 12768 37080 12909 37108
rect 12768 37068 12774 37080
rect 12897 37077 12909 37080
rect 12943 37077 12955 37111
rect 12897 37071 12955 37077
rect 13170 37068 13176 37120
rect 13228 37068 13234 37120
rect 13630 37068 13636 37120
rect 13688 37068 13694 37120
rect 14366 37068 14372 37120
rect 14424 37068 14430 37120
rect 1104 37018 14971 37040
rect 1104 36966 4376 37018
rect 4428 36966 4440 37018
rect 4492 36966 4504 37018
rect 4556 36966 4568 37018
rect 4620 36966 4632 37018
rect 4684 36966 7803 37018
rect 7855 36966 7867 37018
rect 7919 36966 7931 37018
rect 7983 36966 7995 37018
rect 8047 36966 8059 37018
rect 8111 36966 11230 37018
rect 11282 36966 11294 37018
rect 11346 36966 11358 37018
rect 11410 36966 11422 37018
rect 11474 36966 11486 37018
rect 11538 36966 14657 37018
rect 14709 36966 14721 37018
rect 14773 36966 14785 37018
rect 14837 36966 14849 37018
rect 14901 36966 14913 37018
rect 14965 36966 14971 37018
rect 1104 36944 14971 36966
rect 2133 36907 2191 36913
rect 2133 36873 2145 36907
rect 2179 36904 2191 36907
rect 2222 36904 2228 36916
rect 2179 36876 2228 36904
rect 2179 36873 2191 36876
rect 2133 36867 2191 36873
rect 2222 36864 2228 36876
rect 2280 36864 2286 36916
rect 9953 36907 10011 36913
rect 9953 36873 9965 36907
rect 9999 36904 10011 36907
rect 10962 36904 10968 36916
rect 9999 36876 10968 36904
rect 9999 36873 10011 36876
rect 9953 36867 10011 36873
rect 10962 36864 10968 36876
rect 11020 36864 11026 36916
rect 11606 36864 11612 36916
rect 11664 36864 11670 36916
rect 11882 36864 11888 36916
rect 11940 36864 11946 36916
rect 12161 36907 12219 36913
rect 12161 36873 12173 36907
rect 12207 36904 12219 36907
rect 12342 36904 12348 36916
rect 12207 36876 12348 36904
rect 12207 36873 12219 36876
rect 12161 36867 12219 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 13170 36904 13176 36916
rect 12544 36876 13176 36904
rect 12544 36836 12572 36876
rect 13170 36864 13176 36876
rect 13228 36864 13234 36916
rect 12084 36808 12572 36836
rect 750 36728 756 36780
rect 808 36768 814 36780
rect 1397 36771 1455 36777
rect 1397 36768 1409 36771
rect 808 36740 1409 36768
rect 808 36728 814 36740
rect 1397 36737 1409 36740
rect 1443 36737 1455 36771
rect 1397 36731 1455 36737
rect 2317 36771 2375 36777
rect 2317 36737 2329 36771
rect 2363 36768 2375 36771
rect 4246 36768 4252 36780
rect 2363 36740 4252 36768
rect 2363 36737 2375 36740
rect 2317 36731 2375 36737
rect 4246 36728 4252 36740
rect 4304 36728 4310 36780
rect 12084 36777 12112 36808
rect 10137 36771 10195 36777
rect 10137 36737 10149 36771
rect 10183 36737 10195 36771
rect 10137 36731 10195 36737
rect 11793 36771 11851 36777
rect 11793 36737 11805 36771
rect 11839 36737 11851 36771
rect 11793 36731 11851 36737
rect 12069 36771 12127 36777
rect 12069 36737 12081 36771
rect 12115 36737 12127 36771
rect 12321 36771 12379 36777
rect 12321 36768 12333 36771
rect 12069 36731 12127 36737
rect 12176 36740 12333 36768
rect 5166 36700 5172 36712
rect 2746 36672 5172 36700
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 2746 36564 2774 36672
rect 5166 36660 5172 36672
rect 5224 36700 5230 36712
rect 10152 36700 10180 36731
rect 5224 36672 10180 36700
rect 5224 36660 5230 36672
rect 8294 36592 8300 36644
rect 8352 36632 8358 36644
rect 11330 36632 11336 36644
rect 8352 36604 11336 36632
rect 8352 36592 8358 36604
rect 11330 36592 11336 36604
rect 11388 36592 11394 36644
rect 1627 36536 2774 36564
rect 11808 36564 11836 36731
rect 11882 36660 11888 36712
rect 11940 36700 11946 36712
rect 12176 36700 12204 36740
rect 12321 36737 12333 36740
rect 12367 36737 12379 36771
rect 12321 36731 12379 36737
rect 12710 36728 12716 36780
rect 12768 36728 12774 36780
rect 12986 36728 12992 36780
rect 13044 36728 13050 36780
rect 13357 36771 13415 36777
rect 13357 36737 13369 36771
rect 13403 36768 13415 36771
rect 13446 36768 13452 36780
rect 13403 36740 13452 36768
rect 13403 36737 13415 36740
rect 13357 36731 13415 36737
rect 13446 36728 13452 36740
rect 13504 36728 13510 36780
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 14093 36771 14151 36777
rect 14093 36737 14105 36771
rect 14139 36737 14151 36771
rect 14093 36731 14151 36737
rect 11940 36672 12204 36700
rect 11940 36660 11946 36672
rect 13173 36635 13231 36641
rect 13173 36632 13185 36635
rect 12452 36604 13185 36632
rect 12452 36564 12480 36604
rect 13173 36601 13185 36604
rect 13219 36601 13231 36635
rect 13173 36595 13231 36601
rect 13354 36592 13360 36644
rect 13412 36592 13418 36644
rect 13446 36592 13452 36644
rect 13504 36632 13510 36644
rect 13556 36632 13584 36731
rect 13630 36660 13636 36712
rect 13688 36700 13694 36712
rect 14108 36700 14136 36731
rect 13688 36672 14136 36700
rect 13688 36660 13694 36672
rect 13504 36604 13584 36632
rect 13504 36592 13510 36604
rect 11808 36536 12480 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 12526 36524 12532 36576
rect 12584 36524 12590 36576
rect 12805 36567 12863 36573
rect 12805 36533 12817 36567
rect 12851 36564 12863 36567
rect 13372 36564 13400 36592
rect 12851 36536 13400 36564
rect 12851 36533 12863 36536
rect 12805 36527 12863 36533
rect 13814 36524 13820 36576
rect 13872 36524 13878 36576
rect 14369 36567 14427 36573
rect 14369 36533 14381 36567
rect 14415 36564 14427 36567
rect 15286 36564 15292 36576
rect 14415 36536 15292 36564
rect 14415 36533 14427 36536
rect 14369 36527 14427 36533
rect 15286 36524 15292 36536
rect 15344 36524 15350 36576
rect 1104 36474 14812 36496
rect 1104 36422 2663 36474
rect 2715 36422 2727 36474
rect 2779 36422 2791 36474
rect 2843 36422 2855 36474
rect 2907 36422 2919 36474
rect 2971 36422 6090 36474
rect 6142 36422 6154 36474
rect 6206 36422 6218 36474
rect 6270 36422 6282 36474
rect 6334 36422 6346 36474
rect 6398 36422 9517 36474
rect 9569 36422 9581 36474
rect 9633 36422 9645 36474
rect 9697 36422 9709 36474
rect 9761 36422 9773 36474
rect 9825 36422 12944 36474
rect 12996 36422 13008 36474
rect 13060 36422 13072 36474
rect 13124 36422 13136 36474
rect 13188 36422 13200 36474
rect 13252 36422 14812 36474
rect 1104 36400 14812 36422
rect 1581 36363 1639 36369
rect 1581 36329 1593 36363
rect 1627 36360 1639 36363
rect 7282 36360 7288 36372
rect 1627 36332 7288 36360
rect 1627 36329 1639 36332
rect 1581 36323 1639 36329
rect 7282 36320 7288 36332
rect 7340 36320 7346 36372
rect 12158 36320 12164 36372
rect 12216 36320 12222 36372
rect 12526 36320 12532 36372
rect 12584 36320 12590 36372
rect 12710 36320 12716 36372
rect 12768 36360 12774 36372
rect 13446 36360 13452 36372
rect 12768 36332 13452 36360
rect 12768 36320 12774 36332
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 12544 36224 12572 36320
rect 12618 36252 12624 36304
rect 12676 36292 12682 36304
rect 12894 36292 12900 36304
rect 12676 36264 12900 36292
rect 12676 36252 12682 36264
rect 12894 36252 12900 36264
rect 12952 36252 12958 36304
rect 12544 36196 13124 36224
rect 1394 36116 1400 36168
rect 1452 36116 1458 36168
rect 12345 36159 12403 36165
rect 12345 36125 12357 36159
rect 12391 36156 12403 36159
rect 12434 36156 12440 36168
rect 12391 36128 12440 36156
rect 12391 36125 12403 36128
rect 12345 36119 12403 36125
rect 12434 36116 12440 36128
rect 12492 36116 12498 36168
rect 12618 36116 12624 36168
rect 12676 36116 12682 36168
rect 12710 36116 12716 36168
rect 12768 36116 12774 36168
rect 12802 36116 12808 36168
rect 12860 36116 12866 36168
rect 13096 36165 13124 36196
rect 13081 36159 13139 36165
rect 13081 36125 13093 36159
rect 13127 36125 13139 36159
rect 13081 36119 13139 36125
rect 13170 36116 13176 36168
rect 13228 36156 13234 36168
rect 13357 36159 13415 36165
rect 13357 36156 13369 36159
rect 13228 36128 13369 36156
rect 13228 36116 13234 36128
rect 13357 36125 13369 36128
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 13446 36116 13452 36168
rect 13504 36156 13510 36168
rect 14185 36159 14243 36165
rect 14185 36156 14197 36159
rect 13504 36128 14197 36156
rect 13504 36116 13510 36128
rect 14185 36125 14197 36128
rect 14231 36125 14243 36159
rect 14185 36119 14243 36125
rect 10962 36048 10968 36100
rect 11020 36088 11026 36100
rect 12728 36088 12756 36116
rect 11020 36060 12756 36088
rect 11020 36048 11026 36060
rect 12437 36023 12495 36029
rect 12437 35989 12449 36023
rect 12483 36020 12495 36023
rect 12820 36020 12848 36116
rect 13541 36091 13599 36097
rect 13541 36088 13553 36091
rect 12912 36060 13553 36088
rect 12912 36029 12940 36060
rect 13541 36057 13553 36060
rect 13587 36057 13599 36091
rect 13541 36051 13599 36057
rect 12483 35992 12848 36020
rect 12897 36023 12955 36029
rect 12483 35989 12495 35992
rect 12437 35983 12495 35989
rect 12897 35989 12909 36023
rect 12943 35989 12955 36023
rect 12897 35983 12955 35989
rect 13173 36023 13231 36029
rect 13173 35989 13185 36023
rect 13219 36020 13231 36023
rect 13354 36020 13360 36032
rect 13219 35992 13360 36020
rect 13219 35989 13231 35992
rect 13173 35983 13231 35989
rect 13354 35980 13360 35992
rect 13412 35980 13418 36032
rect 13722 35980 13728 36032
rect 13780 36020 13786 36032
rect 13817 36023 13875 36029
rect 13817 36020 13829 36023
rect 13780 35992 13829 36020
rect 13780 35980 13786 35992
rect 13817 35989 13829 35992
rect 13863 35989 13875 36023
rect 13817 35983 13875 35989
rect 14369 36023 14427 36029
rect 14369 35989 14381 36023
rect 14415 36020 14427 36023
rect 15102 36020 15108 36032
rect 14415 35992 15108 36020
rect 14415 35989 14427 35992
rect 14369 35983 14427 35989
rect 15102 35980 15108 35992
rect 15160 35980 15166 36032
rect 1104 35930 14971 35952
rect 1104 35878 4376 35930
rect 4428 35878 4440 35930
rect 4492 35878 4504 35930
rect 4556 35878 4568 35930
rect 4620 35878 4632 35930
rect 4684 35878 7803 35930
rect 7855 35878 7867 35930
rect 7919 35878 7931 35930
rect 7983 35878 7995 35930
rect 8047 35878 8059 35930
rect 8111 35878 11230 35930
rect 11282 35878 11294 35930
rect 11346 35878 11358 35930
rect 11410 35878 11422 35930
rect 11474 35878 11486 35930
rect 11538 35878 14657 35930
rect 14709 35878 14721 35930
rect 14773 35878 14785 35930
rect 14837 35878 14849 35930
rect 14901 35878 14913 35930
rect 14965 35878 14971 35930
rect 1104 35856 14971 35878
rect 10229 35819 10287 35825
rect 10229 35785 10241 35819
rect 10275 35816 10287 35819
rect 10275 35788 12434 35816
rect 10275 35785 10287 35788
rect 10229 35779 10287 35785
rect 11974 35748 11980 35760
rect 11808 35720 11980 35748
rect 10410 35640 10416 35692
rect 10468 35640 10474 35692
rect 10686 35640 10692 35692
rect 10744 35640 10750 35692
rect 11808 35689 11836 35720
rect 11974 35708 11980 35720
rect 12032 35708 12038 35760
rect 12406 35748 12434 35788
rect 13446 35748 13452 35760
rect 12406 35720 13452 35748
rect 13446 35708 13452 35720
rect 13504 35708 13510 35760
rect 11791 35683 11849 35689
rect 11791 35649 11803 35683
rect 11837 35649 11849 35683
rect 11791 35643 11849 35649
rect 11882 35640 11888 35692
rect 11940 35680 11946 35692
rect 12989 35683 13047 35689
rect 12989 35680 13001 35683
rect 11940 35652 13001 35680
rect 11940 35640 11946 35652
rect 12989 35649 13001 35652
rect 13035 35649 13047 35683
rect 12989 35643 13047 35649
rect 13541 35683 13599 35689
rect 13541 35649 13553 35683
rect 13587 35649 13599 35683
rect 13541 35643 13599 35649
rect 11514 35572 11520 35624
rect 11572 35572 11578 35624
rect 12434 35572 12440 35624
rect 12492 35612 12498 35624
rect 13170 35612 13176 35624
rect 12492 35584 13176 35612
rect 12492 35572 12498 35584
rect 13170 35572 13176 35584
rect 13228 35572 13234 35624
rect 10962 35504 10968 35556
rect 11020 35504 11026 35556
rect 13556 35544 13584 35643
rect 13998 35640 14004 35692
rect 14056 35680 14062 35692
rect 14093 35683 14151 35689
rect 14093 35680 14105 35683
rect 14056 35652 14105 35680
rect 14056 35640 14062 35652
rect 14093 35649 14105 35652
rect 14139 35649 14151 35683
rect 14093 35643 14151 35649
rect 15102 35544 15108 35556
rect 12406 35516 13584 35544
rect 13740 35516 15108 35544
rect 10505 35479 10563 35485
rect 10505 35445 10517 35479
rect 10551 35476 10563 35479
rect 10980 35476 11008 35504
rect 10551 35448 11008 35476
rect 10551 35445 10563 35448
rect 10505 35439 10563 35445
rect 11146 35436 11152 35488
rect 11204 35476 11210 35488
rect 12406 35476 12434 35516
rect 11204 35448 12434 35476
rect 11204 35436 11210 35448
rect 12526 35436 12532 35488
rect 12584 35436 12590 35488
rect 13265 35479 13323 35485
rect 13265 35445 13277 35479
rect 13311 35476 13323 35479
rect 13740 35476 13768 35516
rect 15102 35504 15108 35516
rect 15160 35504 15166 35556
rect 13311 35448 13768 35476
rect 13311 35445 13323 35448
rect 13265 35439 13323 35445
rect 13814 35436 13820 35488
rect 13872 35436 13878 35488
rect 14366 35436 14372 35488
rect 14424 35436 14430 35488
rect 1104 35386 14812 35408
rect 1104 35334 2663 35386
rect 2715 35334 2727 35386
rect 2779 35334 2791 35386
rect 2843 35334 2855 35386
rect 2907 35334 2919 35386
rect 2971 35334 6090 35386
rect 6142 35334 6154 35386
rect 6206 35334 6218 35386
rect 6270 35334 6282 35386
rect 6334 35334 6346 35386
rect 6398 35334 9517 35386
rect 9569 35334 9581 35386
rect 9633 35334 9645 35386
rect 9697 35334 9709 35386
rect 9761 35334 9773 35386
rect 9825 35334 12944 35386
rect 12996 35334 13008 35386
rect 13060 35334 13072 35386
rect 13124 35334 13136 35386
rect 13188 35334 13200 35386
rect 13252 35334 14812 35386
rect 1104 35312 14812 35334
rect 1762 35232 1768 35284
rect 1820 35232 1826 35284
rect 9493 35275 9551 35281
rect 9493 35241 9505 35275
rect 9539 35272 9551 35275
rect 10410 35272 10416 35284
rect 9539 35244 10416 35272
rect 9539 35241 9551 35244
rect 9493 35235 9551 35241
rect 10410 35232 10416 35244
rect 10468 35232 10474 35284
rect 10686 35232 10692 35284
rect 10744 35232 10750 35284
rect 11977 35275 12035 35281
rect 11977 35241 11989 35275
rect 12023 35272 12035 35275
rect 13630 35272 13636 35284
rect 12023 35244 13636 35272
rect 12023 35241 12035 35244
rect 11977 35235 12035 35241
rect 13630 35232 13636 35244
rect 13688 35232 13694 35284
rect 1581 35207 1639 35213
rect 1581 35173 1593 35207
rect 1627 35204 1639 35207
rect 9769 35207 9827 35213
rect 1627 35176 2774 35204
rect 1627 35173 1639 35176
rect 1581 35167 1639 35173
rect 2746 35136 2774 35176
rect 9769 35173 9781 35207
rect 9815 35204 9827 35207
rect 10704 35204 10732 35232
rect 9815 35176 10732 35204
rect 12253 35207 12311 35213
rect 9815 35173 9827 35176
rect 9769 35167 9827 35173
rect 12253 35173 12265 35207
rect 12299 35173 12311 35207
rect 12253 35167 12311 35173
rect 12621 35207 12679 35213
rect 12621 35173 12633 35207
rect 12667 35204 12679 35207
rect 12667 35176 13400 35204
rect 12667 35173 12679 35176
rect 12621 35167 12679 35173
rect 5902 35136 5908 35148
rect 2746 35108 5908 35136
rect 5902 35096 5908 35108
rect 5960 35136 5966 35148
rect 11790 35136 11796 35148
rect 5960 35108 11796 35136
rect 5960 35096 5966 35108
rect 11790 35096 11796 35108
rect 11848 35096 11854 35148
rect 750 35028 756 35080
rect 808 35068 814 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 808 35040 1409 35068
rect 808 35028 814 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1946 35028 1952 35080
rect 2004 35028 2010 35080
rect 9674 35028 9680 35080
rect 9732 35028 9738 35080
rect 9953 35071 10011 35077
rect 9953 35037 9965 35071
rect 9999 35037 10011 35071
rect 9953 35031 10011 35037
rect 9030 34960 9036 35012
rect 9088 35000 9094 35012
rect 9968 35000 9996 35031
rect 11054 35028 11060 35080
rect 11112 35068 11118 35080
rect 11885 35071 11943 35077
rect 11885 35068 11897 35071
rect 11112 35040 11897 35068
rect 11112 35028 11118 35040
rect 11885 35037 11897 35040
rect 11931 35037 11943 35071
rect 11885 35031 11943 35037
rect 12161 35071 12219 35077
rect 12161 35037 12173 35071
rect 12207 35068 12219 35071
rect 12268 35068 12296 35167
rect 12342 35096 12348 35148
rect 12400 35136 12406 35148
rect 12400 35108 13124 35136
rect 12400 35096 12406 35108
rect 12207 35040 12296 35068
rect 12437 35071 12495 35077
rect 12207 35037 12219 35040
rect 12161 35031 12219 35037
rect 12437 35037 12449 35071
rect 12483 35037 12495 35071
rect 12437 35031 12495 35037
rect 9088 34972 9996 35000
rect 9088 34960 9094 34972
rect 12066 34960 12072 35012
rect 12124 35000 12130 35012
rect 12452 35000 12480 35031
rect 12618 35028 12624 35080
rect 12676 35068 12682 35080
rect 13096 35077 13124 35108
rect 13372 35077 13400 35176
rect 12805 35071 12863 35077
rect 12805 35068 12817 35071
rect 12676 35040 12817 35068
rect 12676 35028 12682 35040
rect 12805 35037 12817 35040
rect 12851 35037 12863 35071
rect 12805 35031 12863 35037
rect 13081 35071 13139 35077
rect 13081 35037 13093 35071
rect 13127 35037 13139 35071
rect 13081 35031 13139 35037
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35037 13415 35071
rect 13357 35031 13415 35037
rect 13722 35028 13728 35080
rect 13780 35068 13786 35080
rect 14277 35071 14335 35077
rect 14277 35068 14289 35071
rect 13780 35040 14289 35068
rect 13780 35028 13786 35040
rect 14277 35037 14289 35040
rect 14323 35037 14335 35071
rect 14277 35031 14335 35037
rect 12124 34972 12480 35000
rect 12124 34960 12130 34972
rect 13538 34960 13544 35012
rect 13596 34960 13602 35012
rect 13906 34960 13912 35012
rect 13964 34960 13970 35012
rect 11698 34892 11704 34944
rect 11756 34892 11762 34944
rect 12894 34892 12900 34944
rect 12952 34892 12958 34944
rect 13170 34892 13176 34944
rect 13228 34892 13234 34944
rect 14090 34892 14096 34944
rect 14148 34892 14154 34944
rect 1104 34842 14971 34864
rect 1104 34790 4376 34842
rect 4428 34790 4440 34842
rect 4492 34790 4504 34842
rect 4556 34790 4568 34842
rect 4620 34790 4632 34842
rect 4684 34790 7803 34842
rect 7855 34790 7867 34842
rect 7919 34790 7931 34842
rect 7983 34790 7995 34842
rect 8047 34790 8059 34842
rect 8111 34790 11230 34842
rect 11282 34790 11294 34842
rect 11346 34790 11358 34842
rect 11410 34790 11422 34842
rect 11474 34790 11486 34842
rect 11538 34790 14657 34842
rect 14709 34790 14721 34842
rect 14773 34790 14785 34842
rect 14837 34790 14849 34842
rect 14901 34790 14913 34842
rect 14965 34790 14971 34842
rect 1104 34768 14971 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 1765 34731 1823 34737
rect 1765 34697 1777 34731
rect 1811 34728 1823 34731
rect 1946 34728 1952 34740
rect 1811 34700 1952 34728
rect 1811 34697 1823 34700
rect 1765 34691 1823 34697
rect 1596 34660 1624 34691
rect 1946 34688 1952 34700
rect 2004 34688 2010 34740
rect 8757 34731 8815 34737
rect 8757 34697 8769 34731
rect 8803 34728 8815 34731
rect 9674 34728 9680 34740
rect 8803 34700 9680 34728
rect 8803 34697 8815 34700
rect 8757 34691 8815 34697
rect 9674 34688 9680 34700
rect 9732 34688 9738 34740
rect 9769 34731 9827 34737
rect 9769 34697 9781 34731
rect 9815 34697 9827 34731
rect 9769 34691 9827 34697
rect 10505 34731 10563 34737
rect 10505 34697 10517 34731
rect 10551 34728 10563 34731
rect 10551 34700 10916 34728
rect 10551 34697 10563 34700
rect 10505 34691 10563 34697
rect 4798 34660 4804 34672
rect 1596 34632 4804 34660
rect 4798 34620 4804 34632
rect 4856 34660 4862 34672
rect 5442 34660 5448 34672
rect 4856 34632 5448 34660
rect 4856 34620 4862 34632
rect 5442 34620 5448 34632
rect 5500 34620 5506 34672
rect 9030 34620 9036 34672
rect 9088 34620 9094 34672
rect 9784 34660 9812 34691
rect 10888 34660 10916 34700
rect 10962 34688 10968 34740
rect 11020 34688 11026 34740
rect 11146 34688 11152 34740
rect 11204 34688 11210 34740
rect 11609 34731 11667 34737
rect 11609 34697 11621 34731
rect 11655 34728 11667 34731
rect 12066 34728 12072 34740
rect 11655 34700 12072 34728
rect 11655 34697 11667 34700
rect 11609 34691 11667 34697
rect 12066 34688 12072 34700
rect 12124 34688 12130 34740
rect 12894 34688 12900 34740
rect 12952 34688 12958 34740
rect 12989 34731 13047 34737
rect 12989 34697 13001 34731
rect 13035 34697 13047 34731
rect 12989 34691 13047 34697
rect 11164 34660 11192 34688
rect 9784 34632 10732 34660
rect 10888 34632 11192 34660
rect 1394 34552 1400 34604
rect 1452 34552 1458 34604
rect 1946 34552 1952 34604
rect 2004 34552 2010 34604
rect 5810 34552 5816 34604
rect 5868 34592 5874 34604
rect 8941 34595 8999 34601
rect 8941 34592 8953 34595
rect 5868 34564 8953 34592
rect 5868 34552 5874 34564
rect 8941 34561 8953 34564
rect 8987 34561 8999 34595
rect 8941 34555 8999 34561
rect 6454 34484 6460 34536
rect 6512 34524 6518 34536
rect 8294 34524 8300 34536
rect 6512 34496 8300 34524
rect 6512 34484 6518 34496
rect 8294 34484 8300 34496
rect 8352 34484 8358 34536
rect 9048 34465 9076 34620
rect 9214 34552 9220 34604
rect 9272 34552 9278 34604
rect 9306 34552 9312 34604
rect 9364 34592 9370 34604
rect 9493 34595 9551 34601
rect 9493 34592 9505 34595
rect 9364 34564 9505 34592
rect 9364 34552 9370 34564
rect 9493 34561 9505 34564
rect 9539 34561 9551 34595
rect 9493 34555 9551 34561
rect 9950 34552 9956 34604
rect 10008 34552 10014 34604
rect 10704 34601 10732 34632
rect 11882 34620 11888 34672
rect 11940 34620 11946 34672
rect 12912 34660 12940 34688
rect 12544 34632 12940 34660
rect 10689 34595 10747 34601
rect 10689 34561 10701 34595
rect 10735 34561 10747 34595
rect 10689 34555 10747 34561
rect 10778 34552 10784 34604
rect 10836 34592 10842 34604
rect 11149 34595 11207 34601
rect 11149 34592 11161 34595
rect 10836 34564 11161 34592
rect 10836 34552 10842 34564
rect 11149 34561 11161 34564
rect 11195 34561 11207 34595
rect 11149 34555 11207 34561
rect 11790 34552 11796 34604
rect 11848 34552 11854 34604
rect 11900 34524 11928 34620
rect 12250 34552 12256 34604
rect 12308 34552 12314 34604
rect 12544 34601 12572 34632
rect 12529 34595 12587 34601
rect 12529 34561 12541 34595
rect 12575 34561 12587 34595
rect 12529 34555 12587 34561
rect 12805 34595 12863 34601
rect 12805 34561 12817 34595
rect 12851 34592 12863 34595
rect 13004 34592 13032 34691
rect 13170 34688 13176 34740
rect 13228 34728 13234 34740
rect 13228 34700 13952 34728
rect 13228 34688 13234 34700
rect 13924 34669 13952 34700
rect 13909 34663 13967 34669
rect 13909 34629 13921 34663
rect 13955 34629 13967 34663
rect 13909 34623 13967 34629
rect 12851 34564 13032 34592
rect 13173 34595 13231 34601
rect 12851 34561 12863 34564
rect 12805 34555 12863 34561
rect 13173 34561 13185 34595
rect 13219 34561 13231 34595
rect 13173 34555 13231 34561
rect 13357 34595 13415 34601
rect 13357 34561 13369 34595
rect 13403 34592 13415 34595
rect 13446 34592 13452 34604
rect 13403 34564 13452 34592
rect 13403 34561 13415 34564
rect 13357 34555 13415 34561
rect 9324 34496 11928 34524
rect 12084 34496 12664 34524
rect 9324 34465 9352 34496
rect 9033 34459 9091 34465
rect 9033 34425 9045 34459
rect 9079 34425 9091 34459
rect 9033 34419 9091 34425
rect 9309 34459 9367 34465
rect 9309 34425 9321 34459
rect 9355 34425 9367 34459
rect 9309 34419 9367 34425
rect 10134 34416 10140 34468
rect 10192 34456 10198 34468
rect 11974 34456 11980 34468
rect 10192 34428 11980 34456
rect 10192 34416 10198 34428
rect 11974 34416 11980 34428
rect 12032 34416 12038 34468
rect 12084 34465 12112 34496
rect 12069 34459 12127 34465
rect 12069 34425 12081 34459
rect 12115 34425 12127 34459
rect 12069 34419 12127 34425
rect 12345 34459 12403 34465
rect 12345 34425 12357 34459
rect 12391 34456 12403 34459
rect 12434 34456 12440 34468
rect 12391 34428 12440 34456
rect 12391 34425 12403 34428
rect 12345 34419 12403 34425
rect 12434 34416 12440 34428
rect 12492 34416 12498 34468
rect 12636 34456 12664 34496
rect 12710 34484 12716 34536
rect 12768 34524 12774 34536
rect 13188 34524 13216 34555
rect 13446 34552 13452 34564
rect 13504 34552 13510 34604
rect 12768 34496 13216 34524
rect 12768 34484 12774 34496
rect 12802 34456 12808 34468
rect 12636 34428 12808 34456
rect 12802 34416 12808 34428
rect 12860 34416 12866 34468
rect 12621 34391 12679 34397
rect 12621 34357 12633 34391
rect 12667 34388 12679 34391
rect 13262 34388 13268 34400
rect 12667 34360 13268 34388
rect 12667 34357 12679 34360
rect 12621 34351 12679 34357
rect 13262 34348 13268 34360
rect 13320 34348 13326 34400
rect 13630 34348 13636 34400
rect 13688 34348 13694 34400
rect 14182 34348 14188 34400
rect 14240 34348 14246 34400
rect 1104 34298 14812 34320
rect 1104 34246 2663 34298
rect 2715 34246 2727 34298
rect 2779 34246 2791 34298
rect 2843 34246 2855 34298
rect 2907 34246 2919 34298
rect 2971 34246 6090 34298
rect 6142 34246 6154 34298
rect 6206 34246 6218 34298
rect 6270 34246 6282 34298
rect 6334 34246 6346 34298
rect 6398 34246 9517 34298
rect 9569 34246 9581 34298
rect 9633 34246 9645 34298
rect 9697 34246 9709 34298
rect 9761 34246 9773 34298
rect 9825 34246 12944 34298
rect 12996 34246 13008 34298
rect 13060 34246 13072 34298
rect 13124 34246 13136 34298
rect 13188 34246 13200 34298
rect 13252 34246 14812 34298
rect 1104 34224 14812 34246
rect 1581 34187 1639 34193
rect 1581 34153 1593 34187
rect 1627 34184 1639 34187
rect 1946 34184 1952 34196
rect 1627 34156 1952 34184
rect 1627 34153 1639 34156
rect 1581 34147 1639 34153
rect 1946 34144 1952 34156
rect 2004 34144 2010 34196
rect 9217 34187 9275 34193
rect 9217 34153 9229 34187
rect 9263 34184 9275 34187
rect 9306 34184 9312 34196
rect 9263 34156 9312 34184
rect 9263 34153 9275 34156
rect 9217 34147 9275 34153
rect 9306 34144 9312 34156
rect 9364 34144 9370 34196
rect 9950 34144 9956 34196
rect 10008 34144 10014 34196
rect 10505 34187 10563 34193
rect 10505 34153 10517 34187
rect 10551 34184 10563 34187
rect 10778 34184 10784 34196
rect 10551 34156 10784 34184
rect 10551 34153 10563 34156
rect 10505 34147 10563 34153
rect 10778 34144 10784 34156
rect 10836 34144 10842 34196
rect 11698 34144 11704 34196
rect 11756 34184 11762 34196
rect 11756 34156 14228 34184
rect 11756 34144 11762 34156
rect 8941 34119 8999 34125
rect 8941 34085 8953 34119
rect 8987 34116 8999 34119
rect 9968 34116 9996 34144
rect 8987 34088 9996 34116
rect 10229 34119 10287 34125
rect 8987 34085 8999 34088
rect 8941 34079 8999 34085
rect 10229 34085 10241 34119
rect 10275 34085 10287 34119
rect 10229 34079 10287 34085
rect 12621 34119 12679 34125
rect 12621 34085 12633 34119
rect 12667 34085 12679 34119
rect 12621 34079 12679 34085
rect 12989 34119 13047 34125
rect 12989 34085 13001 34119
rect 13035 34116 13047 34119
rect 13722 34116 13728 34128
rect 13035 34088 13728 34116
rect 13035 34085 13047 34088
rect 12989 34079 13047 34085
rect 10244 34048 10272 34079
rect 12636 34048 12664 34079
rect 13722 34076 13728 34088
rect 13780 34076 13786 34128
rect 13814 34048 13820 34060
rect 10244 34020 11008 34048
rect 12636 34020 13820 34048
rect 1765 33983 1823 33989
rect 1765 33949 1777 33983
rect 1811 33980 1823 33983
rect 7098 33980 7104 33992
rect 1811 33952 7104 33980
rect 1811 33949 1823 33952
rect 1765 33943 1823 33949
rect 7098 33940 7104 33952
rect 7156 33940 7162 33992
rect 9122 33940 9128 33992
rect 9180 33940 9186 33992
rect 9398 33940 9404 33992
rect 9456 33940 9462 33992
rect 9582 33940 9588 33992
rect 9640 33980 9646 33992
rect 10980 33989 11008 34020
rect 13814 34008 13820 34020
rect 13872 34008 13878 34060
rect 10413 33983 10471 33989
rect 10413 33980 10425 33983
rect 9640 33952 10425 33980
rect 9640 33940 9646 33952
rect 10413 33949 10425 33952
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10689 33983 10747 33989
rect 10689 33949 10701 33983
rect 10735 33949 10747 33983
rect 10689 33943 10747 33949
rect 10965 33983 11023 33989
rect 10965 33949 10977 33983
rect 11011 33949 11023 33983
rect 10965 33943 11023 33949
rect 9858 33872 9864 33924
rect 9916 33912 9922 33924
rect 10704 33912 10732 33943
rect 11606 33940 11612 33992
rect 11664 33940 11670 33992
rect 11883 33983 11941 33989
rect 11883 33949 11895 33983
rect 11929 33980 11941 33983
rect 12250 33980 12256 33992
rect 11929 33952 12256 33980
rect 11929 33949 11941 33952
rect 11883 33943 11941 33949
rect 12250 33940 12256 33952
rect 12308 33940 12314 33992
rect 12406 33952 12848 33980
rect 12406 33912 12434 33952
rect 12820 33912 12848 33952
rect 13170 33940 13176 33992
rect 13228 33940 13234 33992
rect 13354 33940 13360 33992
rect 13412 33980 13418 33992
rect 14200 33989 14228 34156
rect 13541 33983 13599 33989
rect 13541 33980 13553 33983
rect 13412 33952 13553 33980
rect 13412 33940 13418 33952
rect 13541 33949 13553 33952
rect 13587 33949 13599 33983
rect 13541 33943 13599 33949
rect 14185 33983 14243 33989
rect 14185 33949 14197 33983
rect 14231 33949 14243 33983
rect 14185 33943 14243 33949
rect 9916 33884 10732 33912
rect 10796 33884 12434 33912
rect 12544 33884 12756 33912
rect 12820 33884 13308 33912
rect 9916 33872 9922 33884
rect 10796 33853 10824 33884
rect 10781 33847 10839 33853
rect 10781 33813 10793 33847
rect 10827 33813 10839 33847
rect 10781 33807 10839 33813
rect 11698 33804 11704 33856
rect 11756 33844 11762 33856
rect 12544 33844 12572 33884
rect 12728 33856 12756 33884
rect 11756 33816 12572 33844
rect 11756 33804 11762 33816
rect 12710 33804 12716 33856
rect 12768 33804 12774 33856
rect 13280 33844 13308 33884
rect 13906 33872 13912 33924
rect 13964 33872 13970 33924
rect 13998 33872 14004 33924
rect 14056 33872 14062 33924
rect 14016 33844 14044 33872
rect 13280 33816 14044 33844
rect 14366 33804 14372 33856
rect 14424 33804 14430 33856
rect 1104 33754 14971 33776
rect 1104 33702 4376 33754
rect 4428 33702 4440 33754
rect 4492 33702 4504 33754
rect 4556 33702 4568 33754
rect 4620 33702 4632 33754
rect 4684 33702 7803 33754
rect 7855 33702 7867 33754
rect 7919 33702 7931 33754
rect 7983 33702 7995 33754
rect 8047 33702 8059 33754
rect 8111 33702 11230 33754
rect 11282 33702 11294 33754
rect 11346 33702 11358 33754
rect 11410 33702 11422 33754
rect 11474 33702 11486 33754
rect 11538 33702 14657 33754
rect 14709 33702 14721 33754
rect 14773 33702 14785 33754
rect 14837 33702 14849 33754
rect 14901 33702 14913 33754
rect 14965 33702 14971 33754
rect 1104 33680 14971 33702
rect 1581 33643 1639 33649
rect 1581 33609 1593 33643
rect 1627 33640 1639 33643
rect 3694 33640 3700 33652
rect 1627 33612 3700 33640
rect 1627 33609 1639 33612
rect 1581 33603 1639 33609
rect 3694 33600 3700 33612
rect 3752 33640 3758 33652
rect 6454 33640 6460 33652
rect 3752 33612 6460 33640
rect 3752 33600 3758 33612
rect 6454 33600 6460 33612
rect 6512 33600 6518 33652
rect 8113 33643 8171 33649
rect 8113 33609 8125 33643
rect 8159 33640 8171 33643
rect 9398 33640 9404 33652
rect 8159 33612 9404 33640
rect 8159 33609 8171 33612
rect 8113 33603 8171 33609
rect 9398 33600 9404 33612
rect 9456 33600 9462 33652
rect 9582 33600 9588 33652
rect 9640 33600 9646 33652
rect 9858 33600 9864 33652
rect 9916 33600 9922 33652
rect 10413 33643 10471 33649
rect 10413 33609 10425 33643
rect 10459 33609 10471 33643
rect 10413 33603 10471 33609
rect 10428 33572 10456 33603
rect 13262 33600 13268 33652
rect 13320 33600 13326 33652
rect 10428 33544 11192 33572
rect 750 33464 756 33516
rect 808 33504 814 33516
rect 1397 33507 1455 33513
rect 1397 33504 1409 33507
rect 808 33476 1409 33504
rect 808 33464 814 33476
rect 1397 33473 1409 33476
rect 1443 33473 1455 33507
rect 1397 33467 1455 33473
rect 8294 33464 8300 33516
rect 8352 33464 8358 33516
rect 9769 33507 9827 33513
rect 9769 33473 9781 33507
rect 9815 33473 9827 33507
rect 9769 33467 9827 33473
rect 10045 33507 10103 33513
rect 10045 33473 10057 33507
rect 10091 33473 10103 33507
rect 10045 33467 10103 33473
rect 6454 33396 6460 33448
rect 6512 33436 6518 33448
rect 9784 33436 9812 33467
rect 6512 33408 9812 33436
rect 6512 33396 6518 33408
rect 7006 33328 7012 33380
rect 7064 33368 7070 33380
rect 10060 33368 10088 33467
rect 10594 33464 10600 33516
rect 10652 33464 10658 33516
rect 11164 33513 11192 33544
rect 11149 33507 11207 33513
rect 11149 33473 11161 33507
rect 11195 33473 11207 33507
rect 11149 33467 11207 33473
rect 11791 33507 11849 33513
rect 11791 33473 11803 33507
rect 11837 33504 11849 33507
rect 11882 33504 11888 33516
rect 11837 33476 11888 33504
rect 11837 33473 11849 33476
rect 11791 33467 11849 33473
rect 11882 33464 11888 33476
rect 11940 33504 11946 33516
rect 12342 33504 12348 33516
rect 11940 33476 12348 33504
rect 11940 33464 11946 33476
rect 12342 33464 12348 33476
rect 12400 33464 12406 33516
rect 12710 33464 12716 33516
rect 12768 33504 12774 33516
rect 13173 33507 13231 33513
rect 13173 33504 13185 33507
rect 12768 33476 13185 33504
rect 12768 33464 12774 33476
rect 13173 33473 13185 33476
rect 13219 33473 13231 33507
rect 13280 33504 13308 33600
rect 13722 33532 13728 33584
rect 13780 33572 13786 33584
rect 13909 33575 13967 33581
rect 13909 33572 13921 33575
rect 13780 33544 13921 33572
rect 13780 33532 13786 33544
rect 13909 33541 13921 33544
rect 13955 33541 13967 33575
rect 13909 33535 13967 33541
rect 13357 33507 13415 33513
rect 13357 33504 13369 33507
rect 13280 33476 13369 33504
rect 13173 33467 13231 33473
rect 13357 33473 13369 33476
rect 13403 33473 13415 33507
rect 13357 33467 13415 33473
rect 11514 33396 11520 33448
rect 11572 33396 11578 33448
rect 13446 33436 13452 33448
rect 12406 33408 13452 33436
rect 7064 33340 10088 33368
rect 10965 33371 11023 33377
rect 7064 33328 7070 33340
rect 10965 33337 10977 33371
rect 11011 33337 11023 33371
rect 10965 33331 11023 33337
rect 10980 33300 11008 33331
rect 12406 33300 12434 33408
rect 13446 33396 13452 33408
rect 13504 33396 13510 33448
rect 14274 33368 14280 33380
rect 13004 33340 14280 33368
rect 10980 33272 12434 33300
rect 12529 33303 12587 33309
rect 12529 33269 12541 33303
rect 12575 33300 12587 33303
rect 12802 33300 12808 33312
rect 12575 33272 12808 33300
rect 12575 33269 12587 33272
rect 12529 33263 12587 33269
rect 12802 33260 12808 33272
rect 12860 33260 12866 33312
rect 13004 33309 13032 33340
rect 14274 33328 14280 33340
rect 14332 33328 14338 33380
rect 12989 33303 13047 33309
rect 12989 33269 13001 33303
rect 13035 33269 13047 33303
rect 12989 33263 13047 33269
rect 13630 33260 13636 33312
rect 13688 33260 13694 33312
rect 14182 33260 14188 33312
rect 14240 33260 14246 33312
rect 1104 33210 14812 33232
rect 1104 33158 2663 33210
rect 2715 33158 2727 33210
rect 2779 33158 2791 33210
rect 2843 33158 2855 33210
rect 2907 33158 2919 33210
rect 2971 33158 6090 33210
rect 6142 33158 6154 33210
rect 6206 33158 6218 33210
rect 6270 33158 6282 33210
rect 6334 33158 6346 33210
rect 6398 33158 9517 33210
rect 9569 33158 9581 33210
rect 9633 33158 9645 33210
rect 9697 33158 9709 33210
rect 9761 33158 9773 33210
rect 9825 33158 12944 33210
rect 12996 33158 13008 33210
rect 13060 33158 13072 33210
rect 13124 33158 13136 33210
rect 13188 33158 13200 33210
rect 13252 33158 14812 33210
rect 1104 33136 14812 33158
rect 10045 33099 10103 33105
rect 10045 33065 10057 33099
rect 10091 33096 10103 33099
rect 10594 33096 10600 33108
rect 10091 33068 10600 33096
rect 10091 33065 10103 33068
rect 10045 33059 10103 33065
rect 10594 33056 10600 33068
rect 10652 33056 10658 33108
rect 10873 33099 10931 33105
rect 10873 33065 10885 33099
rect 10919 33096 10931 33099
rect 11054 33096 11060 33108
rect 10919 33068 11060 33096
rect 10919 33065 10931 33068
rect 10873 33059 10931 33065
rect 11054 33056 11060 33068
rect 11112 33056 11118 33108
rect 11149 33099 11207 33105
rect 11149 33065 11161 33099
rect 11195 33096 11207 33099
rect 12253 33099 12311 33105
rect 11195 33068 11928 33096
rect 11195 33065 11207 33068
rect 11149 33059 11207 33065
rect 11422 32988 11428 33040
rect 11480 32988 11486 33040
rect 11701 33031 11759 33037
rect 11701 32997 11713 33031
rect 11747 32997 11759 33031
rect 11701 32991 11759 32997
rect 11716 32960 11744 32991
rect 11072 32932 11744 32960
rect 11900 32960 11928 33068
rect 12253 33065 12265 33099
rect 12299 33096 12311 33099
rect 13722 33096 13728 33108
rect 12299 33068 13728 33096
rect 12299 33065 12311 33068
rect 12253 33059 12311 33065
rect 13722 33056 13728 33068
rect 13780 33056 13786 33108
rect 11977 33031 12035 33037
rect 11977 32997 11989 33031
rect 12023 33028 12035 33031
rect 13173 33031 13231 33037
rect 12023 33000 12434 33028
rect 12023 32997 12035 33000
rect 11977 32991 12035 32997
rect 12406 32960 12434 33000
rect 13173 32997 13185 33031
rect 13219 33028 13231 33031
rect 15562 33028 15568 33040
rect 13219 33000 15568 33028
rect 13219 32997 13231 33000
rect 13173 32991 13231 32997
rect 15562 32988 15568 33000
rect 15620 32988 15626 33040
rect 11900 32932 12204 32960
rect 12406 32932 12480 32960
rect 750 32852 756 32904
rect 808 32892 814 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 808 32864 1409 32892
rect 808 32852 814 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 9950 32852 9956 32904
rect 10008 32892 10014 32904
rect 11072 32901 11100 32932
rect 10229 32895 10287 32901
rect 10229 32892 10241 32895
rect 10008 32864 10241 32892
rect 10008 32852 10014 32864
rect 10229 32861 10241 32864
rect 10275 32861 10287 32895
rect 10229 32855 10287 32861
rect 11057 32895 11115 32901
rect 11057 32861 11069 32895
rect 11103 32861 11115 32895
rect 11057 32855 11115 32861
rect 11333 32895 11391 32901
rect 11333 32861 11345 32895
rect 11379 32861 11391 32895
rect 11333 32855 11391 32861
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 1670 32756 1676 32768
rect 1627 32728 1676 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 1670 32716 1676 32728
rect 1728 32716 1734 32768
rect 10962 32716 10968 32768
rect 11020 32756 11026 32768
rect 11348 32756 11376 32855
rect 11422 32852 11428 32904
rect 11480 32892 11486 32904
rect 12176 32901 12204 32932
rect 12452 32901 12480 32932
rect 12636 32932 13032 32960
rect 11609 32895 11667 32901
rect 11609 32892 11621 32895
rect 11480 32864 11621 32892
rect 11480 32852 11486 32864
rect 11609 32861 11621 32864
rect 11655 32861 11667 32895
rect 11885 32895 11943 32901
rect 11885 32892 11897 32895
rect 11609 32855 11667 32861
rect 11808 32864 11897 32892
rect 11808 32768 11836 32864
rect 11885 32861 11897 32864
rect 11931 32861 11943 32895
rect 11885 32855 11943 32861
rect 12161 32895 12219 32901
rect 12161 32861 12173 32895
rect 12207 32861 12219 32895
rect 12161 32855 12219 32861
rect 12437 32895 12495 32901
rect 12437 32861 12449 32895
rect 12483 32861 12495 32895
rect 12437 32855 12495 32861
rect 12066 32784 12072 32836
rect 12124 32824 12130 32836
rect 12636 32824 12664 32932
rect 12713 32895 12771 32901
rect 12713 32861 12725 32895
rect 12759 32892 12771 32895
rect 12894 32892 12900 32904
rect 12759 32864 12900 32892
rect 12759 32861 12771 32864
rect 12713 32855 12771 32861
rect 12894 32852 12900 32864
rect 12952 32852 12958 32904
rect 13004 32901 13032 32932
rect 12989 32895 13047 32901
rect 12989 32861 13001 32895
rect 13035 32861 13047 32895
rect 12989 32855 13047 32861
rect 13354 32852 13360 32904
rect 13412 32852 13418 32904
rect 14090 32852 14096 32904
rect 14148 32852 14154 32904
rect 13541 32827 13599 32833
rect 13541 32824 13553 32827
rect 12124 32796 12664 32824
rect 12820 32796 13553 32824
rect 12124 32784 12130 32796
rect 11020 32728 11376 32756
rect 11020 32716 11026 32728
rect 11790 32716 11796 32768
rect 11848 32716 11854 32768
rect 12529 32759 12587 32765
rect 12529 32725 12541 32759
rect 12575 32756 12587 32759
rect 12618 32756 12624 32768
rect 12575 32728 12624 32756
rect 12575 32725 12587 32728
rect 12529 32719 12587 32725
rect 12618 32716 12624 32728
rect 12676 32716 12682 32768
rect 12820 32765 12848 32796
rect 13541 32793 13553 32796
rect 13587 32793 13599 32827
rect 13541 32787 13599 32793
rect 13909 32827 13967 32833
rect 13909 32793 13921 32827
rect 13955 32824 13967 32827
rect 15102 32824 15108 32836
rect 13955 32796 15108 32824
rect 13955 32793 13967 32796
rect 13909 32787 13967 32793
rect 15102 32784 15108 32796
rect 15160 32784 15166 32836
rect 12805 32759 12863 32765
rect 12805 32725 12817 32759
rect 12851 32725 12863 32759
rect 12805 32719 12863 32725
rect 14274 32716 14280 32768
rect 14332 32716 14338 32768
rect 1104 32666 14971 32688
rect 1104 32614 4376 32666
rect 4428 32614 4440 32666
rect 4492 32614 4504 32666
rect 4556 32614 4568 32666
rect 4620 32614 4632 32666
rect 4684 32614 7803 32666
rect 7855 32614 7867 32666
rect 7919 32614 7931 32666
rect 7983 32614 7995 32666
rect 8047 32614 8059 32666
rect 8111 32614 11230 32666
rect 11282 32614 11294 32666
rect 11346 32614 11358 32666
rect 11410 32614 11422 32666
rect 11474 32614 11486 32666
rect 11538 32614 14657 32666
rect 14709 32614 14721 32666
rect 14773 32614 14785 32666
rect 14837 32614 14849 32666
rect 14901 32614 14913 32666
rect 14965 32614 14971 32666
rect 1104 32592 14971 32614
rect 1670 32512 1676 32564
rect 1728 32552 1734 32564
rect 11054 32552 11060 32564
rect 1728 32524 11060 32552
rect 1728 32512 1734 32524
rect 11054 32512 11060 32524
rect 11112 32512 11118 32564
rect 11330 32512 11336 32564
rect 11388 32552 11394 32564
rect 13262 32552 13268 32564
rect 11388 32524 13268 32552
rect 11388 32512 11394 32524
rect 13262 32512 13268 32524
rect 13320 32512 13326 32564
rect 8386 32484 8392 32496
rect 8312 32456 8392 32484
rect 8312 32455 8340 32456
rect 8279 32449 8340 32455
rect 7098 32376 7104 32428
rect 7156 32416 7162 32428
rect 7650 32416 7656 32428
rect 7156 32388 7656 32416
rect 7156 32376 7162 32388
rect 7650 32376 7656 32388
rect 7708 32416 7714 32428
rect 8021 32419 8079 32425
rect 8021 32416 8033 32419
rect 7708 32388 8033 32416
rect 7708 32376 7714 32388
rect 8021 32385 8033 32388
rect 8067 32385 8079 32419
rect 8279 32415 8291 32449
rect 8325 32418 8340 32449
rect 8386 32444 8392 32456
rect 8444 32484 8450 32496
rect 9122 32484 9128 32496
rect 8444 32456 9128 32484
rect 8444 32444 8450 32456
rect 9122 32444 9128 32456
rect 9180 32444 9186 32496
rect 10042 32484 10048 32496
rect 9692 32456 10048 32484
rect 9692 32455 9720 32456
rect 9659 32449 9720 32455
rect 8325 32415 8337 32418
rect 8279 32409 8337 32415
rect 9659 32415 9671 32449
rect 9705 32418 9720 32449
rect 10042 32444 10048 32456
rect 10100 32484 10106 32496
rect 10962 32484 10968 32496
rect 10100 32456 10968 32484
rect 10100 32444 10106 32456
rect 10962 32444 10968 32456
rect 11020 32444 11026 32496
rect 12434 32484 12440 32496
rect 11348 32456 12440 32484
rect 11348 32425 11376 32456
rect 12434 32444 12440 32456
rect 12492 32444 12498 32496
rect 11333 32419 11391 32425
rect 9705 32415 9717 32418
rect 9659 32409 9717 32415
rect 8021 32379 8079 32385
rect 11333 32385 11345 32419
rect 11379 32385 11391 32419
rect 11790 32416 11796 32428
rect 11751 32388 11796 32416
rect 11333 32379 11391 32385
rect 8036 32212 8064 32379
rect 11790 32376 11796 32388
rect 11848 32376 11854 32428
rect 12158 32376 12164 32428
rect 12216 32416 12222 32428
rect 13173 32419 13231 32425
rect 13173 32416 13185 32419
rect 12216 32388 13185 32416
rect 12216 32376 12222 32388
rect 13173 32385 13185 32388
rect 13219 32385 13231 32419
rect 13173 32379 13231 32385
rect 13722 32376 13728 32428
rect 13780 32376 13786 32428
rect 14182 32376 14188 32428
rect 14240 32376 14246 32428
rect 9401 32351 9459 32357
rect 9401 32348 9413 32351
rect 8680 32320 9413 32348
rect 8680 32212 8708 32320
rect 9401 32317 9413 32320
rect 9447 32317 9459 32351
rect 9401 32311 9459 32317
rect 11517 32351 11575 32357
rect 11517 32317 11529 32351
rect 11563 32317 11575 32351
rect 11517 32311 11575 32317
rect 11532 32280 11560 32311
rect 12710 32308 12716 32360
rect 12768 32348 12774 32360
rect 13630 32348 13636 32360
rect 12768 32320 13636 32348
rect 12768 32308 12774 32320
rect 13630 32308 13636 32320
rect 13688 32308 13694 32360
rect 11532 32252 11652 32280
rect 11624 32224 11652 32252
rect 8036 32184 8708 32212
rect 9030 32172 9036 32224
rect 9088 32172 9094 32224
rect 10410 32172 10416 32224
rect 10468 32172 10474 32224
rect 11146 32172 11152 32224
rect 11204 32172 11210 32224
rect 11606 32172 11612 32224
rect 11664 32172 11670 32224
rect 12529 32215 12587 32221
rect 12529 32181 12541 32215
rect 12575 32212 12587 32215
rect 12710 32212 12716 32224
rect 12575 32184 12716 32212
rect 12575 32181 12587 32184
rect 12529 32175 12587 32181
rect 12710 32172 12716 32184
rect 12768 32172 12774 32224
rect 13449 32215 13507 32221
rect 13449 32181 13461 32215
rect 13495 32212 13507 32215
rect 13906 32212 13912 32224
rect 13495 32184 13912 32212
rect 13495 32181 13507 32184
rect 13449 32175 13507 32181
rect 13906 32172 13912 32184
rect 13964 32172 13970 32224
rect 13998 32172 14004 32224
rect 14056 32172 14062 32224
rect 14366 32172 14372 32224
rect 14424 32172 14430 32224
rect 1104 32122 14812 32144
rect 1104 32070 2663 32122
rect 2715 32070 2727 32122
rect 2779 32070 2791 32122
rect 2843 32070 2855 32122
rect 2907 32070 2919 32122
rect 2971 32070 6090 32122
rect 6142 32070 6154 32122
rect 6206 32070 6218 32122
rect 6270 32070 6282 32122
rect 6334 32070 6346 32122
rect 6398 32070 9517 32122
rect 9569 32070 9581 32122
rect 9633 32070 9645 32122
rect 9697 32070 9709 32122
rect 9761 32070 9773 32122
rect 9825 32070 12944 32122
rect 12996 32070 13008 32122
rect 13060 32070 13072 32122
rect 13124 32070 13136 32122
rect 13188 32070 13200 32122
rect 13252 32070 14812 32122
rect 1104 32048 14812 32070
rect 1581 32011 1639 32017
rect 1581 31977 1593 32011
rect 1627 32008 1639 32011
rect 1762 32008 1768 32020
rect 1627 31980 1768 32008
rect 1627 31977 1639 31980
rect 1581 31971 1639 31977
rect 1762 31968 1768 31980
rect 1820 32008 1826 32020
rect 10134 32008 10140 32020
rect 1820 31980 10140 32008
rect 1820 31968 1826 31980
rect 10134 31968 10140 31980
rect 10192 31968 10198 32020
rect 11146 31968 11152 32020
rect 11204 32008 11210 32020
rect 11204 31980 11836 32008
rect 11204 31968 11210 31980
rect 7929 31943 7987 31949
rect 7929 31909 7941 31943
rect 7975 31940 7987 31943
rect 8202 31940 8208 31952
rect 7975 31912 8208 31940
rect 7975 31909 7987 31912
rect 7929 31903 7987 31909
rect 8202 31900 8208 31912
rect 8260 31900 8266 31952
rect 11330 31900 11336 31952
rect 11388 31900 11394 31952
rect 11609 31943 11667 31949
rect 11609 31909 11621 31943
rect 11655 31940 11667 31943
rect 11698 31940 11704 31952
rect 11655 31912 11704 31940
rect 11655 31909 11667 31912
rect 11609 31903 11667 31909
rect 11698 31900 11704 31912
rect 11756 31900 11762 31952
rect 6914 31832 6920 31884
rect 6972 31832 6978 31884
rect 11808 31872 11836 31980
rect 12158 31968 12164 32020
rect 12216 31968 12222 32020
rect 12434 31968 12440 32020
rect 12492 32008 12498 32020
rect 12621 32011 12679 32017
rect 12621 32008 12633 32011
rect 12492 31980 12633 32008
rect 12492 31968 12498 31980
rect 12621 31977 12633 31980
rect 12667 31977 12679 32011
rect 14182 32008 14188 32020
rect 12621 31971 12679 31977
rect 12912 31980 14188 32008
rect 11885 31943 11943 31949
rect 11885 31909 11897 31943
rect 11931 31940 11943 31943
rect 12912 31940 12940 31980
rect 14182 31968 14188 31980
rect 14240 31968 14246 32020
rect 11931 31912 12940 31940
rect 11931 31909 11943 31912
rect 11885 31903 11943 31909
rect 12526 31872 12532 31884
rect 9646 31844 11652 31872
rect 11808 31844 12112 31872
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 7191 31807 7249 31813
rect 7191 31773 7203 31807
rect 7237 31804 7249 31807
rect 8110 31804 8116 31816
rect 7237 31776 8116 31804
rect 7237 31773 7249 31776
rect 7191 31767 7249 31773
rect 7484 31748 7512 31776
rect 8110 31764 8116 31776
rect 8168 31764 8174 31816
rect 9214 31764 9220 31816
rect 9272 31804 9278 31816
rect 9646 31804 9674 31844
rect 9272 31776 9674 31804
rect 9272 31764 9278 31776
rect 11514 31764 11520 31816
rect 11572 31764 11578 31816
rect 11624 31804 11652 31844
rect 12084 31813 12112 31844
rect 12360 31844 12532 31872
rect 12360 31813 12388 31844
rect 12526 31832 12532 31844
rect 12584 31832 12590 31884
rect 11793 31807 11851 31813
rect 11793 31804 11805 31807
rect 11624 31776 11805 31804
rect 11793 31773 11805 31776
rect 11839 31773 11851 31807
rect 11793 31767 11851 31773
rect 12069 31807 12127 31813
rect 12069 31773 12081 31807
rect 12115 31773 12127 31807
rect 12069 31767 12127 31773
rect 12345 31807 12403 31813
rect 12345 31773 12357 31807
rect 12391 31773 12403 31807
rect 12345 31767 12403 31773
rect 12618 31764 12624 31816
rect 12676 31804 12682 31816
rect 12805 31807 12863 31813
rect 12805 31804 12817 31807
rect 12676 31776 12817 31804
rect 12676 31764 12682 31776
rect 12805 31773 12817 31776
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 12986 31764 12992 31816
rect 13044 31764 13050 31816
rect 14369 31807 14427 31813
rect 14369 31773 14381 31807
rect 14415 31804 14427 31807
rect 15654 31804 15660 31816
rect 14415 31776 15660 31804
rect 14415 31773 14427 31776
rect 14369 31767 14427 31773
rect 15654 31764 15660 31776
rect 15712 31764 15718 31816
rect 7466 31696 7472 31748
rect 7524 31696 7530 31748
rect 13541 31739 13599 31745
rect 13541 31736 13553 31739
rect 13004 31708 13553 31736
rect 11514 31628 11520 31680
rect 11572 31668 11578 31680
rect 11698 31668 11704 31680
rect 11572 31640 11704 31668
rect 11572 31628 11578 31640
rect 11698 31628 11704 31640
rect 11756 31628 11762 31680
rect 11790 31628 11796 31680
rect 11848 31668 11854 31680
rect 12250 31668 12256 31680
rect 11848 31640 12256 31668
rect 11848 31628 11854 31640
rect 12250 31628 12256 31640
rect 12308 31628 12314 31680
rect 12434 31628 12440 31680
rect 12492 31668 12498 31680
rect 13004 31668 13032 31708
rect 13541 31705 13553 31708
rect 13587 31705 13599 31739
rect 13541 31699 13599 31705
rect 12492 31640 13032 31668
rect 13265 31671 13323 31677
rect 12492 31628 12498 31640
rect 13265 31637 13277 31671
rect 13311 31668 13323 31671
rect 13354 31668 13360 31680
rect 13311 31640 13360 31668
rect 13311 31637 13323 31640
rect 13265 31631 13323 31637
rect 13354 31628 13360 31640
rect 13412 31628 13418 31680
rect 13817 31671 13875 31677
rect 13817 31637 13829 31671
rect 13863 31668 13875 31671
rect 13906 31668 13912 31680
rect 13863 31640 13912 31668
rect 13863 31637 13875 31640
rect 13817 31631 13875 31637
rect 13906 31628 13912 31640
rect 13964 31628 13970 31680
rect 14182 31628 14188 31680
rect 14240 31628 14246 31680
rect 1104 31578 14971 31600
rect 1104 31526 4376 31578
rect 4428 31526 4440 31578
rect 4492 31526 4504 31578
rect 4556 31526 4568 31578
rect 4620 31526 4632 31578
rect 4684 31526 7803 31578
rect 7855 31526 7867 31578
rect 7919 31526 7931 31578
rect 7983 31526 7995 31578
rect 8047 31526 8059 31578
rect 8111 31526 11230 31578
rect 11282 31526 11294 31578
rect 11346 31526 11358 31578
rect 11410 31526 11422 31578
rect 11474 31526 11486 31578
rect 11538 31526 14657 31578
rect 14709 31526 14721 31578
rect 14773 31526 14785 31578
rect 14837 31526 14849 31578
rect 14901 31526 14913 31578
rect 14965 31526 14971 31578
rect 1104 31504 14971 31526
rect 10962 31424 10968 31476
rect 11020 31424 11026 31476
rect 11974 31424 11980 31476
rect 12032 31424 12038 31476
rect 9214 31396 9220 31408
rect 8956 31368 9220 31396
rect 8956 31367 8984 31368
rect 8923 31361 8984 31367
rect 750 31288 756 31340
rect 808 31328 814 31340
rect 1397 31331 1455 31337
rect 1397 31328 1409 31331
rect 808 31300 1409 31328
rect 808 31288 814 31300
rect 1397 31297 1409 31300
rect 1443 31297 1455 31331
rect 1397 31291 1455 31297
rect 5442 31288 5448 31340
rect 5500 31328 5506 31340
rect 7527 31331 7585 31337
rect 7527 31328 7539 31331
rect 5500 31300 7539 31328
rect 5500 31288 5506 31300
rect 7527 31297 7539 31300
rect 7573 31328 7585 31331
rect 8294 31328 8300 31340
rect 7573 31300 8300 31328
rect 7573 31297 7585 31300
rect 7527 31291 7585 31297
rect 8294 31288 8300 31300
rect 8352 31288 8358 31340
rect 8923 31327 8935 31361
rect 8969 31330 8984 31361
rect 9214 31356 9220 31368
rect 9272 31356 9278 31408
rect 10520 31368 11376 31396
rect 10520 31340 10548 31368
rect 8969 31327 8981 31330
rect 8923 31321 8981 31327
rect 10502 31288 10508 31340
rect 10560 31288 10566 31340
rect 11146 31288 11152 31340
rect 11204 31288 11210 31340
rect 11348 31328 11376 31368
rect 11759 31331 11817 31337
rect 11759 31328 11771 31331
rect 11348 31300 11771 31328
rect 11759 31297 11771 31300
rect 11805 31328 11817 31331
rect 11992 31328 12020 31424
rect 12158 31356 12164 31408
rect 12216 31396 12222 31408
rect 13357 31399 13415 31405
rect 13357 31396 13369 31399
rect 12216 31368 13369 31396
rect 12216 31356 12222 31368
rect 13357 31365 13369 31368
rect 13403 31365 13415 31399
rect 13357 31359 13415 31365
rect 13909 31399 13967 31405
rect 13909 31365 13921 31399
rect 13955 31396 13967 31399
rect 14274 31396 14280 31408
rect 13955 31368 14280 31396
rect 13955 31365 13967 31368
rect 13909 31359 13967 31365
rect 14274 31356 14280 31368
rect 14332 31356 14338 31408
rect 11805 31300 12020 31328
rect 13081 31331 13139 31337
rect 11805 31297 11817 31300
rect 11759 31291 11817 31297
rect 13081 31297 13093 31331
rect 13127 31328 13139 31331
rect 15378 31328 15384 31340
rect 13127 31300 15384 31328
rect 13127 31297 13139 31300
rect 13081 31291 13139 31297
rect 15378 31288 15384 31300
rect 15436 31288 15442 31340
rect 7285 31263 7343 31269
rect 7285 31229 7297 31263
rect 7331 31229 7343 31263
rect 8665 31263 8723 31269
rect 8665 31260 8677 31263
rect 7285 31223 7343 31229
rect 8220 31232 8677 31260
rect 1578 31084 1584 31136
rect 1636 31084 1642 31136
rect 7300 31124 7328 31223
rect 7558 31124 7564 31136
rect 7300 31096 7564 31124
rect 7558 31084 7564 31096
rect 7616 31124 7622 31136
rect 8220 31124 8248 31232
rect 8665 31229 8677 31232
rect 8711 31229 8723 31263
rect 11514 31260 11520 31272
rect 8665 31223 8723 31229
rect 9324 31232 11520 31260
rect 7616 31096 8248 31124
rect 7616 31084 7622 31096
rect 8294 31084 8300 31136
rect 8352 31084 8358 31136
rect 8680 31124 8708 31223
rect 9324 31124 9352 31232
rect 11514 31220 11520 31232
rect 11572 31220 11578 31272
rect 12250 31220 12256 31272
rect 12308 31260 12314 31272
rect 12308 31232 13584 31260
rect 12308 31220 12314 31232
rect 13262 31192 13268 31204
rect 12176 31164 13268 31192
rect 8680 31096 9352 31124
rect 9677 31127 9735 31133
rect 9677 31093 9689 31127
rect 9723 31124 9735 31127
rect 9858 31124 9864 31136
rect 9723 31096 9864 31124
rect 9723 31093 9735 31096
rect 9677 31087 9735 31093
rect 9858 31084 9864 31096
rect 9916 31084 9922 31136
rect 11790 31084 11796 31136
rect 11848 31124 11854 31136
rect 12176 31124 12204 31164
rect 13262 31152 13268 31164
rect 13320 31152 13326 31204
rect 13556 31136 13584 31232
rect 11848 31096 12204 31124
rect 11848 31084 11854 31096
rect 12250 31084 12256 31136
rect 12308 31124 12314 31136
rect 12529 31127 12587 31133
rect 12529 31124 12541 31127
rect 12308 31096 12541 31124
rect 12308 31084 12314 31096
rect 12529 31093 12541 31096
rect 12575 31093 12587 31127
rect 12529 31087 12587 31093
rect 12618 31084 12624 31136
rect 12676 31124 12682 31136
rect 12897 31127 12955 31133
rect 12897 31124 12909 31127
rect 12676 31096 12909 31124
rect 12676 31084 12682 31096
rect 12897 31093 12909 31096
rect 12943 31093 12955 31127
rect 12897 31087 12955 31093
rect 13538 31084 13544 31136
rect 13596 31084 13602 31136
rect 13630 31084 13636 31136
rect 13688 31084 13694 31136
rect 14185 31127 14243 31133
rect 14185 31093 14197 31127
rect 14231 31124 14243 31127
rect 15286 31124 15292 31136
rect 14231 31096 15292 31124
rect 14231 31093 14243 31096
rect 14185 31087 14243 31093
rect 15286 31084 15292 31096
rect 15344 31084 15350 31136
rect 1104 31034 14812 31056
rect 1104 30982 2663 31034
rect 2715 30982 2727 31034
rect 2779 30982 2791 31034
rect 2843 30982 2855 31034
rect 2907 30982 2919 31034
rect 2971 30982 6090 31034
rect 6142 30982 6154 31034
rect 6206 30982 6218 31034
rect 6270 30982 6282 31034
rect 6334 30982 6346 31034
rect 6398 30982 9517 31034
rect 9569 30982 9581 31034
rect 9633 30982 9645 31034
rect 9697 30982 9709 31034
rect 9761 30982 9773 31034
rect 9825 30982 12944 31034
rect 12996 30982 13008 31034
rect 13060 30982 13072 31034
rect 13124 30982 13136 31034
rect 13188 30982 13200 31034
rect 13252 30982 14812 31034
rect 1104 30960 14812 30982
rect 1578 30880 1584 30932
rect 1636 30920 1642 30932
rect 1636 30892 2774 30920
rect 1636 30880 1642 30892
rect 2746 30580 2774 30892
rect 5350 30880 5356 30932
rect 5408 30920 5414 30932
rect 5408 30892 9628 30920
rect 5408 30880 5414 30892
rect 9493 30855 9551 30861
rect 9493 30821 9505 30855
rect 9539 30821 9551 30855
rect 9600 30852 9628 30892
rect 10318 30880 10324 30932
rect 10376 30880 10382 30932
rect 10965 30923 11023 30929
rect 10965 30889 10977 30923
rect 11011 30920 11023 30923
rect 11146 30920 11152 30932
rect 11011 30892 11152 30920
rect 11011 30889 11023 30892
rect 10965 30883 11023 30889
rect 11146 30880 11152 30892
rect 11204 30880 11210 30932
rect 11514 30880 11520 30932
rect 11572 30880 11578 30932
rect 11790 30880 11796 30932
rect 11848 30880 11854 30932
rect 12066 30880 12072 30932
rect 12124 30880 12130 30932
rect 12618 30920 12624 30932
rect 12268 30892 12624 30920
rect 9600 30824 10640 30852
rect 9493 30815 9551 30821
rect 9508 30784 9536 30815
rect 10612 30784 10640 30824
rect 9508 30756 10548 30784
rect 10612 30756 12020 30784
rect 9674 30676 9680 30728
rect 9732 30676 9738 30728
rect 10520 30725 10548 30756
rect 10229 30719 10287 30725
rect 10229 30716 10241 30719
rect 9968 30688 10241 30716
rect 9968 30592 9996 30688
rect 10229 30685 10241 30688
rect 10275 30685 10287 30719
rect 10229 30679 10287 30685
rect 10505 30719 10563 30725
rect 10505 30685 10517 30719
rect 10551 30685 10563 30719
rect 10505 30679 10563 30685
rect 10870 30676 10876 30728
rect 10928 30676 10934 30728
rect 11992 30725 12020 30756
rect 12268 30725 12296 30892
rect 12618 30880 12624 30892
rect 12676 30880 12682 30932
rect 13446 30784 13452 30796
rect 12360 30756 13452 30784
rect 11149 30719 11207 30725
rect 11149 30685 11161 30719
rect 11195 30685 11207 30719
rect 11149 30679 11207 30685
rect 11701 30719 11759 30725
rect 11701 30685 11713 30719
rect 11747 30685 11759 30719
rect 11701 30679 11759 30685
rect 11977 30719 12035 30725
rect 11977 30685 11989 30719
rect 12023 30685 12035 30719
rect 11977 30679 12035 30685
rect 12253 30719 12311 30725
rect 12253 30685 12265 30719
rect 12299 30685 12311 30719
rect 12253 30679 12311 30685
rect 11164 30648 11192 30679
rect 10060 30620 11192 30648
rect 11716 30648 11744 30679
rect 12360 30648 12388 30756
rect 13446 30744 13452 30756
rect 13504 30744 13510 30796
rect 12434 30676 12440 30728
rect 12492 30676 12498 30728
rect 14185 30719 14243 30725
rect 14185 30716 14197 30719
rect 12636 30688 14197 30716
rect 12636 30648 12664 30688
rect 14185 30685 14197 30688
rect 14231 30685 14243 30719
rect 14185 30679 14243 30685
rect 11716 30620 12388 30648
rect 12452 30620 12664 30648
rect 12805 30651 12863 30657
rect 3786 30580 3792 30592
rect 2746 30552 3792 30580
rect 3786 30540 3792 30552
rect 3844 30540 3850 30592
rect 9950 30540 9956 30592
rect 10008 30540 10014 30592
rect 10060 30589 10088 30620
rect 10045 30583 10103 30589
rect 10045 30549 10057 30583
rect 10091 30549 10103 30583
rect 10045 30543 10103 30549
rect 10689 30583 10747 30589
rect 10689 30549 10701 30583
rect 10735 30580 10747 30583
rect 12452 30580 12480 30620
rect 12805 30617 12817 30651
rect 12851 30648 12863 30651
rect 12894 30648 12900 30660
rect 12851 30620 12900 30648
rect 12851 30617 12863 30620
rect 12805 30611 12863 30617
rect 12894 30608 12900 30620
rect 12952 30608 12958 30660
rect 12986 30608 12992 30660
rect 13044 30608 13050 30660
rect 13354 30608 13360 30660
rect 13412 30608 13418 30660
rect 13541 30651 13599 30657
rect 13541 30617 13553 30651
rect 13587 30617 13599 30651
rect 13541 30611 13599 30617
rect 13909 30651 13967 30657
rect 13909 30617 13921 30651
rect 13955 30648 13967 30651
rect 14550 30648 14556 30660
rect 13955 30620 14556 30648
rect 13955 30617 13967 30620
rect 13909 30611 13967 30617
rect 10735 30552 12480 30580
rect 10735 30549 10747 30552
rect 10689 30543 10747 30549
rect 12710 30540 12716 30592
rect 12768 30580 12774 30592
rect 13556 30580 13584 30611
rect 14550 30608 14556 30620
rect 14608 30608 14614 30660
rect 12768 30552 13584 30580
rect 14369 30583 14427 30589
rect 12768 30540 12774 30552
rect 14369 30549 14381 30583
rect 14415 30580 14427 30583
rect 15102 30580 15108 30592
rect 14415 30552 15108 30580
rect 14415 30549 14427 30552
rect 14369 30543 14427 30549
rect 15102 30540 15108 30552
rect 15160 30540 15166 30592
rect 1104 30490 14971 30512
rect 1104 30438 4376 30490
rect 4428 30438 4440 30490
rect 4492 30438 4504 30490
rect 4556 30438 4568 30490
rect 4620 30438 4632 30490
rect 4684 30438 7803 30490
rect 7855 30438 7867 30490
rect 7919 30438 7931 30490
rect 7983 30438 7995 30490
rect 8047 30438 8059 30490
rect 8111 30438 11230 30490
rect 11282 30438 11294 30490
rect 11346 30438 11358 30490
rect 11410 30438 11422 30490
rect 11474 30438 11486 30490
rect 11538 30438 14657 30490
rect 14709 30438 14721 30490
rect 14773 30438 14785 30490
rect 14837 30438 14849 30490
rect 14901 30438 14913 30490
rect 14965 30438 14971 30490
rect 1104 30416 14971 30438
rect 7098 30336 7104 30388
rect 7156 30376 7162 30388
rect 9122 30376 9128 30388
rect 7156 30348 9128 30376
rect 7156 30336 7162 30348
rect 9122 30336 9128 30348
rect 9180 30336 9186 30388
rect 13449 30379 13507 30385
rect 13449 30345 13461 30379
rect 13495 30376 13507 30379
rect 13722 30376 13728 30388
rect 13495 30348 13728 30376
rect 13495 30345 13507 30348
rect 13449 30339 13507 30345
rect 13722 30336 13728 30348
rect 13780 30336 13786 30388
rect 6822 30308 6828 30320
rect 6380 30280 6828 30308
rect 750 30200 756 30252
rect 808 30240 814 30252
rect 6380 30249 6408 30280
rect 6822 30268 6828 30280
rect 6880 30308 6886 30320
rect 7190 30308 7196 30320
rect 6880 30280 7196 30308
rect 6880 30268 6886 30280
rect 7190 30268 7196 30280
rect 7248 30268 7254 30320
rect 8478 30268 8484 30320
rect 8536 30308 8542 30320
rect 8536 30280 9260 30308
rect 8536 30268 8542 30280
rect 1397 30243 1455 30249
rect 1397 30240 1409 30243
rect 808 30212 1409 30240
rect 808 30200 814 30212
rect 1397 30209 1409 30212
rect 1443 30209 1455 30243
rect 1397 30203 1455 30209
rect 6365 30243 6423 30249
rect 6365 30209 6377 30243
rect 6411 30209 6423 30243
rect 6365 30203 6423 30209
rect 6639 30243 6697 30249
rect 6639 30209 6651 30243
rect 6685 30240 6697 30243
rect 7006 30240 7012 30252
rect 6685 30212 7012 30240
rect 6685 30209 6697 30212
rect 6639 30203 6697 30209
rect 7006 30200 7012 30212
rect 7064 30240 7070 30252
rect 7374 30240 7380 30252
rect 7064 30212 7380 30240
rect 7064 30200 7070 30212
rect 7374 30200 7380 30212
rect 7432 30200 7438 30252
rect 9125 30243 9183 30249
rect 9125 30240 9137 30243
rect 9048 30212 9137 30240
rect 9048 30184 9076 30212
rect 9125 30209 9137 30212
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 9030 30132 9036 30184
rect 9088 30132 9094 30184
rect 9232 30181 9260 30280
rect 10410 30200 10416 30252
rect 10468 30200 10474 30252
rect 12802 30200 12808 30252
rect 12860 30200 12866 30252
rect 13998 30200 14004 30252
rect 14056 30200 14062 30252
rect 9217 30175 9275 30181
rect 9217 30141 9229 30175
rect 9263 30141 9275 30175
rect 9217 30135 9275 30141
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 9401 30175 9459 30181
rect 9401 30172 9413 30175
rect 9364 30144 9413 30172
rect 9364 30132 9370 30144
rect 9401 30141 9413 30144
rect 9447 30141 9459 30175
rect 9401 30135 9459 30141
rect 9766 30132 9772 30184
rect 9824 30132 9830 30184
rect 9858 30132 9864 30184
rect 9916 30132 9922 30184
rect 10318 30181 10324 30184
rect 10137 30175 10195 30181
rect 10137 30172 10149 30175
rect 9968 30144 10149 30172
rect 1581 30107 1639 30113
rect 1581 30073 1593 30107
rect 1627 30104 1639 30107
rect 3878 30104 3884 30116
rect 1627 30076 3884 30104
rect 1627 30073 1639 30076
rect 1581 30067 1639 30073
rect 3878 30064 3884 30076
rect 3936 30064 3942 30116
rect 8941 30107 8999 30113
rect 7300 30076 8892 30104
rect 2406 29996 2412 30048
rect 2464 30036 2470 30048
rect 7300 30036 7328 30076
rect 2464 30008 7328 30036
rect 2464 29996 2470 30008
rect 7374 29996 7380 30048
rect 7432 29996 7438 30048
rect 8864 30036 8892 30076
rect 8941 30073 8953 30107
rect 8987 30104 8999 30107
rect 9674 30104 9680 30116
rect 8987 30076 9680 30104
rect 8987 30073 8999 30076
rect 8941 30067 8999 30073
rect 9674 30064 9680 30076
rect 9732 30064 9738 30116
rect 9784 30104 9812 30132
rect 9968 30104 9996 30144
rect 10137 30141 10149 30144
rect 10183 30141 10195 30175
rect 10137 30135 10195 30141
rect 10275 30175 10324 30181
rect 10275 30141 10287 30175
rect 10321 30141 10324 30175
rect 10275 30135 10324 30141
rect 10318 30132 10324 30135
rect 10376 30132 10382 30184
rect 11606 30132 11612 30184
rect 11664 30132 11670 30184
rect 11790 30132 11796 30184
rect 11848 30132 11854 30184
rect 12529 30175 12587 30181
rect 12529 30172 12541 30175
rect 12084 30144 12541 30172
rect 11882 30104 11888 30116
rect 9784 30076 9996 30104
rect 10980 30076 11888 30104
rect 10980 30036 11008 30076
rect 11882 30064 11888 30076
rect 11940 30064 11946 30116
rect 12084 30048 12112 30144
rect 12529 30141 12541 30144
rect 12575 30141 12587 30175
rect 12529 30135 12587 30141
rect 12667 30175 12725 30181
rect 12667 30141 12679 30175
rect 12713 30172 12725 30175
rect 13354 30172 13360 30184
rect 12713 30144 13360 30172
rect 12713 30141 12725 30144
rect 12667 30135 12725 30141
rect 13354 30132 13360 30144
rect 13412 30132 13418 30184
rect 12253 30107 12311 30113
rect 12253 30073 12265 30107
rect 12299 30073 12311 30107
rect 12253 30067 12311 30073
rect 13817 30107 13875 30113
rect 13817 30073 13829 30107
rect 13863 30104 13875 30107
rect 13906 30104 13912 30116
rect 13863 30076 13912 30104
rect 13863 30073 13875 30076
rect 13817 30067 13875 30073
rect 8864 30008 11008 30036
rect 11054 29996 11060 30048
rect 11112 29996 11118 30048
rect 12066 29996 12072 30048
rect 12124 29996 12130 30048
rect 12268 30036 12296 30067
rect 13906 30064 13912 30076
rect 13964 30104 13970 30116
rect 13964 30076 15792 30104
rect 13964 30064 13970 30076
rect 15764 30048 15792 30076
rect 12618 30036 12624 30048
rect 12268 30008 12624 30036
rect 12618 29996 12624 30008
rect 12676 29996 12682 30048
rect 14274 29996 14280 30048
rect 14332 29996 14338 30048
rect 15746 29996 15752 30048
rect 15804 29996 15810 30048
rect 1104 29946 14812 29968
rect 1104 29894 2663 29946
rect 2715 29894 2727 29946
rect 2779 29894 2791 29946
rect 2843 29894 2855 29946
rect 2907 29894 2919 29946
rect 2971 29894 6090 29946
rect 6142 29894 6154 29946
rect 6206 29894 6218 29946
rect 6270 29894 6282 29946
rect 6334 29894 6346 29946
rect 6398 29894 9517 29946
rect 9569 29894 9581 29946
rect 9633 29894 9645 29946
rect 9697 29894 9709 29946
rect 9761 29894 9773 29946
rect 9825 29894 12944 29946
rect 12996 29894 13008 29946
rect 13060 29894 13072 29946
rect 13124 29894 13136 29946
rect 13188 29894 13200 29946
rect 13252 29894 14812 29946
rect 1104 29872 14812 29894
rect 1581 29835 1639 29841
rect 1581 29801 1593 29835
rect 1627 29832 1639 29835
rect 2038 29832 2044 29844
rect 1627 29804 2044 29832
rect 1627 29801 1639 29804
rect 1581 29795 1639 29801
rect 2038 29792 2044 29804
rect 2096 29832 2102 29844
rect 2406 29832 2412 29844
rect 2096 29804 2412 29832
rect 2096 29792 2102 29804
rect 2406 29792 2412 29804
rect 2464 29792 2470 29844
rect 7374 29792 7380 29844
rect 7432 29832 7438 29844
rect 7432 29804 7604 29832
rect 7432 29792 7438 29804
rect 7576 29773 7604 29804
rect 8294 29792 8300 29844
rect 8352 29832 8358 29844
rect 10781 29835 10839 29841
rect 8352 29804 9628 29832
rect 8352 29792 8358 29804
rect 7561 29767 7619 29773
rect 7561 29733 7573 29767
rect 7607 29733 7619 29767
rect 7561 29727 7619 29733
rect 8754 29724 8760 29776
rect 8812 29724 8818 29776
rect 8938 29724 8944 29776
rect 8996 29764 9002 29776
rect 9600 29773 9628 29804
rect 9692 29804 10548 29832
rect 9585 29767 9643 29773
rect 8996 29736 9352 29764
rect 8996 29724 9002 29736
rect 4246 29656 4252 29708
rect 4304 29696 4310 29708
rect 5534 29696 5540 29708
rect 4304 29668 5540 29696
rect 4304 29656 4310 29668
rect 5534 29656 5540 29668
rect 5592 29656 5598 29708
rect 7650 29656 7656 29708
rect 7708 29696 7714 29708
rect 7954 29699 8012 29705
rect 7954 29696 7966 29699
rect 7708 29668 7966 29696
rect 7708 29656 7714 29668
rect 7954 29665 7966 29668
rect 8000 29665 8012 29699
rect 7954 29659 8012 29665
rect 9125 29699 9183 29705
rect 9125 29665 9137 29699
rect 9171 29696 9183 29699
rect 9214 29696 9220 29708
rect 9171 29668 9220 29696
rect 9171 29665 9183 29668
rect 9125 29659 9183 29665
rect 9214 29656 9220 29668
rect 9272 29656 9278 29708
rect 9324 29696 9352 29736
rect 9585 29733 9597 29767
rect 9631 29733 9643 29767
rect 9585 29727 9643 29733
rect 9692 29696 9720 29804
rect 9324 29668 9720 29696
rect 10137 29699 10195 29705
rect 10137 29665 10149 29699
rect 10183 29696 10195 29699
rect 10520 29696 10548 29804
rect 10781 29801 10793 29835
rect 10827 29832 10839 29835
rect 10870 29832 10876 29844
rect 10827 29804 10876 29832
rect 10827 29801 10839 29804
rect 10781 29795 10839 29801
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 11054 29792 11060 29844
rect 11112 29792 11118 29844
rect 11333 29835 11391 29841
rect 11333 29801 11345 29835
rect 11379 29832 11391 29835
rect 12158 29832 12164 29844
rect 11379 29804 12164 29832
rect 11379 29801 11391 29804
rect 11333 29795 11391 29801
rect 12158 29792 12164 29804
rect 12216 29792 12222 29844
rect 13446 29792 13452 29844
rect 13504 29792 13510 29844
rect 10183 29668 10548 29696
rect 11072 29696 11100 29792
rect 12250 29724 12256 29776
rect 12308 29724 12314 29776
rect 13814 29724 13820 29776
rect 13872 29724 13878 29776
rect 11793 29699 11851 29705
rect 11072 29668 11560 29696
rect 10183 29665 10195 29668
rect 10137 29659 10195 29665
rect 750 29588 756 29640
rect 808 29628 814 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 808 29600 1409 29628
rect 808 29588 814 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 5810 29628 5816 29640
rect 1397 29591 1455 29597
rect 5644 29600 5816 29628
rect 3878 29520 3884 29572
rect 3936 29560 3942 29572
rect 5644 29560 5672 29600
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 6822 29588 6828 29640
rect 6880 29628 6886 29640
rect 6917 29631 6975 29637
rect 6917 29628 6929 29631
rect 6880 29600 6929 29628
rect 6880 29588 6886 29600
rect 6917 29597 6929 29600
rect 6963 29597 6975 29631
rect 6917 29591 6975 29597
rect 7101 29631 7159 29637
rect 7101 29597 7113 29631
rect 7147 29597 7159 29631
rect 7101 29591 7159 29597
rect 3936 29532 5672 29560
rect 3936 29520 3942 29532
rect 6546 29452 6552 29504
rect 6604 29452 6610 29504
rect 6730 29452 6736 29504
rect 6788 29492 6794 29504
rect 7116 29492 7144 29591
rect 7834 29588 7840 29640
rect 7892 29588 7898 29640
rect 8110 29588 8116 29640
rect 8168 29588 8174 29640
rect 8938 29588 8944 29640
rect 8996 29588 9002 29640
rect 9858 29588 9864 29640
rect 9916 29588 9922 29640
rect 10042 29637 10048 29640
rect 9999 29631 10048 29637
rect 9999 29597 10011 29631
rect 10045 29597 10048 29631
rect 9999 29591 10048 29597
rect 10042 29588 10048 29591
rect 10100 29588 10106 29640
rect 11054 29588 11060 29640
rect 11112 29588 11118 29640
rect 11532 29637 11560 29668
rect 11793 29665 11805 29699
rect 11839 29665 11851 29699
rect 11793 29659 11851 29665
rect 11517 29631 11575 29637
rect 11517 29597 11529 29631
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11606 29588 11612 29640
rect 11664 29588 11670 29640
rect 11808 29572 11836 29659
rect 12158 29656 12164 29708
rect 12216 29696 12222 29708
rect 12529 29699 12587 29705
rect 12529 29696 12541 29699
rect 12216 29668 12541 29696
rect 12216 29656 12222 29668
rect 12529 29665 12541 29668
rect 12575 29665 12587 29699
rect 12529 29659 12587 29665
rect 12805 29699 12863 29705
rect 12805 29665 12817 29699
rect 12851 29696 12863 29699
rect 13832 29696 13860 29724
rect 12851 29668 13860 29696
rect 12851 29665 12863 29668
rect 12805 29659 12863 29665
rect 12618 29588 12624 29640
rect 12676 29637 12682 29640
rect 12676 29631 12704 29637
rect 12692 29597 12704 29631
rect 12676 29591 12704 29597
rect 13725 29631 13783 29637
rect 13725 29597 13737 29631
rect 13771 29597 13783 29631
rect 13725 29591 13783 29597
rect 12676 29588 12682 29591
rect 11790 29520 11796 29572
rect 11848 29520 11854 29572
rect 13740 29560 13768 29591
rect 13814 29588 13820 29640
rect 13872 29628 13878 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 13872 29600 14289 29628
rect 13872 29588 13878 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 14366 29560 14372 29572
rect 13740 29532 14372 29560
rect 14366 29520 14372 29532
rect 14424 29520 14430 29572
rect 10042 29492 10048 29504
rect 6788 29464 10048 29492
rect 6788 29452 6794 29464
rect 10042 29452 10048 29464
rect 10100 29492 10106 29504
rect 10410 29492 10416 29504
rect 10100 29464 10416 29492
rect 10100 29452 10106 29464
rect 10410 29452 10416 29464
rect 10468 29452 10474 29504
rect 10873 29495 10931 29501
rect 10873 29461 10885 29495
rect 10919 29492 10931 29495
rect 12434 29492 12440 29504
rect 10919 29464 12440 29492
rect 10919 29461 10931 29464
rect 10873 29455 10931 29461
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 13541 29495 13599 29501
rect 13541 29461 13553 29495
rect 13587 29492 13599 29495
rect 13906 29492 13912 29504
rect 13587 29464 13912 29492
rect 13587 29461 13599 29464
rect 13541 29455 13599 29461
rect 13906 29452 13912 29464
rect 13964 29452 13970 29504
rect 14090 29452 14096 29504
rect 14148 29452 14154 29504
rect 1104 29402 14971 29424
rect 1104 29350 4376 29402
rect 4428 29350 4440 29402
rect 4492 29350 4504 29402
rect 4556 29350 4568 29402
rect 4620 29350 4632 29402
rect 4684 29350 7803 29402
rect 7855 29350 7867 29402
rect 7919 29350 7931 29402
rect 7983 29350 7995 29402
rect 8047 29350 8059 29402
rect 8111 29350 11230 29402
rect 11282 29350 11294 29402
rect 11346 29350 11358 29402
rect 11410 29350 11422 29402
rect 11474 29350 11486 29402
rect 11538 29350 14657 29402
rect 14709 29350 14721 29402
rect 14773 29350 14785 29402
rect 14837 29350 14849 29402
rect 14901 29350 14913 29402
rect 14965 29350 14971 29402
rect 1104 29328 14971 29350
rect 6546 29248 6552 29300
rect 6604 29248 6610 29300
rect 8294 29248 8300 29300
rect 8352 29288 8358 29300
rect 9858 29288 9864 29300
rect 8352 29260 9864 29288
rect 8352 29248 8358 29260
rect 6564 29152 6592 29248
rect 6564 29124 7142 29152
rect 6730 29044 6736 29096
rect 6788 29044 6794 29096
rect 6822 29044 6828 29096
rect 6880 29044 6886 29096
rect 7009 29087 7067 29093
rect 7009 29053 7021 29087
rect 7055 29053 7067 29087
rect 7114 29084 7142 29124
rect 7834 29112 7840 29164
rect 7892 29161 7898 29164
rect 7892 29155 7920 29161
rect 7908 29121 7920 29155
rect 7892 29115 7920 29121
rect 7892 29112 7898 29115
rect 8018 29112 8024 29164
rect 8076 29112 8082 29164
rect 7469 29087 7527 29093
rect 7469 29084 7481 29087
rect 7114 29056 7481 29084
rect 7009 29047 7067 29053
rect 7469 29053 7481 29056
rect 7515 29053 7527 29087
rect 7469 29047 7527 29053
rect 7745 29087 7803 29093
rect 7745 29053 7757 29087
rect 7791 29084 7803 29087
rect 8588 29084 8616 29260
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 12069 29291 12127 29297
rect 12069 29257 12081 29291
rect 12115 29288 12127 29291
rect 12115 29260 12434 29288
rect 12115 29257 12127 29260
rect 12069 29251 12127 29257
rect 8665 29223 8723 29229
rect 8665 29189 8677 29223
rect 8711 29220 8723 29223
rect 12406 29220 12434 29260
rect 12710 29248 12716 29300
rect 12768 29248 12774 29300
rect 12802 29248 12808 29300
rect 12860 29248 12866 29300
rect 12989 29291 13047 29297
rect 12989 29257 13001 29291
rect 13035 29288 13047 29291
rect 13035 29260 13400 29288
rect 13035 29257 13047 29260
rect 12989 29251 13047 29257
rect 12820 29220 12848 29248
rect 13372 29229 13400 29260
rect 8711 29192 12020 29220
rect 12406 29192 12848 29220
rect 13357 29223 13415 29229
rect 8711 29189 8723 29192
rect 8665 29183 8723 29189
rect 9030 29161 9036 29164
rect 8999 29155 9036 29161
rect 8999 29152 9011 29155
rect 7791 29056 8616 29084
rect 8680 29124 9011 29152
rect 7791 29053 7803 29056
rect 7745 29047 7803 29053
rect 5258 28976 5264 29028
rect 5316 29016 5322 29028
rect 6748 29016 6776 29044
rect 7024 29016 7052 29047
rect 8680 29028 8708 29124
rect 8999 29121 9011 29124
rect 8999 29115 9036 29121
rect 9030 29112 9036 29115
rect 9088 29112 9094 29164
rect 11790 29152 11796 29164
rect 9416 29124 11796 29152
rect 8754 29044 8760 29096
rect 8812 29044 8818 29096
rect 5316 28988 6684 29016
rect 6748 28988 7052 29016
rect 5316 28976 5322 28988
rect 6656 28948 6684 28988
rect 8662 28976 8668 29028
rect 8720 28976 8726 29028
rect 9416 28948 9444 29124
rect 11790 29112 11796 29124
rect 11848 29112 11854 29164
rect 11992 29161 12020 29192
rect 13357 29189 13369 29223
rect 13403 29189 13415 29223
rect 13357 29183 13415 29189
rect 13909 29223 13967 29229
rect 13909 29189 13921 29223
rect 13955 29220 13967 29223
rect 14182 29220 14188 29232
rect 13955 29192 14188 29220
rect 13955 29189 13967 29192
rect 13909 29183 13967 29189
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 12253 29155 12311 29161
rect 12253 29121 12265 29155
rect 12299 29121 12311 29155
rect 12253 29115 12311 29121
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 11882 29044 11888 29096
rect 11940 29084 11946 29096
rect 12268 29084 12296 29115
rect 11940 29056 12296 29084
rect 12636 29084 12664 29115
rect 12894 29112 12900 29164
rect 12952 29112 12958 29164
rect 12986 29112 12992 29164
rect 13044 29152 13050 29164
rect 13173 29155 13231 29161
rect 13173 29152 13185 29155
rect 13044 29124 13185 29152
rect 13044 29112 13050 29124
rect 13173 29121 13185 29124
rect 13219 29121 13231 29155
rect 13173 29115 13231 29121
rect 13998 29112 14004 29164
rect 14056 29112 14062 29164
rect 13262 29084 13268 29096
rect 12636 29056 13268 29084
rect 11940 29044 11946 29056
rect 13262 29044 13268 29056
rect 13320 29044 13326 29096
rect 11790 28976 11796 29028
rect 11848 28976 11854 29028
rect 12437 29019 12495 29025
rect 12437 28985 12449 29019
rect 12483 29016 12495 29019
rect 14016 29016 14044 29112
rect 12483 28988 14044 29016
rect 12483 28985 12495 28988
rect 12437 28979 12495 28985
rect 6656 28920 9444 28948
rect 9769 28951 9827 28957
rect 9769 28917 9781 28951
rect 9815 28948 9827 28951
rect 10134 28948 10140 28960
rect 9815 28920 10140 28948
rect 9815 28917 9827 28920
rect 9769 28911 9827 28917
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 10686 28908 10692 28960
rect 10744 28948 10750 28960
rect 12250 28948 12256 28960
rect 10744 28920 12256 28948
rect 10744 28908 10750 28920
rect 12250 28908 12256 28920
rect 12308 28908 12314 28960
rect 13630 28908 13636 28960
rect 13688 28908 13694 28960
rect 14182 28908 14188 28960
rect 14240 28908 14246 28960
rect 1104 28858 14812 28880
rect 1104 28806 2663 28858
rect 2715 28806 2727 28858
rect 2779 28806 2791 28858
rect 2843 28806 2855 28858
rect 2907 28806 2919 28858
rect 2971 28806 6090 28858
rect 6142 28806 6154 28858
rect 6206 28806 6218 28858
rect 6270 28806 6282 28858
rect 6334 28806 6346 28858
rect 6398 28806 9517 28858
rect 9569 28806 9581 28858
rect 9633 28806 9645 28858
rect 9697 28806 9709 28858
rect 9761 28806 9773 28858
rect 9825 28806 12944 28858
rect 12996 28806 13008 28858
rect 13060 28806 13072 28858
rect 13124 28806 13136 28858
rect 13188 28806 13200 28858
rect 13252 28806 14812 28858
rect 1104 28784 14812 28806
rect 5534 28704 5540 28756
rect 5592 28744 5598 28756
rect 5994 28744 6000 28756
rect 5592 28716 6000 28744
rect 5592 28704 5598 28716
rect 5994 28704 6000 28716
rect 6052 28744 6058 28756
rect 7653 28747 7711 28753
rect 6052 28716 7326 28744
rect 6052 28704 6058 28716
rect 6702 28676 6730 28716
rect 6656 28648 6730 28676
rect 7298 28676 7326 28716
rect 7653 28713 7665 28747
rect 7699 28744 7711 28747
rect 8018 28744 8024 28756
rect 7699 28716 8024 28744
rect 7699 28713 7711 28716
rect 7653 28707 7711 28713
rect 8018 28704 8024 28716
rect 8076 28704 8082 28756
rect 10778 28704 10784 28756
rect 10836 28744 10842 28756
rect 10836 28716 12204 28744
rect 10836 28704 10842 28716
rect 8754 28676 8760 28688
rect 7298 28648 8760 28676
rect 6656 28617 6684 28648
rect 8754 28636 8760 28648
rect 8812 28676 8818 28688
rect 8812 28648 9674 28676
rect 8812 28636 8818 28648
rect 9646 28620 9674 28648
rect 10134 28636 10140 28688
rect 10192 28676 10198 28688
rect 10413 28679 10471 28685
rect 10413 28676 10425 28679
rect 10192 28648 10425 28676
rect 10192 28636 10198 28648
rect 10413 28645 10425 28648
rect 10459 28645 10471 28679
rect 10413 28639 10471 28645
rect 6641 28611 6699 28617
rect 6641 28577 6653 28611
rect 6687 28577 6699 28611
rect 9646 28580 9680 28620
rect 6641 28571 6699 28577
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 9769 28611 9827 28617
rect 9769 28577 9781 28611
rect 9815 28608 9827 28611
rect 10318 28608 10324 28620
rect 9815 28580 10324 28608
rect 9815 28577 9827 28580
rect 9769 28571 9827 28577
rect 10318 28568 10324 28580
rect 10376 28608 10382 28620
rect 11701 28611 11759 28617
rect 11701 28608 11713 28611
rect 10376 28580 11713 28608
rect 10376 28568 10382 28580
rect 11701 28577 11713 28580
rect 11747 28608 11759 28611
rect 12176 28608 12204 28716
rect 12250 28704 12256 28756
rect 12308 28744 12314 28756
rect 12618 28744 12624 28756
rect 12308 28716 12624 28744
rect 12308 28704 12314 28716
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 13541 28747 13599 28753
rect 13541 28713 13553 28747
rect 13587 28744 13599 28747
rect 13814 28744 13820 28756
rect 13587 28716 13820 28744
rect 13587 28713 13599 28716
rect 13541 28707 13599 28713
rect 13814 28704 13820 28716
rect 13872 28704 13878 28756
rect 12342 28636 12348 28688
rect 12400 28636 12406 28688
rect 12738 28611 12796 28617
rect 12738 28608 12750 28611
rect 11747 28580 12112 28608
rect 12176 28580 12750 28608
rect 11747 28577 11759 28580
rect 11701 28571 11759 28577
rect 12084 28552 12112 28580
rect 12738 28577 12750 28580
rect 12784 28577 12796 28611
rect 12738 28571 12796 28577
rect 750 28500 756 28552
rect 808 28540 814 28552
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 808 28512 1409 28540
rect 808 28500 814 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 6899 28543 6957 28549
rect 6899 28540 6911 28543
rect 1397 28503 1455 28509
rect 6840 28512 6911 28540
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 3786 28364 3792 28416
rect 3844 28404 3850 28416
rect 6840 28404 6868 28512
rect 6899 28509 6911 28512
rect 6945 28509 6957 28543
rect 6899 28503 6957 28509
rect 8846 28500 8852 28552
rect 8904 28540 8910 28552
rect 9953 28543 10011 28549
rect 9953 28540 9965 28543
rect 8904 28512 9965 28540
rect 8904 28500 8910 28512
rect 9953 28509 9965 28512
rect 9999 28509 10011 28543
rect 9953 28503 10011 28509
rect 7098 28404 7104 28416
rect 3844 28376 7104 28404
rect 3844 28364 3850 28376
rect 7098 28364 7104 28376
rect 7156 28364 7162 28416
rect 9968 28404 9996 28503
rect 10686 28500 10692 28552
rect 10744 28500 10750 28552
rect 10778 28500 10784 28552
rect 10836 28549 10842 28552
rect 10836 28543 10864 28549
rect 10852 28509 10864 28543
rect 10836 28503 10864 28509
rect 10836 28500 10842 28503
rect 10962 28500 10968 28552
rect 11020 28500 11026 28552
rect 11885 28543 11943 28549
rect 11885 28509 11897 28543
rect 11931 28509 11943 28543
rect 11885 28503 11943 28509
rect 11900 28472 11928 28503
rect 12066 28500 12072 28552
rect 12124 28500 12130 28552
rect 12618 28500 12624 28552
rect 12676 28500 12682 28552
rect 12894 28500 12900 28552
rect 12952 28500 12958 28552
rect 13538 28500 13544 28552
rect 13596 28540 13602 28552
rect 13633 28543 13691 28549
rect 13633 28540 13645 28543
rect 13596 28512 13645 28540
rect 13596 28500 13602 28512
rect 13633 28509 13645 28512
rect 13679 28509 13691 28543
rect 13633 28503 13691 28509
rect 13998 28500 14004 28552
rect 14056 28540 14062 28552
rect 14185 28543 14243 28549
rect 14185 28540 14197 28543
rect 14056 28512 14197 28540
rect 14056 28500 14062 28512
rect 14185 28509 14197 28512
rect 14231 28509 14243 28543
rect 14185 28503 14243 28509
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 14550 28540 14556 28552
rect 14424 28512 14556 28540
rect 14424 28500 14430 28512
rect 14550 28500 14556 28512
rect 14608 28500 14614 28552
rect 11440 28444 11928 28472
rect 11440 28404 11468 28444
rect 9968 28376 11468 28404
rect 11609 28407 11667 28413
rect 11609 28373 11621 28407
rect 11655 28404 11667 28407
rect 12342 28404 12348 28416
rect 11655 28376 12348 28404
rect 11655 28373 11667 28376
rect 11609 28367 11667 28373
rect 12342 28364 12348 28376
rect 12400 28364 12406 28416
rect 13814 28364 13820 28416
rect 13872 28364 13878 28416
rect 14366 28364 14372 28416
rect 14424 28364 14430 28416
rect 1104 28314 14971 28336
rect 1104 28262 4376 28314
rect 4428 28262 4440 28314
rect 4492 28262 4504 28314
rect 4556 28262 4568 28314
rect 4620 28262 4632 28314
rect 4684 28262 7803 28314
rect 7855 28262 7867 28314
rect 7919 28262 7931 28314
rect 7983 28262 7995 28314
rect 8047 28262 8059 28314
rect 8111 28262 11230 28314
rect 11282 28262 11294 28314
rect 11346 28262 11358 28314
rect 11410 28262 11422 28314
rect 11474 28262 11486 28314
rect 11538 28262 14657 28314
rect 14709 28262 14721 28314
rect 14773 28262 14785 28314
rect 14837 28262 14849 28314
rect 14901 28262 14913 28314
rect 14965 28262 14971 28314
rect 1104 28240 14971 28262
rect 1578 28160 1584 28212
rect 1636 28200 1642 28212
rect 1946 28200 1952 28212
rect 1636 28172 1952 28200
rect 1636 28160 1642 28172
rect 1946 28160 1952 28172
rect 2004 28200 2010 28212
rect 10134 28200 10140 28212
rect 2004 28172 10140 28200
rect 2004 28160 2010 28172
rect 10134 28160 10140 28172
rect 10192 28200 10198 28212
rect 10502 28200 10508 28212
rect 10192 28172 10508 28200
rect 10192 28160 10198 28172
rect 10502 28160 10508 28172
rect 10560 28160 10566 28212
rect 10689 28203 10747 28209
rect 10689 28169 10701 28203
rect 10735 28200 10747 28203
rect 10962 28200 10968 28212
rect 10735 28172 10968 28200
rect 10735 28169 10747 28172
rect 10689 28163 10747 28169
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11698 28160 11704 28212
rect 11756 28200 11762 28212
rect 12713 28203 12771 28209
rect 11756 28172 12434 28200
rect 11756 28160 11762 28172
rect 9766 28092 9772 28144
rect 9824 28132 9830 28144
rect 10870 28132 10876 28144
rect 9824 28104 10876 28132
rect 9824 28092 9830 28104
rect 10870 28092 10876 28104
rect 10928 28132 10934 28144
rect 10928 28104 11744 28132
rect 10928 28092 10934 28104
rect 1486 28024 1492 28076
rect 1544 28024 1550 28076
rect 7558 28024 7564 28076
rect 7616 28064 7622 28076
rect 8021 28067 8079 28073
rect 8021 28064 8033 28067
rect 7616 28036 8033 28064
rect 7616 28024 7622 28036
rect 8021 28033 8033 28036
rect 8067 28064 8079 28067
rect 8202 28064 8208 28076
rect 8067 28036 8208 28064
rect 8067 28033 8079 28036
rect 8021 28027 8079 28033
rect 8202 28024 8208 28036
rect 8260 28024 8266 28076
rect 8295 28067 8353 28073
rect 8295 28033 8307 28067
rect 8341 28064 8353 28067
rect 9784 28064 9812 28092
rect 8341 28036 9260 28064
rect 8341 28033 8353 28036
rect 8295 28027 8353 28033
rect 1581 27863 1639 27869
rect 1581 27829 1593 27863
rect 1627 27860 1639 27863
rect 1670 27860 1676 27872
rect 1627 27832 1676 27860
rect 1627 27829 1639 27832
rect 1581 27823 1639 27829
rect 1670 27820 1676 27832
rect 1728 27860 1734 27872
rect 6638 27860 6644 27872
rect 1728 27832 6644 27860
rect 1728 27820 1734 27832
rect 6638 27820 6644 27832
rect 6696 27860 6702 27872
rect 8386 27860 8392 27872
rect 6696 27832 8392 27860
rect 6696 27820 6702 27832
rect 8386 27820 8392 27832
rect 8444 27820 8450 27872
rect 9033 27863 9091 27869
rect 9033 27829 9045 27863
rect 9079 27860 9091 27863
rect 9122 27860 9128 27872
rect 9079 27832 9128 27860
rect 9079 27829 9091 27832
rect 9033 27823 9091 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 9232 27860 9260 28036
rect 9692 28036 9812 28064
rect 9692 28005 9720 28036
rect 9858 28024 9864 28076
rect 9916 28064 9922 28076
rect 9951 28067 10009 28073
rect 9951 28064 9963 28067
rect 9916 28036 9963 28064
rect 9916 28024 9922 28036
rect 9951 28033 9963 28036
rect 9997 28033 10009 28067
rect 9951 28027 10009 28033
rect 11716 28008 11744 28104
rect 11974 28103 11980 28144
rect 11959 28097 11980 28103
rect 11959 28063 11971 28097
rect 12032 28092 12038 28144
rect 12406 28132 12434 28172
rect 12713 28169 12725 28203
rect 12759 28200 12771 28203
rect 12894 28200 12900 28212
rect 12759 28172 12900 28200
rect 12759 28169 12771 28172
rect 12713 28163 12771 28169
rect 12894 28160 12900 28172
rect 12952 28160 12958 28212
rect 14274 28200 14280 28212
rect 13004 28172 14280 28200
rect 13004 28132 13032 28172
rect 14274 28160 14280 28172
rect 14332 28160 14338 28212
rect 12406 28104 13032 28132
rect 13906 28092 13912 28144
rect 13964 28092 13970 28144
rect 12005 28066 12020 28092
rect 12005 28063 12017 28066
rect 11959 28057 12017 28063
rect 12066 28024 12072 28076
rect 12124 28064 12130 28076
rect 12124 28036 12434 28064
rect 12124 28024 12130 28036
rect 9677 27999 9735 28005
rect 9677 27965 9689 27999
rect 9723 27965 9735 27999
rect 9677 27959 9735 27965
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 12406 27928 12434 28036
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 13357 28067 13415 28073
rect 13357 28064 13369 28067
rect 12676 28036 13369 28064
rect 12676 28024 12682 28036
rect 13357 28033 13369 28036
rect 13403 28033 13415 28067
rect 13357 28027 13415 28033
rect 15102 27928 15108 27940
rect 12406 27900 15108 27928
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 10042 27860 10048 27872
rect 9232 27832 10048 27860
rect 10042 27820 10048 27832
rect 10100 27820 10106 27872
rect 10502 27820 10508 27872
rect 10560 27860 10566 27872
rect 12802 27860 12808 27872
rect 10560 27832 12808 27860
rect 10560 27820 10566 27832
rect 12802 27820 12808 27832
rect 12860 27820 12866 27872
rect 13630 27820 13636 27872
rect 13688 27820 13694 27872
rect 14182 27820 14188 27872
rect 14240 27820 14246 27872
rect 1104 27770 14812 27792
rect 1104 27718 2663 27770
rect 2715 27718 2727 27770
rect 2779 27718 2791 27770
rect 2843 27718 2855 27770
rect 2907 27718 2919 27770
rect 2971 27718 6090 27770
rect 6142 27718 6154 27770
rect 6206 27718 6218 27770
rect 6270 27718 6282 27770
rect 6334 27718 6346 27770
rect 6398 27718 9517 27770
rect 9569 27718 9581 27770
rect 9633 27718 9645 27770
rect 9697 27718 9709 27770
rect 9761 27718 9773 27770
rect 9825 27718 12944 27770
rect 12996 27718 13008 27770
rect 13060 27718 13072 27770
rect 13124 27718 13136 27770
rect 13188 27718 13200 27770
rect 13252 27718 14812 27770
rect 1104 27696 14812 27718
rect 11333 27659 11391 27665
rect 11333 27625 11345 27659
rect 11379 27656 11391 27659
rect 11885 27659 11943 27665
rect 11379 27628 11836 27656
rect 11379 27625 11391 27628
rect 11333 27619 11391 27625
rect 11808 27588 11836 27628
rect 11885 27625 11897 27659
rect 11931 27656 11943 27659
rect 13538 27656 13544 27668
rect 11931 27628 13544 27656
rect 11931 27625 11943 27628
rect 11885 27619 11943 27625
rect 13538 27616 13544 27628
rect 13596 27616 13602 27668
rect 11808 27560 14228 27588
rect 11992 27492 12873 27520
rect 5994 27412 6000 27464
rect 6052 27452 6058 27464
rect 6089 27455 6147 27461
rect 6089 27452 6101 27455
rect 6052 27424 6101 27452
rect 6052 27412 6058 27424
rect 6089 27421 6101 27424
rect 6135 27421 6147 27455
rect 6089 27415 6147 27421
rect 6347 27425 6405 27431
rect 6347 27391 6359 27425
rect 6393 27422 6405 27425
rect 6393 27391 6408 27422
rect 8202 27412 8208 27464
rect 8260 27452 8266 27464
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8260 27424 8953 27452
rect 8260 27412 8266 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 9183 27455 9241 27461
rect 9183 27452 9195 27455
rect 8941 27415 8999 27421
rect 9048 27424 9195 27452
rect 6347 27385 6408 27391
rect 6380 27384 6408 27385
rect 9048 27384 9076 27424
rect 9183 27421 9195 27424
rect 9229 27421 9241 27455
rect 9183 27415 9241 27421
rect 10870 27412 10876 27464
rect 10928 27452 10934 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 10928 27424 11529 27452
rect 10928 27412 10934 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11517 27415 11575 27421
rect 11790 27412 11796 27464
rect 11848 27412 11854 27464
rect 6380 27356 6500 27384
rect 6472 27328 6500 27356
rect 8588 27356 9076 27384
rect 8588 27328 8616 27356
rect 9674 27344 9680 27396
rect 9732 27384 9738 27396
rect 11992 27384 12020 27492
rect 12066 27412 12072 27464
rect 12124 27412 12130 27464
rect 12342 27412 12348 27464
rect 12400 27412 12406 27464
rect 12845 27461 12873 27492
rect 12805 27455 12873 27461
rect 12805 27421 12817 27455
rect 12851 27421 12873 27455
rect 12805 27420 12873 27421
rect 12805 27415 12863 27420
rect 13078 27412 13084 27464
rect 13136 27412 13142 27464
rect 13357 27455 13415 27461
rect 13357 27421 13369 27455
rect 13403 27452 13415 27455
rect 13446 27452 13452 27464
rect 13403 27424 13452 27452
rect 13403 27421 13415 27424
rect 13357 27415 13415 27421
rect 13446 27412 13452 27424
rect 13504 27412 13510 27464
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27452 13599 27455
rect 14090 27452 14096 27464
rect 13587 27424 14096 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 14090 27412 14096 27424
rect 14148 27412 14154 27464
rect 14200 27461 14228 27560
rect 14185 27455 14243 27461
rect 14185 27421 14197 27455
rect 14231 27421 14243 27455
rect 14185 27415 14243 27421
rect 13630 27384 13636 27396
rect 9732 27356 12020 27384
rect 12544 27356 13636 27384
rect 9732 27344 9738 27356
rect 6454 27276 6460 27328
rect 6512 27276 6518 27328
rect 7101 27319 7159 27325
rect 7101 27285 7113 27319
rect 7147 27316 7159 27319
rect 7190 27316 7196 27328
rect 7147 27288 7196 27316
rect 7147 27285 7159 27288
rect 7101 27279 7159 27285
rect 7190 27276 7196 27288
rect 7248 27276 7254 27328
rect 8570 27276 8576 27328
rect 8628 27276 8634 27328
rect 9766 27276 9772 27328
rect 9824 27316 9830 27328
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 9824 27288 9965 27316
rect 9824 27276 9830 27288
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 11609 27319 11667 27325
rect 11609 27285 11621 27319
rect 11655 27316 11667 27319
rect 11974 27316 11980 27328
rect 11655 27288 11980 27316
rect 11655 27285 11667 27288
rect 11609 27279 11667 27285
rect 11974 27276 11980 27288
rect 12032 27276 12038 27328
rect 12161 27319 12219 27325
rect 12161 27285 12173 27319
rect 12207 27316 12219 27319
rect 12544 27316 12572 27356
rect 13630 27344 13636 27356
rect 13688 27344 13694 27396
rect 13906 27344 13912 27396
rect 13964 27344 13970 27396
rect 12207 27288 12572 27316
rect 12207 27285 12219 27288
rect 12161 27279 12219 27285
rect 12618 27276 12624 27328
rect 12676 27276 12682 27328
rect 12894 27276 12900 27328
rect 12952 27276 12958 27328
rect 13173 27319 13231 27325
rect 13173 27285 13185 27319
rect 13219 27316 13231 27319
rect 13722 27316 13728 27328
rect 13219 27288 13728 27316
rect 13219 27285 13231 27288
rect 13173 27279 13231 27285
rect 13722 27276 13728 27288
rect 13780 27276 13786 27328
rect 14369 27319 14427 27325
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14415 27288 15056 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 1104 27226 14971 27248
rect 1104 27174 4376 27226
rect 4428 27174 4440 27226
rect 4492 27174 4504 27226
rect 4556 27174 4568 27226
rect 4620 27174 4632 27226
rect 4684 27174 7803 27226
rect 7855 27174 7867 27226
rect 7919 27174 7931 27226
rect 7983 27174 7995 27226
rect 8047 27174 8059 27226
rect 8111 27174 11230 27226
rect 11282 27174 11294 27226
rect 11346 27174 11358 27226
rect 11410 27174 11422 27226
rect 11474 27174 11486 27226
rect 11538 27174 14657 27226
rect 14709 27174 14721 27226
rect 14773 27174 14785 27226
rect 14837 27174 14849 27226
rect 14901 27174 14913 27226
rect 14965 27174 14971 27226
rect 1104 27152 14971 27174
rect 5534 27072 5540 27124
rect 5592 27112 5598 27124
rect 8294 27112 8300 27124
rect 5592 27084 8300 27112
rect 5592 27072 5598 27084
rect 8294 27072 8300 27084
rect 8352 27072 8358 27124
rect 8481 27115 8539 27121
rect 8481 27081 8493 27115
rect 8527 27112 8539 27115
rect 9674 27112 9680 27124
rect 8527 27084 9680 27112
rect 8527 27081 8539 27084
rect 8481 27075 8539 27081
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 10413 27115 10471 27121
rect 10413 27081 10425 27115
rect 10459 27112 10471 27115
rect 11054 27112 11060 27124
rect 10459 27084 11060 27112
rect 10459 27081 10471 27084
rect 10413 27075 10471 27081
rect 11054 27072 11060 27084
rect 11112 27072 11118 27124
rect 11974 27072 11980 27124
rect 12032 27072 12038 27124
rect 12069 27115 12127 27121
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12342 27112 12348 27124
rect 12115 27084 12348 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12342 27072 12348 27084
rect 12400 27072 12406 27124
rect 12618 27072 12624 27124
rect 12676 27072 12682 27124
rect 12894 27072 12900 27124
rect 12952 27112 12958 27124
rect 12952 27084 13032 27112
rect 12952 27072 12958 27084
rect 8312 27044 8340 27072
rect 11992 27044 12020 27072
rect 12437 27047 12495 27053
rect 8312 27016 8432 27044
rect 11992 27016 12388 27044
rect 750 26936 756 26988
rect 808 26976 814 26988
rect 1489 26979 1547 26985
rect 1489 26976 1501 26979
rect 808 26948 1501 26976
rect 808 26936 814 26948
rect 1489 26945 1501 26948
rect 1535 26945 1547 26979
rect 1489 26939 1547 26945
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 6788 26948 6837 26976
rect 6788 26936 6794 26948
rect 6825 26945 6837 26948
rect 6871 26945 6883 26979
rect 8404 26976 8432 27016
rect 8404 26948 8892 26976
rect 6825 26939 6883 26945
rect 6641 26911 6699 26917
rect 6641 26877 6653 26911
rect 6687 26877 6699 26911
rect 6641 26871 6699 26877
rect 1581 26775 1639 26781
rect 1581 26741 1593 26775
rect 1627 26772 1639 26775
rect 1854 26772 1860 26784
rect 1627 26744 1860 26772
rect 1627 26741 1639 26744
rect 1581 26735 1639 26741
rect 1854 26732 1860 26744
rect 1912 26732 1918 26784
rect 6656 26772 6684 26871
rect 7190 26868 7196 26920
rect 7248 26908 7254 26920
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 7248 26880 7297 26908
rect 7248 26868 7254 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 7558 26868 7564 26920
rect 7616 26868 7622 26920
rect 7742 26917 7748 26920
rect 7699 26911 7748 26917
rect 7699 26877 7711 26911
rect 7745 26877 7748 26911
rect 7699 26871 7748 26877
rect 7742 26868 7748 26871
rect 7800 26868 7806 26920
rect 7834 26868 7840 26920
rect 7892 26868 7898 26920
rect 8573 26911 8631 26917
rect 8573 26877 8585 26911
rect 8619 26877 8631 26911
rect 8573 26871 8631 26877
rect 8588 26840 8616 26871
rect 8754 26868 8760 26920
rect 8812 26868 8818 26920
rect 8864 26908 8892 26948
rect 9766 26936 9772 26988
rect 9824 26936 9830 26988
rect 11977 26979 12035 26985
rect 11977 26945 11989 26979
rect 12023 26945 12035 26979
rect 11977 26939 12035 26945
rect 8864 26880 9168 26908
rect 9030 26840 9036 26852
rect 8588 26812 9036 26840
rect 9030 26800 9036 26812
rect 9088 26800 9094 26852
rect 9140 26840 9168 26880
rect 9214 26868 9220 26920
rect 9272 26868 9278 26920
rect 9493 26911 9551 26917
rect 9493 26908 9505 26911
rect 9306 26880 9505 26908
rect 9306 26840 9334 26880
rect 9493 26877 9505 26880
rect 9539 26877 9551 26911
rect 9493 26871 9551 26877
rect 9582 26868 9588 26920
rect 9640 26917 9646 26920
rect 9640 26911 9668 26917
rect 9656 26877 9668 26911
rect 11992 26908 12020 26939
rect 12158 26936 12164 26988
rect 12216 26976 12222 26988
rect 12253 26979 12311 26985
rect 12253 26976 12265 26979
rect 12216 26948 12265 26976
rect 12216 26936 12222 26948
rect 12253 26945 12265 26948
rect 12299 26945 12311 26979
rect 12360 26976 12388 27016
rect 12437 27013 12449 27047
rect 12483 27044 12495 27047
rect 12636 27044 12664 27072
rect 13004 27053 13032 27084
rect 13078 27072 13084 27124
rect 13136 27072 13142 27124
rect 14918 27072 14924 27124
rect 14976 27112 14982 27124
rect 15028 27112 15056 27288
rect 14976 27084 15056 27112
rect 14976 27072 14982 27084
rect 12483 27016 12664 27044
rect 12989 27047 13047 27053
rect 12483 27013 12495 27016
rect 12437 27007 12495 27013
rect 12989 27013 13001 27047
rect 13035 27013 13047 27047
rect 12989 27007 13047 27013
rect 13096 26976 13124 27072
rect 13446 27004 13452 27056
rect 13504 27044 13510 27056
rect 14458 27044 14464 27056
rect 13504 27016 14464 27044
rect 13504 27004 13510 27016
rect 14458 27004 14464 27016
rect 14516 27004 14522 27056
rect 13541 26979 13599 26985
rect 13541 26976 13553 26979
rect 12360 26948 12664 26976
rect 13096 26948 13553 26976
rect 12253 26939 12311 26945
rect 12342 26908 12348 26920
rect 11992 26880 12348 26908
rect 9640 26871 9668 26877
rect 9640 26868 9646 26871
rect 12342 26868 12348 26880
rect 12400 26868 12406 26920
rect 12636 26908 12664 26948
rect 13541 26945 13553 26948
rect 13587 26945 13599 26979
rect 13541 26939 13599 26945
rect 13998 26936 14004 26988
rect 14056 26936 14062 26988
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26945 14151 26979
rect 14093 26939 14151 26945
rect 14016 26908 14044 26936
rect 12636 26880 14044 26908
rect 9140 26812 9334 26840
rect 11793 26843 11851 26849
rect 11793 26809 11805 26843
rect 11839 26840 11851 26843
rect 14108 26840 14136 26939
rect 11839 26812 14136 26840
rect 11839 26809 11851 26812
rect 11793 26803 11851 26809
rect 6822 26772 6828 26784
rect 6656 26744 6828 26772
rect 6822 26732 6828 26744
rect 6880 26772 6886 26784
rect 7650 26772 7656 26784
rect 6880 26744 7656 26772
rect 6880 26732 6886 26744
rect 7650 26732 7656 26744
rect 7708 26732 7714 26784
rect 7742 26732 7748 26784
rect 7800 26772 7806 26784
rect 8938 26772 8944 26784
rect 7800 26744 8944 26772
rect 7800 26732 7806 26744
rect 8938 26732 8944 26744
rect 8996 26772 9002 26784
rect 9582 26772 9588 26784
rect 8996 26744 9588 26772
rect 8996 26732 9002 26744
rect 9582 26732 9588 26744
rect 9640 26732 9646 26784
rect 12342 26732 12348 26784
rect 12400 26772 12406 26784
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 12400 26744 12541 26772
rect 12400 26732 12406 26744
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 12529 26735 12587 26741
rect 13262 26732 13268 26784
rect 13320 26732 13326 26784
rect 13814 26732 13820 26784
rect 13872 26732 13878 26784
rect 14369 26775 14427 26781
rect 14369 26741 14381 26775
rect 14415 26772 14427 26775
rect 15286 26772 15292 26784
rect 14415 26744 15292 26772
rect 14415 26741 14427 26744
rect 14369 26735 14427 26741
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 1104 26682 14812 26704
rect 1104 26630 2663 26682
rect 2715 26630 2727 26682
rect 2779 26630 2791 26682
rect 2843 26630 2855 26682
rect 2907 26630 2919 26682
rect 2971 26630 6090 26682
rect 6142 26630 6154 26682
rect 6206 26630 6218 26682
rect 6270 26630 6282 26682
rect 6334 26630 6346 26682
rect 6398 26630 9517 26682
rect 9569 26630 9581 26682
rect 9633 26630 9645 26682
rect 9697 26630 9709 26682
rect 9761 26630 9773 26682
rect 9825 26630 12944 26682
rect 12996 26630 13008 26682
rect 13060 26630 13072 26682
rect 13124 26630 13136 26682
rect 13188 26630 13200 26682
rect 13252 26630 14812 26682
rect 1104 26608 14812 26630
rect 7469 26571 7527 26577
rect 7469 26537 7481 26571
rect 7515 26568 7527 26571
rect 7834 26568 7840 26580
rect 7515 26540 7840 26568
rect 7515 26537 7527 26540
rect 7469 26531 7527 26537
rect 7834 26528 7840 26540
rect 7892 26528 7898 26580
rect 9950 26528 9956 26580
rect 10008 26568 10014 26580
rect 11698 26568 11704 26580
rect 10008 26540 11704 26568
rect 10008 26528 10014 26540
rect 7558 26460 7564 26512
rect 7616 26500 7622 26512
rect 8846 26500 8852 26512
rect 7616 26472 8852 26500
rect 7616 26460 7622 26472
rect 8846 26460 8852 26472
rect 8904 26460 8910 26512
rect 9966 26500 9994 26528
rect 9876 26472 9994 26500
rect 10873 26503 10931 26509
rect 9876 26441 9904 26472
rect 10873 26469 10885 26503
rect 10919 26500 10931 26503
rect 11146 26500 11152 26512
rect 10919 26472 11152 26500
rect 10919 26469 10931 26472
rect 10873 26463 10931 26469
rect 11146 26460 11152 26472
rect 11204 26460 11210 26512
rect 11256 26441 11284 26540
rect 11698 26528 11704 26540
rect 11756 26568 11762 26580
rect 11756 26540 12664 26568
rect 11756 26528 11762 26540
rect 12636 26441 12664 26540
rect 13722 26528 13728 26580
rect 13780 26528 13786 26580
rect 9861 26435 9919 26441
rect 9861 26401 9873 26435
rect 9907 26401 9919 26435
rect 9861 26395 9919 26401
rect 11241 26435 11299 26441
rect 11241 26401 11253 26435
rect 11287 26401 11299 26435
rect 11241 26395 11299 26401
rect 12621 26435 12679 26441
rect 12621 26401 12633 26435
rect 12667 26401 12679 26435
rect 12621 26395 12679 26401
rect 1854 26324 1860 26376
rect 1912 26364 1918 26376
rect 5442 26364 5448 26376
rect 1912 26336 5448 26364
rect 1912 26324 1918 26336
rect 5442 26324 5448 26336
rect 5500 26324 5506 26376
rect 5994 26324 6000 26376
rect 6052 26364 6058 26376
rect 6362 26364 6368 26376
rect 6052 26336 6368 26364
rect 6052 26324 6058 26336
rect 6362 26324 6368 26336
rect 6420 26364 6426 26376
rect 6730 26373 6736 26376
rect 6457 26367 6515 26373
rect 6457 26364 6469 26367
rect 6420 26336 6469 26364
rect 6420 26324 6426 26336
rect 6457 26333 6469 26336
rect 6503 26333 6515 26367
rect 6699 26367 6736 26373
rect 6699 26364 6711 26367
rect 6457 26327 6515 26333
rect 6556 26336 6711 26364
rect 1486 26256 1492 26308
rect 1544 26256 1550 26308
rect 1673 26299 1731 26305
rect 1673 26265 1685 26299
rect 1719 26296 1731 26299
rect 6556 26296 6584 26336
rect 6699 26333 6711 26336
rect 6699 26327 6736 26333
rect 6730 26324 6736 26327
rect 6788 26324 6794 26376
rect 10042 26324 10048 26376
rect 10100 26364 10106 26376
rect 10135 26367 10193 26373
rect 10135 26364 10147 26367
rect 10100 26336 10147 26364
rect 10100 26324 10106 26336
rect 10135 26333 10147 26336
rect 10181 26333 10193 26367
rect 11499 26367 11557 26373
rect 11499 26364 11511 26367
rect 10135 26327 10193 26333
rect 10980 26336 11511 26364
rect 1719 26268 6584 26296
rect 1719 26265 1731 26268
rect 1673 26259 1731 26265
rect 7558 26256 7564 26308
rect 7616 26296 7622 26308
rect 8570 26296 8576 26308
rect 7616 26268 8576 26296
rect 7616 26256 7622 26268
rect 8570 26256 8576 26268
rect 8628 26296 8634 26308
rect 10980 26296 11008 26336
rect 11499 26333 11511 26336
rect 11545 26333 11557 26367
rect 11499 26327 11557 26333
rect 12863 26367 12921 26373
rect 12863 26333 12875 26367
rect 12909 26364 12921 26367
rect 13538 26364 13544 26376
rect 12909 26336 13544 26364
rect 12909 26333 12921 26336
rect 12863 26327 12921 26333
rect 13538 26324 13544 26336
rect 13596 26324 13602 26376
rect 13740 26364 13768 26528
rect 14185 26367 14243 26373
rect 14185 26364 14197 26367
rect 13740 26336 14197 26364
rect 14185 26333 14197 26336
rect 14231 26333 14243 26367
rect 14185 26327 14243 26333
rect 8628 26268 11008 26296
rect 8628 26256 8634 26268
rect 10980 26240 11008 26268
rect 4062 26188 4068 26240
rect 4120 26228 4126 26240
rect 8478 26228 8484 26240
rect 4120 26200 8484 26228
rect 4120 26188 4126 26200
rect 8478 26188 8484 26200
rect 8536 26188 8542 26240
rect 10962 26188 10968 26240
rect 11020 26188 11026 26240
rect 12253 26231 12311 26237
rect 12253 26197 12265 26231
rect 12299 26228 12311 26231
rect 12710 26228 12716 26240
rect 12299 26200 12716 26228
rect 12299 26197 12311 26200
rect 12253 26191 12311 26197
rect 12710 26188 12716 26200
rect 12768 26188 12774 26240
rect 13630 26188 13636 26240
rect 13688 26188 13694 26240
rect 14366 26188 14372 26240
rect 14424 26188 14430 26240
rect 1104 26138 14971 26160
rect 1104 26086 4376 26138
rect 4428 26086 4440 26138
rect 4492 26086 4504 26138
rect 4556 26086 4568 26138
rect 4620 26086 4632 26138
rect 4684 26086 7803 26138
rect 7855 26086 7867 26138
rect 7919 26086 7931 26138
rect 7983 26086 7995 26138
rect 8047 26086 8059 26138
rect 8111 26086 11230 26138
rect 11282 26086 11294 26138
rect 11346 26086 11358 26138
rect 11410 26086 11422 26138
rect 11474 26086 11486 26138
rect 11538 26086 14657 26138
rect 14709 26086 14721 26138
rect 14773 26086 14785 26138
rect 14837 26086 14849 26138
rect 14901 26086 14913 26138
rect 14965 26086 14971 26138
rect 1104 26064 14971 26086
rect 6638 25984 6644 26036
rect 6696 25984 6702 26036
rect 8202 26024 8208 26036
rect 8036 25996 8208 26024
rect 6656 25927 6684 25984
rect 6623 25921 6684 25927
rect 6623 25887 6635 25921
rect 6669 25890 6684 25921
rect 6669 25887 6681 25890
rect 6623 25881 6681 25887
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 8036 25897 8064 25996
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 9950 25984 9956 26036
rect 10008 25984 10014 26036
rect 12434 25984 12440 26036
rect 12492 26024 12498 26036
rect 13357 26027 13415 26033
rect 13357 26024 13369 26027
rect 12492 25996 13369 26024
rect 12492 25984 12498 25996
rect 13357 25993 13369 25996
rect 13403 25993 13415 26027
rect 13357 25987 13415 25993
rect 9858 25956 9864 25968
rect 9646 25928 9864 25956
rect 8021 25891 8079 25897
rect 8021 25888 8033 25891
rect 7248 25860 8033 25888
rect 7248 25848 7254 25860
rect 8021 25857 8033 25860
rect 8067 25857 8079 25891
rect 8294 25888 8300 25900
rect 8255 25860 8300 25888
rect 8021 25851 8079 25857
rect 8294 25848 8300 25860
rect 8352 25888 8358 25900
rect 9646 25888 9674 25928
rect 9858 25916 9864 25928
rect 9916 25916 9922 25968
rect 8352 25860 9674 25888
rect 9968 25888 9996 25984
rect 10134 25916 10140 25968
rect 10192 25956 10198 25968
rect 10192 25928 10272 25956
rect 10192 25916 10198 25928
rect 10244 25918 10272 25928
rect 10303 25921 10361 25927
rect 10303 25918 10315 25921
rect 10045 25891 10103 25897
rect 10045 25888 10057 25891
rect 9968 25860 10057 25888
rect 8352 25848 8358 25860
rect 10045 25857 10057 25860
rect 10091 25857 10103 25891
rect 10244 25890 10315 25918
rect 10303 25887 10315 25890
rect 10349 25887 10361 25921
rect 11698 25916 11704 25968
rect 11756 25916 11762 25968
rect 13446 25916 13452 25968
rect 13504 25956 13510 25968
rect 14093 25959 14151 25965
rect 14093 25956 14105 25959
rect 13504 25928 14105 25956
rect 13504 25916 13510 25928
rect 14093 25925 14105 25928
rect 14139 25925 14151 25959
rect 14093 25919 14151 25925
rect 10303 25881 10361 25887
rect 10045 25851 10103 25857
rect 10686 25848 10692 25900
rect 10744 25888 10750 25900
rect 11517 25891 11575 25897
rect 10744 25860 11284 25888
rect 10744 25848 10750 25860
rect 6362 25780 6368 25832
rect 6420 25780 6426 25832
rect 11146 25780 11152 25832
rect 11204 25780 11210 25832
rect 11256 25820 11284 25860
rect 11517 25857 11529 25891
rect 11563 25888 11575 25891
rect 11716 25888 11744 25916
rect 11563 25860 11744 25888
rect 11563 25857 11575 25860
rect 11517 25851 11575 25857
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 13354 25848 13360 25900
rect 13412 25888 13418 25900
rect 13541 25891 13599 25897
rect 13541 25888 13553 25891
rect 13412 25860 13553 25888
rect 13412 25848 13418 25860
rect 13541 25857 13553 25860
rect 13587 25857 13599 25891
rect 13541 25851 13599 25857
rect 11701 25823 11759 25829
rect 11701 25820 11713 25823
rect 11256 25792 11713 25820
rect 11701 25789 11713 25792
rect 11747 25789 11759 25823
rect 11701 25783 11759 25789
rect 12434 25780 12440 25832
rect 12492 25780 12498 25832
rect 12526 25780 12532 25832
rect 12584 25829 12590 25832
rect 12584 25823 12612 25829
rect 12600 25789 12612 25823
rect 12584 25783 12612 25789
rect 12584 25780 12590 25783
rect 15102 25780 15108 25832
rect 15160 25820 15166 25832
rect 15160 25792 15332 25820
rect 15160 25780 15166 25792
rect 6380 25684 6408 25780
rect 11164 25752 11192 25780
rect 12161 25755 12219 25761
rect 12161 25752 12173 25755
rect 11164 25724 12173 25752
rect 12161 25721 12173 25724
rect 12207 25721 12219 25755
rect 12161 25715 12219 25721
rect 6638 25684 6644 25696
rect 6380 25656 6644 25684
rect 6638 25644 6644 25656
rect 6696 25644 6702 25696
rect 7374 25644 7380 25696
rect 7432 25644 7438 25696
rect 9033 25687 9091 25693
rect 9033 25653 9045 25687
rect 9079 25684 9091 25687
rect 9214 25684 9220 25696
rect 9079 25656 9220 25684
rect 9079 25653 9091 25656
rect 9033 25647 9091 25653
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 11054 25644 11060 25696
rect 11112 25644 11118 25696
rect 11974 25644 11980 25696
rect 12032 25684 12038 25696
rect 12526 25684 12532 25696
rect 12032 25656 12532 25684
rect 12032 25644 12038 25656
rect 12526 25644 12532 25656
rect 12584 25644 12590 25696
rect 13814 25644 13820 25696
rect 13872 25644 13878 25696
rect 14369 25687 14427 25693
rect 14369 25653 14381 25687
rect 14415 25684 14427 25687
rect 15102 25684 15108 25696
rect 14415 25656 15108 25684
rect 14415 25653 14427 25656
rect 14369 25647 14427 25653
rect 15102 25644 15108 25656
rect 15160 25644 15166 25696
rect 1104 25594 14812 25616
rect 1104 25542 2663 25594
rect 2715 25542 2727 25594
rect 2779 25542 2791 25594
rect 2843 25542 2855 25594
rect 2907 25542 2919 25594
rect 2971 25542 6090 25594
rect 6142 25542 6154 25594
rect 6206 25542 6218 25594
rect 6270 25542 6282 25594
rect 6334 25542 6346 25594
rect 6398 25542 9517 25594
rect 9569 25542 9581 25594
rect 9633 25542 9645 25594
rect 9697 25542 9709 25594
rect 9761 25542 9773 25594
rect 9825 25542 12944 25594
rect 12996 25542 13008 25594
rect 13060 25542 13072 25594
rect 13124 25542 13136 25594
rect 13188 25542 13200 25594
rect 13252 25542 14812 25594
rect 15304 25560 15332 25792
rect 1104 25520 14812 25542
rect 15286 25508 15292 25560
rect 15344 25508 15350 25560
rect 6362 25480 6368 25492
rect 1688 25452 6368 25480
rect 1688 25353 1716 25452
rect 6362 25440 6368 25452
rect 6420 25440 6426 25492
rect 7374 25440 7380 25492
rect 7432 25440 7438 25492
rect 7469 25483 7527 25489
rect 7469 25449 7481 25483
rect 7515 25480 7527 25483
rect 9950 25480 9956 25492
rect 7515 25452 9956 25480
rect 7515 25449 7527 25452
rect 7469 25443 7527 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 11054 25440 11060 25492
rect 11112 25440 11118 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 12802 25480 12808 25492
rect 12492 25452 12808 25480
rect 12492 25440 12498 25452
rect 12802 25440 12808 25452
rect 12860 25440 12866 25492
rect 5261 25415 5319 25421
rect 5261 25381 5273 25415
rect 5307 25412 5319 25415
rect 6273 25415 6331 25421
rect 6273 25412 6285 25415
rect 5307 25384 6285 25412
rect 5307 25381 5319 25384
rect 5261 25375 5319 25381
rect 6273 25381 6285 25384
rect 6319 25381 6331 25415
rect 6273 25375 6331 25381
rect 1673 25347 1731 25353
rect 1673 25313 1685 25347
rect 1719 25313 1731 25347
rect 1673 25307 1731 25313
rect 6825 25347 6883 25353
rect 6825 25313 6837 25347
rect 6871 25344 6883 25347
rect 7392 25344 7420 25440
rect 11072 25412 11100 25440
rect 12529 25415 12587 25421
rect 12529 25412 12541 25415
rect 11072 25384 12541 25412
rect 12529 25381 12541 25384
rect 12575 25381 12587 25415
rect 12529 25375 12587 25381
rect 12069 25347 12127 25353
rect 12069 25344 12081 25347
rect 6871 25316 7420 25344
rect 11716 25316 12081 25344
rect 6871 25313 6883 25316
rect 6825 25307 6883 25313
rect 11716 25288 11744 25316
rect 12069 25313 12081 25316
rect 12115 25313 12127 25347
rect 12805 25347 12863 25353
rect 12805 25344 12817 25347
rect 12069 25307 12127 25313
rect 12268 25316 12817 25344
rect 750 25236 756 25288
rect 808 25276 814 25288
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 808 25248 1409 25276
rect 808 25236 814 25248
rect 1397 25245 1409 25248
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4249 25239 4307 25245
rect 4523 25279 4581 25285
rect 4523 25245 4535 25279
rect 4569 25276 4581 25279
rect 5442 25276 5448 25288
rect 4569 25248 5448 25276
rect 4569 25245 4581 25248
rect 4523 25239 4581 25245
rect 4264 25140 4292 25239
rect 5442 25236 5448 25248
rect 5500 25236 5506 25288
rect 5629 25279 5687 25285
rect 5629 25245 5641 25279
rect 5675 25276 5687 25279
rect 5718 25276 5724 25288
rect 5675 25248 5724 25276
rect 5675 25245 5687 25248
rect 5629 25239 5687 25245
rect 5718 25236 5724 25248
rect 5776 25236 5782 25288
rect 5810 25236 5816 25288
rect 5868 25236 5874 25288
rect 6546 25236 6552 25288
rect 6604 25236 6610 25288
rect 6730 25285 6736 25288
rect 6687 25279 6736 25285
rect 6687 25245 6699 25279
rect 6733 25245 6736 25279
rect 6687 25239 6736 25245
rect 6730 25236 6736 25239
rect 6788 25236 6794 25288
rect 9950 25236 9956 25288
rect 10008 25236 10014 25288
rect 10502 25236 10508 25288
rect 10560 25276 10566 25288
rect 10962 25276 10968 25288
rect 10560 25248 10968 25276
rect 10560 25236 10566 25248
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 11698 25236 11704 25288
rect 11756 25236 11762 25288
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25276 11943 25279
rect 11974 25276 11980 25288
rect 11931 25248 11980 25276
rect 11931 25245 11943 25248
rect 11885 25239 11943 25245
rect 11974 25236 11980 25248
rect 12032 25236 12038 25288
rect 12268 25276 12296 25316
rect 12805 25313 12817 25316
rect 12851 25313 12863 25347
rect 12805 25307 12863 25313
rect 13081 25347 13139 25353
rect 13081 25313 13093 25347
rect 13127 25344 13139 25347
rect 13630 25344 13636 25356
rect 13127 25316 13636 25344
rect 13127 25313 13139 25316
rect 13081 25307 13139 25313
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 12084 25248 12296 25276
rect 7374 25168 7380 25220
rect 7432 25208 7438 25220
rect 8662 25208 8668 25220
rect 7432 25180 8668 25208
rect 7432 25168 7438 25180
rect 8662 25168 8668 25180
rect 8720 25168 8726 25220
rect 9968 25208 9996 25236
rect 12084 25208 12112 25248
rect 12894 25236 12900 25288
rect 12952 25285 12958 25288
rect 12952 25279 12980 25285
rect 12968 25245 12980 25279
rect 12952 25239 12980 25245
rect 12952 25236 12958 25239
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 14185 25279 14243 25285
rect 14185 25276 14197 25279
rect 13780 25248 14197 25276
rect 13780 25236 13786 25248
rect 14185 25245 14197 25248
rect 14231 25245 14243 25279
rect 14185 25239 14243 25245
rect 9968 25180 12112 25208
rect 13814 25168 13820 25220
rect 13872 25208 13878 25220
rect 15562 25208 15568 25220
rect 13872 25180 15568 25208
rect 13872 25168 13878 25180
rect 15562 25168 15568 25180
rect 15620 25168 15626 25220
rect 6638 25140 6644 25152
rect 4264 25112 6644 25140
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 10686 25140 10692 25152
rect 6788 25112 10692 25140
rect 6788 25100 6794 25112
rect 10686 25100 10692 25112
rect 10744 25100 10750 25152
rect 10870 25100 10876 25152
rect 10928 25140 10934 25152
rect 13725 25143 13783 25149
rect 13725 25140 13737 25143
rect 10928 25112 13737 25140
rect 10928 25100 10934 25112
rect 13725 25109 13737 25112
rect 13771 25109 13783 25143
rect 13725 25103 13783 25109
rect 14366 25100 14372 25152
rect 14424 25100 14430 25152
rect 1104 25050 14971 25072
rect 1104 24998 4376 25050
rect 4428 24998 4440 25050
rect 4492 24998 4504 25050
rect 4556 24998 4568 25050
rect 4620 24998 4632 25050
rect 4684 24998 7803 25050
rect 7855 24998 7867 25050
rect 7919 24998 7931 25050
rect 7983 24998 7995 25050
rect 8047 24998 8059 25050
rect 8111 24998 11230 25050
rect 11282 24998 11294 25050
rect 11346 24998 11358 25050
rect 11410 24998 11422 25050
rect 11474 24998 11486 25050
rect 11538 24998 14657 25050
rect 14709 24998 14721 25050
rect 14773 24998 14785 25050
rect 14837 24998 14849 25050
rect 14901 24998 14913 25050
rect 14965 24998 14971 25050
rect 1104 24976 14971 24998
rect 10134 24896 10140 24948
rect 10192 24896 10198 24948
rect 12268 24908 12848 24936
rect 1673 24871 1731 24877
rect 1673 24837 1685 24871
rect 1719 24868 1731 24871
rect 7558 24868 7564 24880
rect 1719 24840 7564 24868
rect 1719 24837 1731 24840
rect 1673 24831 1731 24837
rect 7558 24828 7564 24840
rect 7616 24828 7622 24880
rect 750 24760 756 24812
rect 808 24800 814 24812
rect 1489 24803 1547 24809
rect 1489 24800 1501 24803
rect 808 24772 1501 24800
rect 808 24760 814 24772
rect 1489 24769 1501 24772
rect 1535 24769 1547 24803
rect 1489 24763 1547 24769
rect 6915 24803 6973 24809
rect 6915 24769 6927 24803
rect 6961 24800 6973 24803
rect 7374 24800 7380 24812
rect 6961 24772 7380 24800
rect 6961 24769 6973 24772
rect 6915 24763 6973 24769
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24800 8079 24803
rect 8067 24772 8432 24800
rect 8067 24769 8079 24772
rect 8021 24763 8079 24769
rect 5994 24692 6000 24744
rect 6052 24732 6058 24744
rect 6641 24735 6699 24741
rect 6641 24732 6653 24735
rect 6052 24704 6653 24732
rect 6052 24692 6058 24704
rect 6641 24701 6653 24704
rect 6687 24701 6699 24735
rect 6641 24695 6699 24701
rect 7558 24692 7564 24744
rect 7616 24732 7622 24744
rect 8205 24735 8263 24741
rect 8205 24732 8217 24735
rect 7616 24704 8217 24732
rect 7616 24692 7622 24704
rect 8205 24701 8217 24704
rect 8251 24701 8263 24735
rect 8404 24732 8432 24772
rect 9214 24760 9220 24812
rect 9272 24760 9278 24812
rect 10134 24800 10162 24896
rect 12268 24868 12296 24908
rect 11992 24840 12296 24868
rect 10195 24803 10253 24809
rect 10195 24800 10207 24803
rect 10134 24772 10207 24800
rect 10195 24769 10207 24772
rect 10241 24769 10253 24803
rect 11992 24800 12020 24840
rect 10195 24763 10253 24769
rect 11624 24772 12020 24800
rect 8570 24732 8576 24744
rect 8404 24704 8576 24732
rect 8205 24695 8263 24701
rect 8570 24692 8576 24704
rect 8628 24692 8634 24744
rect 9122 24741 9128 24744
rect 8941 24735 8999 24741
rect 8941 24732 8953 24735
rect 8772 24704 8953 24732
rect 8772 24676 8800 24704
rect 8941 24701 8953 24704
rect 8987 24701 8999 24735
rect 8941 24695 8999 24701
rect 9079 24735 9128 24741
rect 9079 24701 9091 24735
rect 9125 24701 9128 24735
rect 9079 24695 9128 24701
rect 9122 24692 9128 24695
rect 9180 24692 9186 24744
rect 9398 24692 9404 24744
rect 9456 24732 9462 24744
rect 9766 24732 9772 24744
rect 9456 24704 9772 24732
rect 9456 24692 9462 24704
rect 9766 24692 9772 24704
rect 9824 24692 9830 24744
rect 9953 24735 10011 24741
rect 9953 24701 9965 24735
rect 9999 24701 10011 24735
rect 9953 24695 10011 24701
rect 7653 24667 7711 24673
rect 7653 24633 7665 24667
rect 7699 24664 7711 24667
rect 8665 24667 8723 24673
rect 8665 24664 8677 24667
rect 7699 24636 8677 24664
rect 7699 24633 7711 24636
rect 7653 24627 7711 24633
rect 8665 24633 8677 24636
rect 8711 24633 8723 24667
rect 8665 24627 8723 24633
rect 8754 24624 8760 24676
rect 8812 24624 8818 24676
rect 9968 24664 9996 24695
rect 11624 24664 11652 24772
rect 12066 24760 12072 24812
rect 12124 24760 12130 24812
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 12820 24800 12848 24908
rect 13648 24840 14044 24868
rect 13648 24800 13676 24840
rect 12492 24772 12781 24800
rect 12820 24772 13676 24800
rect 12492 24760 12498 24772
rect 12161 24735 12219 24741
rect 12161 24701 12173 24735
rect 12207 24701 12219 24735
rect 12753 24732 12781 24772
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 13909 24803 13967 24809
rect 13909 24769 13921 24803
rect 13955 24769 13967 24803
rect 14016 24800 14044 24840
rect 15654 24800 15660 24812
rect 14016 24772 15660 24800
rect 13909 24763 13967 24769
rect 12753 24704 13492 24732
rect 12161 24695 12219 24701
rect 12176 24664 12204 24695
rect 9646 24636 9996 24664
rect 10796 24636 11652 24664
rect 11716 24636 12204 24664
rect 13004 24636 13400 24664
rect 8478 24556 8484 24608
rect 8536 24596 8542 24608
rect 9122 24596 9128 24608
rect 8536 24568 9128 24596
rect 8536 24556 8542 24568
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 9214 24556 9220 24608
rect 9272 24596 9278 24608
rect 9646 24596 9674 24636
rect 9272 24568 9674 24596
rect 9861 24599 9919 24605
rect 9272 24556 9278 24568
rect 9861 24565 9873 24599
rect 9907 24596 9919 24599
rect 10796 24596 10824 24636
rect 9907 24568 10824 24596
rect 9907 24565 9919 24568
rect 9861 24559 9919 24565
rect 10870 24556 10876 24608
rect 10928 24596 10934 24608
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 10928 24568 10977 24596
rect 10928 24556 10934 24568
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 11146 24556 11152 24608
rect 11204 24596 11210 24608
rect 11514 24596 11520 24608
rect 11204 24568 11520 24596
rect 11204 24556 11210 24568
rect 11514 24556 11520 24568
rect 11572 24596 11578 24608
rect 11716 24596 11744 24636
rect 11572 24568 11744 24596
rect 11885 24599 11943 24605
rect 11572 24556 11578 24568
rect 11885 24565 11897 24599
rect 11931 24596 11943 24599
rect 13004 24596 13032 24636
rect 13372 24608 13400 24636
rect 11931 24568 13032 24596
rect 13173 24599 13231 24605
rect 11931 24565 11943 24568
rect 11885 24559 11943 24565
rect 13173 24565 13185 24599
rect 13219 24596 13231 24599
rect 13262 24596 13268 24608
rect 13219 24568 13268 24596
rect 13219 24565 13231 24568
rect 13173 24559 13231 24565
rect 13262 24556 13268 24568
rect 13320 24556 13326 24608
rect 13354 24556 13360 24608
rect 13412 24556 13418 24608
rect 13464 24596 13492 24704
rect 13541 24667 13599 24673
rect 13541 24633 13553 24667
rect 13587 24664 13599 24667
rect 13924 24664 13952 24763
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 14274 24732 14280 24744
rect 13587 24636 13952 24664
rect 14016 24704 14280 24732
rect 13587 24633 13599 24636
rect 13541 24627 13599 24633
rect 14016 24596 14044 24704
rect 14274 24692 14280 24704
rect 14332 24692 14338 24744
rect 13464 24568 14044 24596
rect 14182 24556 14188 24608
rect 14240 24556 14246 24608
rect 1104 24506 14812 24528
rect 1104 24454 2663 24506
rect 2715 24454 2727 24506
rect 2779 24454 2791 24506
rect 2843 24454 2855 24506
rect 2907 24454 2919 24506
rect 2971 24454 6090 24506
rect 6142 24454 6154 24506
rect 6206 24454 6218 24506
rect 6270 24454 6282 24506
rect 6334 24454 6346 24506
rect 6398 24454 9517 24506
rect 9569 24454 9581 24506
rect 9633 24454 9645 24506
rect 9697 24454 9709 24506
rect 9761 24454 9773 24506
rect 9825 24454 12944 24506
rect 12996 24454 13008 24506
rect 13060 24454 13072 24506
rect 13124 24454 13136 24506
rect 13188 24454 13200 24506
rect 13252 24454 14812 24506
rect 1104 24432 14812 24454
rect 5994 24352 6000 24404
rect 6052 24392 6058 24404
rect 7190 24392 7196 24404
rect 6052 24364 7196 24392
rect 6052 24352 6058 24364
rect 7190 24352 7196 24364
rect 7248 24352 7254 24404
rect 9950 24392 9956 24404
rect 8772 24364 9956 24392
rect 8772 24336 8800 24364
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 10134 24352 10140 24404
rect 10192 24352 10198 24404
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 11517 24395 11575 24401
rect 10468 24364 11376 24392
rect 10468 24352 10474 24364
rect 8754 24284 8760 24336
rect 8812 24284 8818 24336
rect 9214 24284 9220 24336
rect 9272 24324 9278 24336
rect 9766 24324 9772 24336
rect 9272 24296 9772 24324
rect 9272 24284 9278 24296
rect 9766 24284 9772 24296
rect 9824 24284 9830 24336
rect 6362 24216 6368 24268
rect 6420 24256 6426 24268
rect 6638 24256 6644 24268
rect 6420 24228 6644 24256
rect 6420 24216 6426 24228
rect 6638 24216 6644 24228
rect 6696 24216 6702 24268
rect 6914 24216 6920 24268
rect 6972 24256 6978 24268
rect 7098 24256 7104 24268
rect 6972 24228 7104 24256
rect 6972 24216 6978 24228
rect 7098 24216 7104 24228
rect 7156 24256 7162 24268
rect 7469 24259 7527 24265
rect 7469 24256 7481 24259
rect 7156 24228 7481 24256
rect 7156 24216 7162 24228
rect 7469 24225 7481 24228
rect 7515 24225 7527 24259
rect 10152 24256 10180 24352
rect 7469 24219 7527 24225
rect 8128 24228 10180 24256
rect 6822 24148 6828 24200
rect 6880 24188 6886 24200
rect 7711 24191 7769 24197
rect 7711 24188 7723 24191
rect 6880 24160 7723 24188
rect 6880 24148 6886 24160
rect 7711 24157 7723 24160
rect 7757 24188 7769 24191
rect 8128 24188 8156 24228
rect 10318 24216 10324 24268
rect 10376 24216 10382 24268
rect 10410 24216 10416 24268
rect 10468 24256 10474 24268
rect 10686 24256 10692 24268
rect 10744 24265 10750 24268
rect 10744 24259 10772 24265
rect 10468 24228 10692 24256
rect 10468 24216 10474 24228
rect 10686 24216 10692 24228
rect 10760 24225 10772 24259
rect 10744 24219 10772 24225
rect 10744 24216 10750 24219
rect 10870 24216 10876 24268
rect 10928 24216 10934 24268
rect 11348 24256 11376 24364
rect 11517 24361 11529 24395
rect 11563 24392 11575 24395
rect 11882 24392 11888 24404
rect 11563 24364 11888 24392
rect 11563 24361 11575 24364
rect 11517 24355 11575 24361
rect 11882 24352 11888 24364
rect 11940 24352 11946 24404
rect 13081 24327 13139 24333
rect 13081 24293 13093 24327
rect 13127 24324 13139 24327
rect 13446 24324 13452 24336
rect 13127 24296 13452 24324
rect 13127 24293 13139 24296
rect 13081 24287 13139 24293
rect 13446 24284 13452 24296
rect 13504 24284 13510 24336
rect 11348 24228 11468 24256
rect 7757 24160 8156 24188
rect 9677 24191 9735 24197
rect 7757 24157 7769 24160
rect 7711 24151 7769 24157
rect 9677 24157 9689 24191
rect 9723 24157 9735 24191
rect 9677 24151 9735 24157
rect 8662 24120 8668 24132
rect 6656 24092 8668 24120
rect 6656 24064 6684 24092
rect 8662 24080 8668 24092
rect 8720 24080 8726 24132
rect 6638 24012 6644 24064
rect 6696 24012 6702 24064
rect 8481 24055 8539 24061
rect 8481 24021 8493 24055
rect 8527 24052 8539 24055
rect 8846 24052 8852 24064
rect 8527 24024 8852 24052
rect 8527 24021 8539 24024
rect 8481 24015 8539 24021
rect 8846 24012 8852 24024
rect 8904 24012 8910 24064
rect 9692 24052 9720 24151
rect 9766 24148 9772 24200
rect 9824 24188 9830 24200
rect 9861 24191 9919 24197
rect 9861 24188 9873 24191
rect 9824 24160 9873 24188
rect 9824 24148 9830 24160
rect 9861 24157 9873 24160
rect 9907 24157 9919 24191
rect 9861 24151 9919 24157
rect 10594 24148 10600 24200
rect 10652 24148 10658 24200
rect 11440 24188 11468 24228
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 11609 24259 11667 24265
rect 11609 24256 11621 24259
rect 11572 24228 11621 24256
rect 11572 24216 11578 24228
rect 11609 24225 11621 24228
rect 11655 24225 11667 24259
rect 11609 24219 11667 24225
rect 13630 24216 13636 24268
rect 13688 24256 13694 24268
rect 13688 24228 14228 24256
rect 13688 24216 13694 24228
rect 11882 24197 11888 24200
rect 11851 24191 11888 24197
rect 11851 24188 11863 24191
rect 11440 24160 11863 24188
rect 11851 24157 11863 24160
rect 11851 24151 11888 24157
rect 11882 24148 11888 24151
rect 11940 24148 11946 24200
rect 13265 24191 13323 24197
rect 13265 24157 13277 24191
rect 13311 24188 13323 24191
rect 13814 24188 13820 24200
rect 13311 24160 13820 24188
rect 13311 24157 13323 24160
rect 13265 24151 13323 24157
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 14200 24197 14228 24228
rect 14185 24191 14243 24197
rect 14185 24157 14197 24191
rect 14231 24157 14243 24191
rect 14185 24151 14243 24157
rect 13541 24123 13599 24129
rect 13541 24089 13553 24123
rect 13587 24120 13599 24123
rect 13722 24120 13728 24132
rect 13587 24092 13728 24120
rect 13587 24089 13599 24092
rect 13541 24083 13599 24089
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 13909 24123 13967 24129
rect 13909 24089 13921 24123
rect 13955 24120 13967 24123
rect 15102 24120 15108 24132
rect 13955 24092 15108 24120
rect 13955 24089 13967 24092
rect 13909 24083 13967 24089
rect 15102 24080 15108 24092
rect 15160 24080 15166 24132
rect 10962 24052 10968 24064
rect 9692 24024 10968 24052
rect 10962 24012 10968 24024
rect 11020 24012 11026 24064
rect 12618 24012 12624 24064
rect 12676 24012 12682 24064
rect 14366 24012 14372 24064
rect 14424 24012 14430 24064
rect 1104 23962 14971 23984
rect 1104 23910 4376 23962
rect 4428 23910 4440 23962
rect 4492 23910 4504 23962
rect 4556 23910 4568 23962
rect 4620 23910 4632 23962
rect 4684 23910 7803 23962
rect 7855 23910 7867 23962
rect 7919 23910 7931 23962
rect 7983 23910 7995 23962
rect 8047 23910 8059 23962
rect 8111 23910 11230 23962
rect 11282 23910 11294 23962
rect 11346 23910 11358 23962
rect 11410 23910 11422 23962
rect 11474 23910 11486 23962
rect 11538 23910 14657 23962
rect 14709 23910 14721 23962
rect 14773 23910 14785 23962
rect 14837 23910 14849 23962
rect 14901 23910 14913 23962
rect 14965 23910 14971 23962
rect 1104 23888 14971 23910
rect 4982 23808 4988 23860
rect 5040 23848 5046 23860
rect 9858 23848 9864 23860
rect 5040 23820 9864 23848
rect 5040 23808 5046 23820
rect 9858 23808 9864 23820
rect 9916 23808 9922 23860
rect 10137 23851 10195 23857
rect 10137 23817 10149 23851
rect 10183 23848 10195 23851
rect 10318 23848 10324 23860
rect 10183 23820 10324 23848
rect 10183 23817 10195 23820
rect 10137 23811 10195 23817
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 10686 23808 10692 23860
rect 10744 23848 10750 23860
rect 12342 23848 12348 23860
rect 10744 23820 12348 23848
rect 10744 23808 10750 23820
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 8110 23780 8116 23792
rect 1688 23752 8116 23780
rect 1688 23721 1716 23752
rect 8110 23740 8116 23752
rect 8168 23740 8174 23792
rect 8570 23740 8576 23792
rect 8628 23780 8634 23792
rect 8628 23752 9720 23780
rect 8628 23740 8634 23752
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 6454 23672 6460 23724
rect 6512 23712 6518 23724
rect 7191 23715 7249 23721
rect 7191 23712 7203 23715
rect 6512 23684 7203 23712
rect 6512 23672 6518 23684
rect 7191 23681 7203 23684
rect 7237 23712 7249 23715
rect 9367 23715 9425 23721
rect 9367 23712 9379 23715
rect 7237 23684 7604 23712
rect 7237 23681 7249 23684
rect 7191 23675 7249 23681
rect 750 23604 756 23656
rect 808 23644 814 23656
rect 1397 23647 1455 23653
rect 1397 23644 1409 23647
rect 808 23616 1409 23644
rect 808 23604 814 23616
rect 1397 23613 1409 23616
rect 1443 23613 1455 23647
rect 1397 23607 1455 23613
rect 6914 23604 6920 23656
rect 6972 23604 6978 23656
rect 7576 23644 7604 23684
rect 8496 23684 9379 23712
rect 8496 23644 8524 23684
rect 9367 23681 9379 23684
rect 9413 23681 9425 23715
rect 9692 23712 9720 23752
rect 13722 23740 13728 23792
rect 13780 23780 13786 23792
rect 14093 23783 14151 23789
rect 14093 23780 14105 23783
rect 13780 23752 14105 23780
rect 13780 23740 13786 23752
rect 14093 23749 14105 23752
rect 14139 23749 14151 23783
rect 14093 23743 14151 23749
rect 9692 23684 10364 23712
rect 9367 23675 9425 23681
rect 7576 23616 8524 23644
rect 9122 23604 9128 23656
rect 9180 23604 9186 23656
rect 9950 23604 9956 23656
rect 10008 23604 10014 23656
rect 10336 23644 10364 23684
rect 11974 23672 11980 23724
rect 12032 23712 12038 23724
rect 12032 23684 12388 23712
rect 12032 23672 12038 23684
rect 12360 23656 12388 23684
rect 13170 23672 13176 23724
rect 13228 23672 13234 23724
rect 11698 23644 11704 23656
rect 10336 23616 11704 23644
rect 11698 23604 11704 23616
rect 11756 23644 11762 23656
rect 12161 23647 12219 23653
rect 12161 23644 12173 23647
rect 11756 23616 12173 23644
rect 11756 23604 11762 23616
rect 12161 23613 12173 23616
rect 12207 23613 12219 23647
rect 12161 23607 12219 23613
rect 12342 23604 12348 23656
rect 12400 23604 12406 23656
rect 12618 23604 12624 23656
rect 12676 23604 12682 23656
rect 12897 23647 12955 23653
rect 12897 23644 12909 23647
rect 12726 23616 12909 23644
rect 9140 23576 9168 23604
rect 7852 23548 9168 23576
rect 9968 23576 9996 23604
rect 12726 23576 12754 23616
rect 12897 23613 12909 23616
rect 12943 23613 12955 23647
rect 12897 23607 12955 23613
rect 12986 23604 12992 23656
rect 13044 23653 13050 23656
rect 13044 23647 13072 23653
rect 13060 23613 13072 23647
rect 13044 23607 13072 23613
rect 13044 23604 13050 23607
rect 9968 23548 12754 23576
rect 7190 23468 7196 23520
rect 7248 23508 7254 23520
rect 7852 23508 7880 23548
rect 7248 23480 7880 23508
rect 7929 23511 7987 23517
rect 7248 23468 7254 23480
rect 7929 23477 7941 23511
rect 7975 23508 7987 23511
rect 8202 23508 8208 23520
rect 7975 23480 8208 23508
rect 7975 23477 7987 23480
rect 7929 23471 7987 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 9398 23468 9404 23520
rect 9456 23508 9462 23520
rect 10870 23508 10876 23520
rect 9456 23480 10876 23508
rect 9456 23468 9462 23480
rect 10870 23468 10876 23480
rect 10928 23468 10934 23520
rect 12726 23508 12754 23548
rect 13262 23508 13268 23520
rect 12726 23480 13268 23508
rect 13262 23468 13268 23480
rect 13320 23468 13326 23520
rect 13354 23468 13360 23520
rect 13412 23508 13418 23520
rect 13817 23511 13875 23517
rect 13817 23508 13829 23511
rect 13412 23480 13829 23508
rect 13412 23468 13418 23480
rect 13817 23477 13829 23480
rect 13863 23477 13875 23511
rect 13817 23471 13875 23477
rect 14366 23468 14372 23520
rect 14424 23468 14430 23520
rect 1104 23418 14812 23440
rect 1104 23366 2663 23418
rect 2715 23366 2727 23418
rect 2779 23366 2791 23418
rect 2843 23366 2855 23418
rect 2907 23366 2919 23418
rect 2971 23366 6090 23418
rect 6142 23366 6154 23418
rect 6206 23366 6218 23418
rect 6270 23366 6282 23418
rect 6334 23366 6346 23418
rect 6398 23366 9517 23418
rect 9569 23366 9581 23418
rect 9633 23366 9645 23418
rect 9697 23366 9709 23418
rect 9761 23366 9773 23418
rect 9825 23366 12944 23418
rect 12996 23366 13008 23418
rect 13060 23366 13072 23418
rect 13124 23366 13136 23418
rect 13188 23366 13200 23418
rect 13252 23366 14812 23418
rect 1104 23344 14812 23366
rect 5442 23264 5448 23316
rect 5500 23304 5506 23316
rect 6914 23304 6920 23316
rect 5500 23276 6920 23304
rect 5500 23264 5506 23276
rect 6914 23264 6920 23276
rect 6972 23304 6978 23316
rect 6972 23276 8524 23304
rect 6972 23264 6978 23276
rect 8496 23248 8524 23276
rect 9122 23264 9128 23316
rect 9180 23304 9186 23316
rect 9950 23304 9956 23316
rect 9180 23276 9956 23304
rect 9180 23264 9186 23276
rect 9950 23264 9956 23276
rect 10008 23264 10014 23316
rect 11146 23304 11152 23316
rect 10888 23276 11152 23304
rect 5261 23239 5319 23245
rect 5261 23205 5273 23239
rect 5307 23236 5319 23239
rect 6273 23239 6331 23245
rect 6273 23236 6285 23239
rect 5307 23208 6285 23236
rect 5307 23205 5319 23208
rect 5261 23199 5319 23205
rect 6273 23205 6285 23208
rect 6319 23205 6331 23239
rect 6273 23199 6331 23205
rect 8478 23196 8484 23248
rect 8536 23196 8542 23248
rect 6546 23128 6552 23180
rect 6604 23128 6610 23180
rect 6730 23177 6736 23180
rect 6687 23171 6736 23177
rect 6687 23137 6699 23171
rect 6733 23137 6736 23171
rect 6687 23131 6736 23137
rect 6730 23128 6736 23131
rect 6788 23128 6794 23180
rect 4246 23060 4252 23112
rect 4304 23060 4310 23112
rect 4523 23103 4581 23109
rect 4523 23069 4535 23103
rect 4569 23100 4581 23103
rect 5166 23100 5172 23112
rect 4569 23072 5172 23100
rect 4569 23069 4581 23072
rect 4523 23063 4581 23069
rect 5166 23060 5172 23072
rect 5224 23060 5230 23112
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5718 23100 5724 23112
rect 5675 23072 5724 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 750 22992 756 23044
rect 808 23032 814 23044
rect 1489 23035 1547 23041
rect 1489 23032 1501 23035
rect 808 23004 1501 23032
rect 808 22992 814 23004
rect 1489 23001 1501 23004
rect 1535 23001 1547 23035
rect 1489 22995 1547 23001
rect 1578 22924 1584 22976
rect 1636 22924 1642 22976
rect 5644 22964 5672 23063
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5810 23060 5816 23112
rect 5868 23060 5874 23112
rect 6822 23060 6828 23112
rect 6880 23060 6886 23112
rect 8496 23100 8524 23196
rect 10888 23177 10916 23276
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 13357 23307 13415 23313
rect 13357 23273 13369 23307
rect 13403 23304 13415 23307
rect 13722 23304 13728 23316
rect 13403 23276 13728 23304
rect 13403 23273 13415 23276
rect 13357 23267 13415 23273
rect 13722 23264 13728 23276
rect 13780 23264 13786 23316
rect 13081 23239 13139 23245
rect 13081 23205 13093 23239
rect 13127 23236 13139 23239
rect 13630 23236 13636 23248
rect 13127 23208 13636 23236
rect 13127 23205 13139 23208
rect 13081 23199 13139 23205
rect 13630 23196 13636 23208
rect 13688 23196 13694 23248
rect 14366 23196 14372 23248
rect 14424 23196 14430 23248
rect 10873 23171 10931 23177
rect 10873 23137 10885 23171
rect 10919 23137 10931 23171
rect 10873 23131 10931 23137
rect 9122 23100 9128 23112
rect 8496 23072 9128 23100
rect 9122 23060 9128 23072
rect 9180 23100 9186 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 9180 23072 9505 23100
rect 9180 23060 9186 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9766 23060 9772 23112
rect 9824 23070 9830 23112
rect 9824 23060 9904 23070
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 11790 23060 11796 23112
rect 11848 23100 11854 23112
rect 12802 23100 12808 23112
rect 11848 23072 12808 23100
rect 11848 23060 11854 23072
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 13265 23103 13323 23109
rect 13265 23069 13277 23103
rect 13311 23100 13323 23103
rect 13354 23100 13360 23112
rect 13311 23072 13360 23100
rect 13311 23069 13323 23072
rect 13265 23063 13323 23069
rect 13354 23060 13360 23072
rect 13412 23060 13418 23112
rect 13446 23060 13452 23112
rect 13504 23100 13510 23112
rect 13541 23103 13599 23109
rect 13541 23100 13553 23103
rect 13504 23072 13553 23100
rect 13504 23060 13510 23072
rect 13541 23069 13553 23072
rect 13587 23069 13599 23103
rect 13541 23063 13599 23069
rect 13630 23060 13636 23112
rect 13688 23060 13694 23112
rect 14185 23103 14243 23109
rect 14185 23069 14197 23103
rect 14231 23100 14243 23103
rect 14274 23100 14280 23112
rect 14231 23072 14280 23100
rect 14231 23069 14243 23072
rect 14185 23063 14243 23069
rect 14274 23060 14280 23072
rect 14332 23060 14338 23112
rect 9767 23059 9779 23060
rect 9813 23059 9904 23060
rect 9767 23053 9904 23059
rect 7469 23035 7527 23041
rect 7469 23001 7481 23035
rect 7515 23032 7527 23035
rect 8478 23032 8484 23044
rect 7515 23004 8484 23032
rect 7515 23001 7527 23004
rect 7469 22995 7527 23001
rect 8478 22992 8484 23004
rect 8536 22992 8542 23044
rect 9784 23042 9904 23053
rect 9876 23032 9904 23042
rect 10042 23032 10048 23044
rect 9876 23004 10048 23032
rect 10042 22992 10048 23004
rect 10100 22992 10106 23044
rect 13906 22992 13912 23044
rect 13964 23032 13970 23044
rect 15930 23032 15936 23044
rect 13964 23004 15936 23032
rect 13964 22992 13970 23004
rect 15930 22992 15936 23004
rect 15988 22992 15994 23044
rect 6914 22964 6920 22976
rect 5644 22936 6920 22964
rect 6914 22924 6920 22936
rect 6972 22924 6978 22976
rect 8110 22924 8116 22976
rect 8168 22964 8174 22976
rect 9582 22964 9588 22976
rect 8168 22936 9588 22964
rect 8168 22924 8174 22936
rect 9582 22924 9588 22936
rect 9640 22924 9646 22976
rect 10505 22967 10563 22973
rect 10505 22933 10517 22967
rect 10551 22964 10563 22967
rect 10870 22964 10876 22976
rect 10551 22936 10876 22964
rect 10551 22933 10563 22936
rect 10505 22927 10563 22933
rect 10870 22924 10876 22936
rect 10928 22924 10934 22976
rect 11882 22924 11888 22976
rect 11940 22924 11946 22976
rect 13817 22967 13875 22973
rect 13817 22933 13829 22967
rect 13863 22964 13875 22967
rect 15102 22964 15108 22976
rect 13863 22936 15108 22964
rect 13863 22933 13875 22936
rect 13817 22927 13875 22933
rect 15102 22924 15108 22936
rect 15160 22924 15166 22976
rect 1104 22874 14971 22896
rect 1104 22822 4376 22874
rect 4428 22822 4440 22874
rect 4492 22822 4504 22874
rect 4556 22822 4568 22874
rect 4620 22822 4632 22874
rect 4684 22822 7803 22874
rect 7855 22822 7867 22874
rect 7919 22822 7931 22874
rect 7983 22822 7995 22874
rect 8047 22822 8059 22874
rect 8111 22822 11230 22874
rect 11282 22822 11294 22874
rect 11346 22822 11358 22874
rect 11410 22822 11422 22874
rect 11474 22822 11486 22874
rect 11538 22822 14657 22874
rect 14709 22822 14721 22874
rect 14773 22822 14785 22874
rect 14837 22822 14849 22874
rect 14901 22822 14913 22874
rect 14965 22822 14971 22874
rect 1104 22800 14971 22822
rect 1578 22720 1584 22772
rect 1636 22760 1642 22772
rect 10686 22760 10692 22772
rect 1636 22732 10692 22760
rect 1636 22720 1642 22732
rect 10686 22720 10692 22732
rect 10744 22760 10750 22772
rect 11146 22760 11152 22772
rect 10744 22732 11152 22760
rect 10744 22720 10750 22732
rect 11146 22720 11152 22732
rect 11204 22720 11210 22772
rect 13265 22763 13323 22769
rect 13265 22729 13277 22763
rect 13311 22760 13323 22763
rect 13630 22760 13636 22772
rect 13311 22732 13636 22760
rect 13311 22729 13323 22732
rect 13265 22723 13323 22729
rect 13630 22720 13636 22732
rect 13688 22720 13694 22772
rect 14274 22720 14280 22772
rect 14332 22720 14338 22772
rect 14090 22692 14096 22704
rect 13188 22664 14096 22692
rect 5074 22584 5080 22636
rect 5132 22624 5138 22636
rect 5994 22624 6000 22636
rect 5132 22596 6000 22624
rect 5132 22584 5138 22596
rect 5994 22584 6000 22596
rect 6052 22584 6058 22636
rect 7190 22584 7196 22636
rect 7248 22624 7254 22636
rect 7558 22624 7564 22636
rect 7248 22596 7564 22624
rect 7248 22584 7254 22596
rect 7558 22584 7564 22596
rect 7616 22624 7622 22636
rect 7653 22627 7711 22633
rect 7653 22624 7665 22627
rect 7616 22596 7665 22624
rect 7616 22584 7622 22596
rect 7653 22593 7665 22596
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 13188 22633 13216 22664
rect 14090 22652 14096 22664
rect 14148 22652 14154 22704
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22593 13231 22627
rect 13173 22587 13231 22593
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 13722 22584 13728 22636
rect 13780 22584 13786 22636
rect 13906 22584 13912 22636
rect 13964 22584 13970 22636
rect 7837 22559 7895 22565
rect 7837 22525 7849 22559
rect 7883 22525 7895 22559
rect 7837 22519 7895 22525
rect 6638 22448 6644 22500
rect 6696 22488 6702 22500
rect 7852 22488 7880 22519
rect 8202 22516 8208 22568
rect 8260 22556 8266 22568
rect 8297 22559 8355 22565
rect 8297 22556 8309 22559
rect 8260 22528 8309 22556
rect 8260 22516 8266 22528
rect 8297 22525 8309 22528
rect 8343 22525 8355 22559
rect 8297 22519 8355 22525
rect 8570 22516 8576 22568
rect 8628 22516 8634 22568
rect 8662 22516 8668 22568
rect 8720 22565 8726 22568
rect 8720 22559 8748 22565
rect 8736 22525 8748 22559
rect 8720 22519 8748 22525
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22556 9551 22559
rect 13998 22556 14004 22568
rect 9539 22528 14004 22556
rect 9539 22525 9551 22528
rect 9493 22519 9551 22525
rect 8720 22516 8726 22519
rect 13998 22516 14004 22528
rect 14056 22516 14062 22568
rect 13354 22488 13360 22500
rect 6696 22460 7880 22488
rect 12636 22460 13360 22488
rect 6696 22448 6702 22460
rect 12636 22432 12664 22460
rect 13354 22448 13360 22460
rect 13412 22448 13418 22500
rect 13541 22491 13599 22497
rect 13541 22457 13553 22491
rect 13587 22488 13599 22491
rect 14292 22488 14320 22720
rect 13587 22460 14320 22488
rect 13587 22457 13599 22460
rect 13541 22451 13599 22457
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 12618 22420 12624 22432
rect 5868 22392 12624 22420
rect 5868 22380 5874 22392
rect 12618 22380 12624 22392
rect 12676 22380 12682 22432
rect 12989 22423 13047 22429
rect 12989 22389 13001 22423
rect 13035 22420 13047 22423
rect 13998 22420 14004 22432
rect 13035 22392 14004 22420
rect 13035 22389 13047 22392
rect 12989 22383 13047 22389
rect 13998 22380 14004 22392
rect 14056 22380 14062 22432
rect 14185 22423 14243 22429
rect 14185 22389 14197 22423
rect 14231 22420 14243 22423
rect 14918 22420 14924 22432
rect 14231 22392 14924 22420
rect 14231 22389 14243 22392
rect 14185 22383 14243 22389
rect 14918 22380 14924 22392
rect 14976 22380 14982 22432
rect 1104 22330 14812 22352
rect 1104 22278 2663 22330
rect 2715 22278 2727 22330
rect 2779 22278 2791 22330
rect 2843 22278 2855 22330
rect 2907 22278 2919 22330
rect 2971 22278 6090 22330
rect 6142 22278 6154 22330
rect 6206 22278 6218 22330
rect 6270 22278 6282 22330
rect 6334 22278 6346 22330
rect 6398 22278 9517 22330
rect 9569 22278 9581 22330
rect 9633 22278 9645 22330
rect 9697 22278 9709 22330
rect 9761 22278 9773 22330
rect 9825 22278 12944 22330
rect 12996 22278 13008 22330
rect 13060 22278 13072 22330
rect 13124 22278 13136 22330
rect 13188 22278 13200 22330
rect 13252 22278 14812 22330
rect 1104 22256 14812 22278
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6822 22216 6828 22228
rect 6503 22188 6828 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 9582 22216 9588 22228
rect 6972 22188 9588 22216
rect 6972 22176 6978 22188
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10686 22216 10692 22228
rect 10008 22188 10692 22216
rect 10008 22176 10014 22188
rect 10226 22108 10232 22160
rect 10284 22108 10290 22160
rect 4246 22040 4252 22092
rect 4304 22080 4310 22092
rect 5442 22080 5448 22092
rect 4304 22052 5448 22080
rect 4304 22040 4310 22052
rect 5442 22040 5448 22052
rect 5500 22040 5506 22092
rect 9674 22040 9680 22092
rect 9732 22080 9738 22092
rect 10244 22080 10272 22108
rect 10428 22089 10456 22188
rect 10686 22176 10692 22188
rect 10744 22176 10750 22228
rect 11425 22219 11483 22225
rect 11425 22185 11437 22219
rect 11471 22216 11483 22219
rect 13170 22216 13176 22228
rect 11471 22188 12480 22216
rect 11471 22185 11483 22188
rect 11425 22179 11483 22185
rect 12452 22157 12480 22188
rect 12544 22188 13176 22216
rect 12437 22151 12495 22157
rect 12437 22117 12449 22151
rect 12483 22117 12495 22151
rect 12437 22111 12495 22117
rect 9732 22052 10272 22080
rect 10413 22083 10471 22089
rect 9732 22040 9738 22052
rect 10060 22024 10088 22052
rect 10413 22049 10425 22083
rect 10459 22049 10471 22083
rect 12066 22080 12072 22092
rect 10413 22043 10471 22049
rect 11348 22052 12072 22080
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 1673 21975 1731 21981
rect 750 21904 756 21956
rect 808 21944 814 21956
rect 1489 21947 1547 21953
rect 1489 21944 1501 21947
rect 808 21916 1501 21944
rect 808 21904 814 21916
rect 1489 21913 1501 21916
rect 1535 21913 1547 21947
rect 1688 21944 1716 21975
rect 3142 21972 3148 22024
rect 3200 21972 3206 22024
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 5719 22015 5777 22021
rect 5719 22012 5731 22015
rect 5684 21984 5731 22012
rect 5684 21972 5690 21984
rect 5719 21981 5731 21984
rect 5765 22012 5777 22015
rect 6270 22012 6276 22024
rect 5765 21984 6276 22012
rect 5765 21981 5777 21984
rect 5719 21975 5777 21981
rect 6270 21972 6276 21984
rect 6328 21972 6334 22024
rect 6454 21972 6460 22024
rect 6512 22012 6518 22024
rect 6822 22012 6828 22024
rect 6512 21984 6828 22012
rect 6512 21972 6518 21984
rect 6822 21972 6828 21984
rect 6880 21972 6886 22024
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 7099 22015 7157 22021
rect 7099 22012 7111 22015
rect 7064 21984 7111 22012
rect 7064 21972 7070 21984
rect 7099 21981 7111 21984
rect 7145 21981 7157 22015
rect 9950 22012 9956 22024
rect 7099 21975 7157 21981
rect 8404 21984 9956 22012
rect 8404 21944 8432 21984
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 10042 21972 10048 22024
rect 10100 21972 10106 22024
rect 10687 22015 10745 22021
rect 10687 22012 10699 22015
rect 10612 21984 10699 22012
rect 1688 21916 8432 21944
rect 1489 21907 1547 21913
rect 9490 21904 9496 21956
rect 9548 21944 9554 21956
rect 10612 21944 10640 21984
rect 10687 21981 10699 21984
rect 10733 22012 10745 22015
rect 11348 22012 11376 22052
rect 12066 22040 12072 22052
rect 12124 22040 12130 22092
rect 12544 22080 12572 22188
rect 13170 22176 13176 22188
rect 13228 22176 13234 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13633 22219 13691 22225
rect 13633 22216 13645 22219
rect 13596 22188 13645 22216
rect 13596 22176 13602 22188
rect 13633 22185 13645 22188
rect 13679 22185 13691 22219
rect 13633 22179 13691 22185
rect 14369 22219 14427 22225
rect 14369 22185 14381 22219
rect 14415 22216 14427 22219
rect 14458 22216 14464 22228
rect 14415 22188 14464 22216
rect 14415 22185 14427 22188
rect 14369 22179 14427 22185
rect 14458 22176 14464 22188
rect 14516 22176 14522 22228
rect 12713 22083 12771 22089
rect 12713 22080 12725 22083
rect 12544 22052 12725 22080
rect 12713 22049 12725 22052
rect 12759 22049 12771 22083
rect 12713 22043 12771 22049
rect 12878 22052 13584 22080
rect 12878 22024 12906 22052
rect 10733 21984 11376 22012
rect 10733 21981 10745 21984
rect 10687 21975 10745 21981
rect 11698 21972 11704 22024
rect 11756 21972 11762 22024
rect 11790 21972 11796 22024
rect 11848 21972 11854 22024
rect 12878 22021 12900 22024
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12851 22015 12900 22021
rect 12851 21981 12863 22015
rect 12897 21981 12900 22015
rect 12851 21975 12900 21981
rect 9548 21916 10640 21944
rect 11716 21944 11744 21972
rect 11992 21944 12020 21975
rect 12894 21972 12900 21975
rect 12952 21972 12958 22024
rect 12986 21972 12992 22024
rect 13044 21972 13050 22024
rect 11716 21916 12020 21944
rect 13556 21944 13584 22052
rect 14090 22040 14096 22092
rect 14148 22080 14154 22092
rect 15194 22080 15200 22092
rect 14148 22052 15200 22080
rect 14148 22040 14154 22052
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15286 22040 15292 22092
rect 15344 22080 15350 22092
rect 15344 22052 15792 22080
rect 15344 22040 15350 22052
rect 13906 21972 13912 22024
rect 13964 21972 13970 22024
rect 13998 21972 14004 22024
rect 14056 22012 14062 22024
rect 14185 22015 14243 22021
rect 14185 22012 14197 22015
rect 14056 21984 14197 22012
rect 14056 21972 14062 21984
rect 14185 21981 14197 21984
rect 14231 21981 14243 22015
rect 14185 21975 14243 21981
rect 13556 21916 14044 21944
rect 9548 21904 9554 21916
rect 14016 21888 14044 21916
rect 15102 21904 15108 21956
rect 15160 21904 15166 21956
rect 15764 21944 15792 22052
rect 15764 21916 15884 21944
rect 3326 21836 3332 21888
rect 3384 21836 3390 21888
rect 7837 21879 7895 21885
rect 7837 21845 7849 21879
rect 7883 21876 7895 21879
rect 8202 21876 8208 21888
rect 7883 21848 8208 21876
rect 7883 21845 7895 21848
rect 7837 21839 7895 21845
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 9582 21836 9588 21888
rect 9640 21876 9646 21888
rect 12894 21876 12900 21888
rect 9640 21848 12900 21876
rect 9640 21836 9646 21848
rect 12894 21836 12900 21848
rect 12952 21836 12958 21888
rect 13078 21836 13084 21888
rect 13136 21876 13142 21888
rect 13725 21879 13783 21885
rect 13725 21876 13737 21879
rect 13136 21848 13737 21876
rect 13136 21836 13142 21848
rect 13725 21845 13737 21848
rect 13771 21845 13783 21879
rect 13725 21839 13783 21845
rect 13998 21836 14004 21888
rect 14056 21836 14062 21888
rect 15120 21808 15148 21904
rect 15856 21888 15884 21916
rect 15838 21836 15844 21888
rect 15896 21836 15902 21888
rect 1104 21786 14971 21808
rect 1104 21734 4376 21786
rect 4428 21734 4440 21786
rect 4492 21734 4504 21786
rect 4556 21734 4568 21786
rect 4620 21734 4632 21786
rect 4684 21734 7803 21786
rect 7855 21734 7867 21786
rect 7919 21734 7931 21786
rect 7983 21734 7995 21786
rect 8047 21734 8059 21786
rect 8111 21734 11230 21786
rect 11282 21734 11294 21786
rect 11346 21734 11358 21786
rect 11410 21734 11422 21786
rect 11474 21734 11486 21786
rect 11538 21734 14657 21786
rect 14709 21734 14721 21786
rect 14773 21734 14785 21786
rect 14837 21734 14849 21786
rect 14901 21734 14913 21786
rect 14965 21734 14971 21786
rect 15120 21780 15424 21808
rect 15396 21752 15424 21780
rect 1104 21712 14971 21734
rect 15378 21700 15384 21752
rect 15436 21700 15442 21752
rect 2682 21632 2688 21684
rect 2740 21632 2746 21684
rect 3142 21632 3148 21684
rect 3200 21672 3206 21684
rect 3237 21675 3295 21681
rect 3237 21672 3249 21675
rect 3200 21644 3249 21672
rect 3200 21632 3206 21644
rect 3237 21641 3249 21644
rect 3283 21641 3295 21675
rect 3237 21635 3295 21641
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5534 21672 5540 21684
rect 5132 21644 5540 21672
rect 5132 21632 5138 21644
rect 5534 21632 5540 21644
rect 5592 21632 5598 21684
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 8386 21672 8392 21684
rect 6604 21644 8392 21672
rect 6604 21632 6610 21644
rect 8386 21632 8392 21644
rect 8444 21632 8450 21684
rect 8478 21632 8484 21684
rect 8536 21672 8542 21684
rect 9309 21675 9367 21681
rect 8536 21644 9168 21672
rect 8536 21632 8542 21644
rect 1397 21607 1455 21613
rect 1397 21573 1409 21607
rect 1443 21604 1455 21607
rect 4154 21604 4160 21616
rect 1443 21576 4160 21604
rect 1443 21573 1455 21576
rect 1397 21567 1455 21573
rect 4154 21564 4160 21576
rect 4212 21564 4218 21616
rect 7190 21564 7196 21616
rect 7248 21604 7254 21616
rect 7374 21604 7380 21616
rect 7248 21576 7380 21604
rect 7248 21564 7254 21576
rect 7374 21564 7380 21576
rect 7432 21564 7438 21616
rect 9140 21604 9168 21644
rect 9309 21641 9321 21675
rect 9355 21672 9367 21675
rect 9398 21672 9404 21684
rect 9355 21644 9404 21672
rect 9355 21641 9367 21644
rect 9309 21635 9367 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 9858 21672 9864 21684
rect 9508 21644 9864 21672
rect 9508 21604 9536 21644
rect 9858 21632 9864 21644
rect 9916 21632 9922 21684
rect 10134 21632 10140 21684
rect 10192 21632 10198 21684
rect 12713 21675 12771 21681
rect 12713 21641 12725 21675
rect 12759 21672 12771 21675
rect 12986 21672 12992 21684
rect 12759 21644 12992 21672
rect 12759 21641 12771 21644
rect 12713 21635 12771 21641
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 13265 21675 13323 21681
rect 13265 21641 13277 21675
rect 13311 21672 13323 21675
rect 14274 21672 14280 21684
rect 13311 21644 14280 21672
rect 13311 21641 13323 21644
rect 13265 21635 13323 21641
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 14369 21675 14427 21681
rect 14369 21641 14381 21675
rect 14415 21672 14427 21675
rect 14458 21672 14464 21684
rect 14415 21644 14464 21672
rect 14415 21641 14427 21644
rect 14369 21635 14427 21641
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 9140 21576 9536 21604
rect 11959 21569 12017 21575
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21536 3479 21539
rect 5626 21536 5632 21548
rect 3467 21508 5632 21536
rect 3467 21505 3479 21508
rect 3421 21499 3479 21505
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 7469 21539 7527 21545
rect 7469 21505 7481 21539
rect 7515 21505 7527 21539
rect 7469 21499 7527 21505
rect 6270 21428 6276 21480
rect 6328 21468 6334 21480
rect 6822 21468 6828 21480
rect 6328 21440 6828 21468
rect 6328 21428 6334 21440
rect 6822 21428 6828 21440
rect 6880 21428 6886 21480
rect 2130 21360 2136 21412
rect 2188 21400 2194 21412
rect 7374 21400 7380 21412
rect 2188 21372 7380 21400
rect 2188 21360 2194 21372
rect 7374 21360 7380 21372
rect 7432 21360 7438 21412
rect 7484 21400 7512 21499
rect 8386 21496 8392 21548
rect 8444 21496 8450 21548
rect 8478 21496 8484 21548
rect 8536 21545 8542 21548
rect 8536 21539 8564 21545
rect 8552 21505 8564 21539
rect 8536 21499 8564 21505
rect 8536 21496 8542 21499
rect 8662 21496 8668 21548
rect 8720 21496 8726 21548
rect 9398 21496 9404 21548
rect 9456 21536 9462 21548
rect 9456 21508 9904 21536
rect 9456 21496 9462 21508
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7616 21440 7665 21468
rect 7616 21428 7622 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 8110 21428 8116 21480
rect 8168 21428 8174 21480
rect 9876 21468 9904 21508
rect 9950 21496 9956 21548
rect 10008 21536 10014 21548
rect 10045 21539 10103 21545
rect 10045 21536 10057 21539
rect 10008 21508 10057 21536
rect 10008 21496 10014 21508
rect 10045 21505 10057 21508
rect 10091 21505 10103 21539
rect 10321 21539 10379 21545
rect 10321 21536 10333 21539
rect 10045 21499 10103 21505
rect 10244 21508 10333 21536
rect 10244 21468 10272 21508
rect 10321 21505 10333 21508
rect 10367 21536 10379 21539
rect 10594 21536 10600 21548
rect 10367 21508 10600 21536
rect 10367 21505 10379 21508
rect 10321 21499 10379 21505
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 10686 21496 10692 21548
rect 10744 21536 10750 21548
rect 11701 21539 11759 21545
rect 11701 21536 11713 21539
rect 10744 21508 11713 21536
rect 10744 21496 10750 21508
rect 11701 21505 11713 21508
rect 11747 21505 11759 21539
rect 11959 21535 11971 21569
rect 12005 21566 12017 21569
rect 12005 21536 12020 21566
rect 12342 21536 12348 21548
rect 12005 21535 12348 21536
rect 11959 21529 12348 21535
rect 11992 21508 12348 21529
rect 11701 21499 11759 21505
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 13078 21496 13084 21548
rect 13136 21496 13142 21548
rect 13354 21496 13360 21548
rect 13412 21536 13418 21548
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 13412 21508 13553 21536
rect 13412 21496 13418 21508
rect 13541 21505 13553 21508
rect 13587 21505 13599 21539
rect 13541 21499 13599 21505
rect 14090 21496 14096 21548
rect 14148 21496 14154 21548
rect 8220 21440 9720 21468
rect 9876 21440 10272 21468
rect 12360 21468 12388 21496
rect 14182 21468 14188 21480
rect 12360 21440 14188 21468
rect 8220 21400 8248 21440
rect 7484 21372 8248 21400
rect 9692 21400 9720 21440
rect 14182 21428 14188 21440
rect 14240 21428 14246 21480
rect 9692 21372 10180 21400
rect 5442 21292 5448 21344
rect 5500 21332 5506 21344
rect 9674 21332 9680 21344
rect 5500 21304 9680 21332
rect 5500 21292 5506 21304
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 9858 21292 9864 21344
rect 9916 21292 9922 21344
rect 10152 21332 10180 21372
rect 11238 21332 11244 21344
rect 10152 21304 11244 21332
rect 11238 21292 11244 21304
rect 11296 21292 11302 21344
rect 11698 21292 11704 21344
rect 11756 21332 11762 21344
rect 12066 21332 12072 21344
rect 11756 21304 12072 21332
rect 11756 21292 11762 21304
rect 12066 21292 12072 21304
rect 12124 21292 12130 21344
rect 13814 21292 13820 21344
rect 13872 21292 13878 21344
rect 1104 21242 14812 21264
rect 1104 21190 2663 21242
rect 2715 21190 2727 21242
rect 2779 21190 2791 21242
rect 2843 21190 2855 21242
rect 2907 21190 2919 21242
rect 2971 21190 6090 21242
rect 6142 21190 6154 21242
rect 6206 21190 6218 21242
rect 6270 21190 6282 21242
rect 6334 21190 6346 21242
rect 6398 21190 9517 21242
rect 9569 21190 9581 21242
rect 9633 21190 9645 21242
rect 9697 21190 9709 21242
rect 9761 21190 9773 21242
rect 9825 21190 12944 21242
rect 12996 21190 13008 21242
rect 13060 21190 13072 21242
rect 13124 21190 13136 21242
rect 13188 21190 13200 21242
rect 13252 21190 14812 21242
rect 1104 21168 14812 21190
rect 1581 21131 1639 21137
rect 1581 21097 1593 21131
rect 1627 21128 1639 21131
rect 5442 21128 5448 21140
rect 1627 21100 5448 21128
rect 1627 21097 1639 21100
rect 1581 21091 1639 21097
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 5813 21131 5871 21137
rect 5813 21097 5825 21131
rect 5859 21128 5871 21131
rect 8481 21131 8539 21137
rect 5859 21100 8432 21128
rect 5859 21097 5871 21100
rect 5813 21091 5871 21097
rect 8404 21060 8432 21100
rect 8481 21097 8493 21131
rect 8527 21128 8539 21131
rect 8662 21128 8668 21140
rect 8527 21100 8668 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 8662 21088 8668 21100
rect 8720 21088 8726 21140
rect 9585 21131 9643 21137
rect 9585 21097 9597 21131
rect 9631 21128 9643 21131
rect 9631 21100 9720 21128
rect 9631 21097 9643 21100
rect 9585 21091 9643 21097
rect 9398 21060 9404 21072
rect 8404 21032 9404 21060
rect 9398 21020 9404 21032
rect 9456 21020 9462 21072
rect 4154 20952 4160 21004
rect 4212 20992 4218 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4212 20964 4445 20992
rect 4212 20952 4218 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5626 20952 5632 21004
rect 5684 20992 5690 21004
rect 5905 20995 5963 21001
rect 5905 20992 5917 20995
rect 5684 20964 5917 20992
rect 5684 20952 5690 20964
rect 5905 20961 5917 20964
rect 5951 20961 5963 20995
rect 5905 20955 5963 20961
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7469 20995 7527 21001
rect 7469 20992 7481 20995
rect 6972 20964 7481 20992
rect 6972 20952 6978 20964
rect 750 20884 756 20936
rect 808 20924 814 20936
rect 1489 20927 1547 20933
rect 1489 20924 1501 20927
rect 808 20896 1501 20924
rect 808 20884 814 20896
rect 1489 20893 1501 20896
rect 1535 20893 1547 20927
rect 1489 20887 1547 20893
rect 5810 20884 5816 20936
rect 5868 20924 5874 20936
rect 6147 20927 6205 20933
rect 6147 20924 6159 20927
rect 5868 20896 6159 20924
rect 5868 20884 5874 20896
rect 6147 20893 6159 20896
rect 6193 20893 6205 20927
rect 7006 20924 7012 20936
rect 6147 20887 6205 20893
rect 6472 20896 7012 20924
rect 6472 20868 6500 20896
rect 7006 20884 7012 20896
rect 7064 20884 7070 20936
rect 4246 20816 4252 20868
rect 4304 20856 4310 20868
rect 4678 20859 4736 20865
rect 4678 20856 4690 20859
rect 4304 20828 4690 20856
rect 4304 20816 4310 20828
rect 4678 20825 4690 20828
rect 4724 20825 4736 20859
rect 4678 20819 4736 20825
rect 6454 20816 6460 20868
rect 6512 20816 6518 20868
rect 6638 20816 6644 20868
rect 6696 20856 6702 20868
rect 7114 20856 7142 20964
rect 7469 20961 7481 20964
rect 7515 20961 7527 20995
rect 9692 21000 9720 21100
rect 9766 21088 9772 21140
rect 9824 21088 9830 21140
rect 9858 21088 9864 21140
rect 9916 21128 9922 21140
rect 14369 21131 14427 21137
rect 9916 21100 14228 21128
rect 9916 21088 9922 21100
rect 9784 21060 9812 21088
rect 10134 21060 10140 21072
rect 9784 21032 10140 21060
rect 10134 21020 10140 21032
rect 10192 21020 10198 21072
rect 10781 21063 10839 21069
rect 10781 21029 10793 21063
rect 10827 21060 10839 21063
rect 10870 21060 10876 21072
rect 10827 21032 10876 21060
rect 10827 21029 10839 21032
rect 10781 21023 10839 21029
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 9692 20992 9994 21000
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9692 20972 10057 20992
rect 9966 20964 10057 20972
rect 7469 20955 7527 20961
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 11333 20995 11391 21001
rect 11333 20961 11345 20995
rect 11379 20992 11391 20995
rect 11882 20992 11888 21004
rect 11379 20964 11888 20992
rect 11379 20961 11391 20964
rect 11333 20955 11391 20961
rect 11882 20952 11888 20964
rect 11940 20952 11946 21004
rect 7374 20884 7380 20936
rect 7432 20924 7438 20936
rect 7743 20927 7801 20933
rect 7743 20924 7755 20927
rect 7432 20896 7755 20924
rect 7432 20884 7438 20896
rect 7743 20893 7755 20896
rect 7789 20893 7801 20927
rect 9493 20927 9551 20933
rect 9493 20924 9505 20927
rect 7743 20887 7801 20893
rect 8680 20896 9505 20924
rect 8680 20868 8708 20896
rect 9493 20893 9505 20896
rect 9539 20893 9551 20927
rect 9493 20887 9551 20893
rect 6696 20828 7142 20856
rect 6696 20816 6702 20828
rect 8662 20816 8668 20868
rect 8720 20816 8726 20868
rect 9508 20856 9536 20887
rect 9674 20884 9680 20936
rect 9732 20884 9738 20936
rect 9769 20927 9827 20933
rect 9769 20893 9781 20927
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 9784 20856 9812 20887
rect 9858 20884 9864 20936
rect 9916 20884 9922 20936
rect 10137 20927 10195 20933
rect 10137 20924 10149 20927
rect 9968 20896 10149 20924
rect 9048 20828 9444 20856
rect 9508 20828 9812 20856
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 6917 20791 6975 20797
rect 6917 20788 6929 20791
rect 6788 20760 6929 20788
rect 6788 20748 6794 20760
rect 6917 20757 6929 20760
rect 6963 20757 6975 20791
rect 6917 20751 6975 20757
rect 7466 20748 7472 20800
rect 7524 20788 7530 20800
rect 9048 20788 9076 20828
rect 7524 20760 9076 20788
rect 9416 20788 9444 20828
rect 9968 20788 9996 20896
rect 10137 20893 10149 20896
rect 10183 20893 10195 20927
rect 10137 20887 10195 20893
rect 10318 20884 10324 20936
rect 10376 20884 10382 20936
rect 11054 20884 11060 20936
rect 11112 20884 11118 20936
rect 11238 20933 11244 20936
rect 11195 20927 11244 20933
rect 11195 20893 11207 20927
rect 11241 20893 11244 20927
rect 11195 20887 11244 20893
rect 11238 20884 11244 20887
rect 11296 20884 11302 20936
rect 11977 20927 12035 20933
rect 11977 20893 11989 20927
rect 12023 20924 12035 20927
rect 12345 20927 12403 20933
rect 12345 20924 12357 20927
rect 12023 20896 12357 20924
rect 12023 20893 12035 20896
rect 11977 20887 12035 20893
rect 12345 20893 12357 20896
rect 12391 20893 12403 20927
rect 12345 20887 12403 20893
rect 12434 20884 12440 20936
rect 12492 20884 12498 20936
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 14200 20933 14228 21100
rect 14369 21097 14381 21131
rect 14415 21128 14427 21131
rect 15102 21128 15108 21140
rect 14415 21100 15108 21128
rect 14415 21097 14427 21100
rect 14369 21091 14427 21097
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 12711 20927 12769 20933
rect 12711 20924 12723 20927
rect 12676 20896 12723 20924
rect 12676 20884 12682 20896
rect 12711 20893 12723 20896
rect 12757 20893 12769 20927
rect 12711 20887 12769 20893
rect 14185 20927 14243 20933
rect 14185 20893 14197 20927
rect 14231 20893 14243 20927
rect 14185 20887 14243 20893
rect 12406 20828 14228 20856
rect 9416 20760 9996 20788
rect 10045 20791 10103 20797
rect 7524 20748 7530 20760
rect 10045 20757 10057 20791
rect 10091 20788 10103 20791
rect 10870 20788 10876 20800
rect 10091 20760 10876 20788
rect 10091 20757 10103 20760
rect 10045 20751 10103 20757
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 11238 20748 11244 20800
rect 11296 20788 11302 20800
rect 11882 20788 11888 20800
rect 11296 20760 11888 20788
rect 11296 20748 11302 20760
rect 11882 20748 11888 20760
rect 11940 20748 11946 20800
rect 12161 20791 12219 20797
rect 12161 20757 12173 20791
rect 12207 20788 12219 20791
rect 12406 20788 12434 20828
rect 14200 20800 14228 20828
rect 12207 20760 12434 20788
rect 13449 20791 13507 20797
rect 12207 20757 12219 20760
rect 12161 20751 12219 20757
rect 13449 20757 13461 20791
rect 13495 20788 13507 20791
rect 13538 20788 13544 20800
rect 13495 20760 13544 20788
rect 13495 20757 13507 20760
rect 13449 20751 13507 20757
rect 13538 20748 13544 20760
rect 13596 20748 13602 20800
rect 14182 20748 14188 20800
rect 14240 20748 14246 20800
rect 1104 20698 14971 20720
rect 1104 20646 4376 20698
rect 4428 20646 4440 20698
rect 4492 20646 4504 20698
rect 4556 20646 4568 20698
rect 4620 20646 4632 20698
rect 4684 20646 7803 20698
rect 7855 20646 7867 20698
rect 7919 20646 7931 20698
rect 7983 20646 7995 20698
rect 8047 20646 8059 20698
rect 8111 20646 11230 20698
rect 11282 20646 11294 20698
rect 11346 20646 11358 20698
rect 11410 20646 11422 20698
rect 11474 20646 11486 20698
rect 11538 20646 14657 20698
rect 14709 20646 14721 20698
rect 14773 20646 14785 20698
rect 14837 20646 14849 20698
rect 14901 20646 14913 20698
rect 14965 20646 14971 20698
rect 1104 20624 14971 20646
rect 5537 20587 5595 20593
rect 5537 20553 5549 20587
rect 5583 20584 5595 20587
rect 6546 20584 6552 20596
rect 5583 20556 6552 20584
rect 5583 20553 5595 20556
rect 5537 20547 5595 20553
rect 6546 20544 6552 20556
rect 6604 20544 6610 20596
rect 7098 20544 7104 20596
rect 7156 20584 7162 20596
rect 7374 20584 7380 20596
rect 7156 20556 7380 20584
rect 7156 20544 7162 20556
rect 7374 20544 7380 20556
rect 7432 20544 7438 20596
rect 8113 20587 8171 20593
rect 8113 20553 8125 20587
rect 8159 20584 8171 20587
rect 8662 20584 8668 20596
rect 8159 20556 8668 20584
rect 8159 20553 8171 20556
rect 8113 20547 8171 20553
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 9858 20544 9864 20596
rect 9916 20584 9922 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 9916 20556 10609 20584
rect 9916 20544 9922 20556
rect 10597 20553 10609 20556
rect 10643 20553 10655 20587
rect 10597 20547 10655 20553
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20584 11759 20587
rect 13354 20584 13360 20596
rect 11747 20556 13360 20584
rect 11747 20553 11759 20556
rect 11701 20547 11759 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 14148 20556 14289 20584
rect 14148 20544 14154 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 6730 20516 6736 20528
rect 1688 20488 2774 20516
rect 750 20408 756 20460
rect 808 20448 814 20460
rect 1688 20457 1716 20488
rect 1489 20451 1547 20457
rect 1489 20448 1501 20451
rect 808 20420 1501 20448
rect 808 20408 814 20420
rect 1489 20417 1501 20420
rect 1535 20417 1547 20451
rect 1489 20411 1547 20417
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 2746 20312 2774 20488
rect 6564 20488 6736 20516
rect 4246 20408 4252 20460
rect 4304 20448 4310 20460
rect 5445 20451 5503 20457
rect 5445 20448 5457 20451
rect 4304 20420 5457 20448
rect 4304 20408 4310 20420
rect 5445 20417 5457 20420
rect 5491 20417 5503 20451
rect 5445 20411 5503 20417
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 6564 20457 6592 20488
rect 6730 20476 6736 20488
rect 6788 20476 6794 20528
rect 11514 20476 11520 20528
rect 11572 20516 11578 20528
rect 12434 20516 12440 20528
rect 11572 20488 12440 20516
rect 11572 20476 11578 20488
rect 12434 20476 12440 20488
rect 12492 20476 12498 20528
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20417 6607 20451
rect 7101 20451 7159 20457
rect 7101 20448 7113 20451
rect 6549 20411 6607 20417
rect 6656 20420 7113 20448
rect 5644 20380 5672 20408
rect 6656 20380 6684 20420
rect 7101 20417 7113 20420
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7375 20451 7433 20457
rect 7375 20448 7387 20451
rect 7340 20420 7387 20448
rect 7340 20408 7346 20420
rect 7375 20417 7387 20420
rect 7421 20417 7433 20451
rect 7375 20411 7433 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20448 10563 20451
rect 11057 20451 11115 20457
rect 10551 20420 10916 20448
rect 10551 20417 10563 20420
rect 10505 20411 10563 20417
rect 5644 20352 6684 20380
rect 6822 20340 6828 20392
rect 6880 20340 6886 20392
rect 7006 20312 7012 20324
rect 2746 20284 7012 20312
rect 7006 20272 7012 20284
rect 7064 20272 7070 20324
rect 10888 20321 10916 20420
rect 11057 20417 11069 20451
rect 11103 20448 11115 20451
rect 11238 20448 11244 20460
rect 11103 20420 11244 20448
rect 11103 20417 11115 20420
rect 11057 20411 11115 20417
rect 11238 20408 11244 20420
rect 11296 20408 11302 20460
rect 11885 20451 11943 20457
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 11900 20380 11928 20411
rect 12158 20408 12164 20460
rect 12216 20408 12222 20460
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 12308 20420 12664 20448
rect 12308 20408 12314 20420
rect 11974 20380 11980 20392
rect 11900 20352 11980 20380
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 12345 20383 12403 20389
rect 12345 20349 12357 20383
rect 12391 20380 12403 20383
rect 12434 20380 12440 20392
rect 12391 20352 12440 20380
rect 12391 20349 12403 20352
rect 12345 20343 12403 20349
rect 12434 20340 12440 20352
rect 12492 20340 12498 20392
rect 12529 20383 12587 20389
rect 12529 20349 12541 20383
rect 12575 20349 12587 20383
rect 12529 20343 12587 20349
rect 10873 20315 10931 20321
rect 10873 20281 10885 20315
rect 10919 20281 10931 20315
rect 10873 20275 10931 20281
rect 12066 20272 12072 20324
rect 12124 20312 12130 20324
rect 12544 20312 12572 20343
rect 12124 20284 12572 20312
rect 12124 20272 12130 20284
rect 6089 20247 6147 20253
rect 6089 20213 6101 20247
rect 6135 20244 6147 20247
rect 6641 20247 6699 20253
rect 6641 20244 6653 20247
rect 6135 20216 6653 20244
rect 6135 20213 6147 20216
rect 6089 20207 6147 20213
rect 6641 20213 6653 20216
rect 6687 20213 6699 20247
rect 6641 20207 6699 20213
rect 6733 20247 6791 20253
rect 6733 20213 6745 20247
rect 6779 20244 6791 20247
rect 7558 20244 7564 20256
rect 6779 20216 7564 20244
rect 6779 20213 6791 20216
rect 6733 20207 6791 20213
rect 7558 20204 7564 20216
rect 7616 20204 7622 20256
rect 11977 20247 12035 20253
rect 11977 20213 11989 20247
rect 12023 20244 12035 20247
rect 12434 20244 12440 20256
rect 12023 20216 12440 20244
rect 12023 20213 12035 20216
rect 11977 20207 12035 20213
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 12636 20244 12664 20420
rect 12710 20408 12716 20460
rect 12768 20408 12774 20460
rect 13262 20408 13268 20460
rect 13320 20408 13326 20460
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 14458 20408 14464 20460
rect 14516 20408 14522 20460
rect 12728 20380 12756 20408
rect 13354 20380 13360 20392
rect 13412 20389 13418 20392
rect 13412 20383 13440 20389
rect 12728 20352 13360 20380
rect 13354 20340 13360 20352
rect 13428 20349 13440 20383
rect 13412 20343 13440 20349
rect 13412 20340 13418 20343
rect 12710 20272 12716 20324
rect 12768 20312 12774 20324
rect 12989 20315 13047 20321
rect 12989 20312 13001 20315
rect 12768 20284 13001 20312
rect 12768 20272 12774 20284
rect 12989 20281 13001 20284
rect 13035 20281 13047 20315
rect 12989 20275 13047 20281
rect 14185 20247 14243 20253
rect 14185 20244 14197 20247
rect 12636 20216 14197 20244
rect 14185 20213 14197 20216
rect 14231 20213 14243 20247
rect 14185 20207 14243 20213
rect 1104 20154 14812 20176
rect 1104 20102 2663 20154
rect 2715 20102 2727 20154
rect 2779 20102 2791 20154
rect 2843 20102 2855 20154
rect 2907 20102 2919 20154
rect 2971 20102 6090 20154
rect 6142 20102 6154 20154
rect 6206 20102 6218 20154
rect 6270 20102 6282 20154
rect 6334 20102 6346 20154
rect 6398 20102 9517 20154
rect 9569 20102 9581 20154
rect 9633 20102 9645 20154
rect 9697 20102 9709 20154
rect 9761 20102 9773 20154
rect 9825 20102 12944 20154
rect 12996 20102 13008 20154
rect 13060 20102 13072 20154
rect 13124 20102 13136 20154
rect 13188 20102 13200 20154
rect 13252 20102 14812 20154
rect 1104 20080 14812 20102
rect 5994 20000 6000 20052
rect 6052 20000 6058 20052
rect 6362 20000 6368 20052
rect 6420 20000 6426 20052
rect 6733 20043 6791 20049
rect 6733 20009 6745 20043
rect 6779 20040 6791 20043
rect 6822 20040 6828 20052
rect 6779 20012 6828 20040
rect 6779 20009 6791 20012
rect 6733 20003 6791 20009
rect 6822 20000 6828 20012
rect 6880 20000 6886 20052
rect 7006 20000 7012 20052
rect 7064 20040 7070 20052
rect 7064 20012 8340 20040
rect 7064 20000 7070 20012
rect 6012 19972 6040 20000
rect 7101 19975 7159 19981
rect 7101 19972 7113 19975
rect 6012 19944 7113 19972
rect 7101 19941 7113 19944
rect 7147 19941 7159 19975
rect 7101 19935 7159 19941
rect 2746 19876 8248 19904
rect 750 19728 756 19780
rect 808 19768 814 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 808 19740 1501 19768
rect 808 19728 814 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 1489 19731 1547 19737
rect 1673 19771 1731 19777
rect 1673 19737 1685 19771
rect 1719 19768 1731 19771
rect 2746 19768 2774 19876
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 6086 19836 6092 19848
rect 5776 19808 6092 19836
rect 5776 19796 5782 19808
rect 6086 19796 6092 19808
rect 6144 19796 6150 19848
rect 6362 19796 6368 19848
rect 6420 19796 6426 19848
rect 6546 19845 6552 19848
rect 6541 19836 6552 19845
rect 6507 19808 6552 19836
rect 6541 19799 6552 19808
rect 6546 19796 6552 19799
rect 6604 19796 6610 19848
rect 6641 19839 6699 19845
rect 6641 19805 6653 19839
rect 6687 19836 6699 19839
rect 6730 19836 6736 19848
rect 6687 19808 6736 19836
rect 6687 19805 6699 19808
rect 6641 19799 6699 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19805 6883 19839
rect 6825 19799 6883 19805
rect 6380 19768 6408 19796
rect 6840 19768 6868 19799
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7285 19839 7343 19845
rect 7285 19836 7297 19839
rect 7156 19808 7297 19836
rect 7156 19796 7162 19808
rect 7285 19805 7297 19808
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 1719 19740 2774 19768
rect 3344 19740 6316 19768
rect 6380 19740 6868 19768
rect 8220 19768 8248 19876
rect 8312 19836 8340 20012
rect 9122 20000 9128 20052
rect 9180 20040 9186 20052
rect 9766 20040 9772 20052
rect 9180 20012 9772 20040
rect 9180 20000 9186 20012
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 11790 20040 11796 20052
rect 9968 20012 11796 20040
rect 9140 19972 9168 20000
rect 9048 19944 9168 19972
rect 9048 19913 9076 19944
rect 9033 19907 9091 19913
rect 9033 19873 9045 19907
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 9306 19836 9312 19848
rect 8312 19809 9312 19836
rect 8312 19808 9303 19809
rect 9291 19775 9303 19808
rect 9364 19796 9370 19848
rect 9337 19778 9352 19796
rect 9337 19775 9349 19778
rect 9291 19769 9349 19775
rect 8220 19740 9260 19768
rect 1719 19737 1731 19740
rect 1673 19731 1731 19737
rect 3344 19712 3372 19740
rect 3326 19660 3332 19712
rect 3384 19660 3390 19712
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 5994 19700 6000 19712
rect 5684 19672 6000 19700
rect 5684 19660 5690 19672
rect 5994 19660 6000 19672
rect 6052 19660 6058 19712
rect 6288 19700 6316 19740
rect 7098 19700 7104 19712
rect 6288 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 8938 19700 8944 19712
rect 8720 19672 8944 19700
rect 8720 19660 8726 19672
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9232 19700 9260 19740
rect 9968 19700 9996 20012
rect 11790 20000 11796 20012
rect 11848 20040 11854 20052
rect 11848 20012 12388 20040
rect 11848 20000 11854 20012
rect 11514 19864 11520 19916
rect 11572 19904 11578 19916
rect 11701 19907 11759 19913
rect 11701 19904 11713 19907
rect 11572 19876 11713 19904
rect 11572 19864 11578 19876
rect 11701 19873 11713 19876
rect 11747 19873 11759 19907
rect 11701 19867 11759 19873
rect 12360 19848 12388 20012
rect 12434 20000 12440 20052
rect 12492 20000 12498 20052
rect 12710 20000 12716 20052
rect 12768 20000 12774 20052
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 13780 20012 14381 20040
rect 13780 20000 13786 20012
rect 14369 20009 14381 20012
rect 14415 20009 14427 20043
rect 14369 20003 14427 20009
rect 15102 20000 15108 20052
rect 15160 20040 15166 20052
rect 15562 20040 15568 20052
rect 15160 20012 15568 20040
rect 15160 20000 15166 20012
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 12452 19972 12480 20000
rect 13814 19972 13820 19984
rect 12452 19944 13820 19972
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 13998 19932 14004 19984
rect 14056 19932 14062 19984
rect 13262 19864 13268 19916
rect 13320 19904 13326 19916
rect 14016 19904 14044 19932
rect 13320 19876 14044 19904
rect 13320 19864 13326 19876
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 11975 19839 12033 19845
rect 11975 19836 11987 19839
rect 11940 19808 11987 19836
rect 11940 19796 11946 19808
rect 11975 19805 11987 19808
rect 12021 19805 12033 19839
rect 11975 19799 12033 19805
rect 12342 19796 12348 19848
rect 12400 19796 12406 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13998 19836 14004 19848
rect 13403 19808 14004 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13998 19796 14004 19808
rect 14056 19796 14062 19848
rect 14182 19796 14188 19848
rect 14240 19796 14246 19848
rect 13725 19771 13783 19777
rect 13725 19737 13737 19771
rect 13771 19768 13783 19771
rect 14642 19768 14648 19780
rect 13771 19740 14648 19768
rect 13771 19737 13783 19740
rect 13725 19731 13783 19737
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 9232 19672 9996 19700
rect 10042 19660 10048 19712
rect 10100 19660 10106 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14458 19700 14464 19712
rect 14240 19672 14464 19700
rect 14240 19660 14246 19672
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 1104 19610 14971 19632
rect 1104 19558 4376 19610
rect 4428 19558 4440 19610
rect 4492 19558 4504 19610
rect 4556 19558 4568 19610
rect 4620 19558 4632 19610
rect 4684 19558 7803 19610
rect 7855 19558 7867 19610
rect 7919 19558 7931 19610
rect 7983 19558 7995 19610
rect 8047 19558 8059 19610
rect 8111 19558 11230 19610
rect 11282 19558 11294 19610
rect 11346 19558 11358 19610
rect 11410 19558 11422 19610
rect 11474 19558 11486 19610
rect 11538 19558 14657 19610
rect 14709 19558 14721 19610
rect 14773 19558 14785 19610
rect 14837 19558 14849 19610
rect 14901 19558 14913 19610
rect 14965 19558 14971 19610
rect 1104 19536 14971 19558
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 6914 19496 6920 19508
rect 5224 19468 6920 19496
rect 5224 19456 5230 19468
rect 6914 19456 6920 19468
rect 6972 19456 6978 19508
rect 9306 19456 9312 19508
rect 9364 19496 9370 19508
rect 11333 19499 11391 19505
rect 9364 19468 11190 19496
rect 9364 19456 9370 19468
rect 6932 19428 6960 19456
rect 6932 19400 7052 19428
rect 7024 19384 7052 19400
rect 7267 19393 7325 19399
rect 7267 19390 7279 19393
rect 7116 19384 7279 19390
rect 5626 19320 5632 19372
rect 5684 19320 5690 19372
rect 5718 19320 5724 19372
rect 5776 19320 5782 19372
rect 5821 19353 5879 19359
rect 4062 19252 4068 19304
rect 4120 19252 4126 19304
rect 5534 19252 5540 19304
rect 5592 19292 5598 19304
rect 5736 19292 5764 19320
rect 5821 19319 5833 19353
rect 5867 19350 5879 19353
rect 5867 19322 5948 19350
rect 5867 19319 5879 19322
rect 5821 19313 5879 19319
rect 5592 19264 5764 19292
rect 5592 19252 5598 19264
rect 4080 19224 4108 19252
rect 5920 19233 5948 19322
rect 6086 19320 6092 19372
rect 6144 19320 6150 19372
rect 7024 19362 7279 19384
rect 7024 19356 7144 19362
rect 7267 19359 7279 19362
rect 7313 19359 7325 19393
rect 8386 19388 8392 19440
rect 8444 19428 8450 19440
rect 8754 19428 8760 19440
rect 8444 19400 8760 19428
rect 8444 19388 8450 19400
rect 8754 19388 8760 19400
rect 8812 19388 8818 19440
rect 11162 19428 11190 19468
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 12158 19496 12164 19508
rect 11379 19468 12164 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 14001 19499 14059 19505
rect 14001 19465 14013 19499
rect 14047 19496 14059 19499
rect 14090 19496 14096 19508
rect 14047 19468 14096 19496
rect 14047 19465 14059 19468
rect 14001 19459 14059 19465
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14366 19456 14372 19508
rect 14424 19456 14430 19508
rect 11162 19400 11894 19428
rect 11866 19399 11894 19400
rect 11866 19393 11925 19399
rect 7267 19353 7325 19359
rect 8772 19360 8800 19388
rect 8849 19363 8907 19369
rect 8849 19360 8861 19363
rect 8772 19332 8861 19360
rect 8849 19329 8861 19332
rect 8895 19329 8907 19363
rect 8849 19323 8907 19329
rect 9122 19320 9128 19372
rect 9180 19360 9186 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9180 19332 9505 19360
rect 9180 19320 9186 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9493 19323 9551 19329
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9858 19360 9864 19372
rect 9723 19332 9864 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 11609 19363 11667 19369
rect 11609 19329 11621 19363
rect 11655 19360 11667 19363
rect 11866 19362 11879 19393
rect 11655 19332 11689 19360
rect 11867 19359 11879 19362
rect 11913 19359 11925 19393
rect 13630 19388 13636 19440
rect 13688 19428 13694 19440
rect 13688 19400 14228 19428
rect 13688 19388 13694 19400
rect 11867 19353 11925 19359
rect 11655 19329 11667 19332
rect 11609 19323 11667 19329
rect 6638 19252 6644 19304
rect 6696 19292 6702 19304
rect 6822 19292 6828 19304
rect 6696 19264 6828 19292
rect 6696 19252 6702 19264
rect 6822 19252 6828 19264
rect 6880 19292 6886 19304
rect 7009 19295 7067 19301
rect 7009 19292 7021 19295
rect 6880 19264 7021 19292
rect 6880 19252 6886 19264
rect 7009 19261 7021 19264
rect 7055 19261 7067 19295
rect 7009 19255 7067 19261
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 7800 19264 9996 19292
rect 7800 19252 7806 19264
rect 5905 19227 5963 19233
rect 4080 19196 5856 19224
rect 3418 19116 3424 19168
rect 3476 19156 3482 19168
rect 4246 19156 4252 19168
rect 3476 19128 4252 19156
rect 3476 19116 3482 19128
rect 4246 19116 4252 19128
rect 4304 19116 4310 19168
rect 5718 19116 5724 19168
rect 5776 19116 5782 19168
rect 5828 19156 5856 19196
rect 5905 19193 5917 19227
rect 5951 19193 5963 19227
rect 9674 19224 9680 19236
rect 5905 19187 5963 19193
rect 7944 19196 9680 19224
rect 7944 19156 7972 19196
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 5828 19128 7972 19156
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 8202 19156 8208 19168
rect 8067 19128 8208 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8665 19159 8723 19165
rect 8665 19125 8677 19159
rect 8711 19156 8723 19159
rect 9030 19156 9036 19168
rect 8711 19128 9036 19156
rect 8711 19125 8723 19128
rect 8665 19119 8723 19125
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9968 19156 9996 19264
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 10137 19295 10195 19301
rect 10137 19292 10149 19295
rect 10100 19264 10149 19292
rect 10100 19252 10106 19264
rect 10137 19261 10149 19264
rect 10183 19261 10195 19295
rect 10137 19255 10195 19261
rect 10410 19252 10416 19304
rect 10468 19252 10474 19304
rect 10502 19252 10508 19304
rect 10560 19301 10566 19304
rect 10560 19295 10588 19301
rect 10576 19261 10588 19295
rect 10560 19255 10588 19261
rect 10560 19252 10566 19255
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 10502 19156 10508 19168
rect 9968 19128 10508 19156
rect 10502 19116 10508 19128
rect 10560 19156 10566 19168
rect 11422 19156 11428 19168
rect 10560 19128 11428 19156
rect 10560 19116 10566 19128
rect 11422 19116 11428 19128
rect 11480 19156 11486 19168
rect 11624 19156 11652 19323
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 14200 19369 14228 19400
rect 13081 19363 13139 19369
rect 13081 19360 13093 19363
rect 12492 19332 13093 19360
rect 12492 19320 12498 19332
rect 13081 19329 13093 19332
rect 13127 19329 13139 19363
rect 13081 19323 13139 19329
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 13740 19292 13768 19323
rect 12400 19264 13768 19292
rect 12400 19252 12406 19264
rect 14458 19224 14464 19236
rect 13372 19196 14464 19224
rect 11480 19128 11652 19156
rect 11480 19116 11486 19128
rect 12618 19116 12624 19168
rect 12676 19116 12682 19168
rect 13372 19165 13400 19196
rect 14458 19184 14464 19196
rect 14516 19184 14522 19236
rect 13357 19159 13415 19165
rect 13357 19125 13369 19159
rect 13403 19125 13415 19159
rect 13357 19119 13415 19125
rect 1104 19066 14812 19088
rect 1104 19014 2663 19066
rect 2715 19014 2727 19066
rect 2779 19014 2791 19066
rect 2843 19014 2855 19066
rect 2907 19014 2919 19066
rect 2971 19014 6090 19066
rect 6142 19014 6154 19066
rect 6206 19014 6218 19066
rect 6270 19014 6282 19066
rect 6334 19014 6346 19066
rect 6398 19014 9517 19066
rect 9569 19014 9581 19066
rect 9633 19014 9645 19066
rect 9697 19014 9709 19066
rect 9761 19014 9773 19066
rect 9825 19014 12944 19066
rect 12996 19014 13008 19066
rect 13060 19014 13072 19066
rect 13124 19014 13136 19066
rect 13188 19014 13200 19066
rect 13252 19014 14812 19066
rect 1104 18992 14812 19014
rect 1578 18912 1584 18964
rect 1636 18912 1642 18964
rect 5718 18912 5724 18964
rect 5776 18912 5782 18964
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 7616 18924 10640 18952
rect 7616 18912 7622 18924
rect 5353 18887 5411 18893
rect 5353 18853 5365 18887
rect 5399 18884 5411 18887
rect 5626 18884 5632 18896
rect 5399 18856 5632 18884
rect 5399 18853 5411 18856
rect 5353 18847 5411 18853
rect 5626 18844 5632 18856
rect 5684 18844 5690 18896
rect 750 18708 756 18760
rect 808 18748 814 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 808 18720 1409 18748
rect 808 18708 814 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 4341 18751 4399 18757
rect 4341 18717 4353 18751
rect 4387 18717 4399 18751
rect 5644 18748 5672 18844
rect 5736 18816 5764 18912
rect 9033 18887 9091 18893
rect 9033 18853 9045 18887
rect 9079 18884 9091 18887
rect 10612 18884 10640 18924
rect 10686 18912 10692 18964
rect 10744 18952 10750 18964
rect 10965 18955 11023 18961
rect 10965 18952 10977 18955
rect 10744 18924 10977 18952
rect 10744 18912 10750 18924
rect 10965 18921 10977 18924
rect 11011 18921 11023 18955
rect 10965 18915 11023 18921
rect 11146 18912 11152 18964
rect 11204 18952 11210 18964
rect 11790 18952 11796 18964
rect 11204 18924 11796 18952
rect 11204 18912 11210 18924
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 12250 18952 12256 18964
rect 12207 18924 12256 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 12406 18924 14320 18952
rect 12406 18884 12434 18924
rect 9079 18856 9536 18884
rect 10612 18856 12434 18884
rect 9079 18853 9091 18856
rect 9033 18847 9091 18853
rect 9508 18825 9536 18856
rect 13630 18844 13636 18896
rect 13688 18884 13694 18896
rect 13725 18887 13783 18893
rect 13725 18884 13737 18887
rect 13688 18856 13737 18884
rect 13688 18844 13694 18856
rect 13725 18853 13737 18856
rect 13771 18853 13783 18887
rect 13725 18847 13783 18853
rect 13906 18844 13912 18896
rect 13964 18884 13970 18896
rect 13964 18856 14228 18884
rect 13964 18844 13970 18856
rect 5997 18819 6055 18825
rect 5997 18816 6009 18819
rect 5736 18788 6009 18816
rect 5997 18785 6009 18788
rect 6043 18785 6055 18819
rect 5997 18779 6055 18785
rect 7469 18819 7527 18825
rect 7469 18785 7481 18819
rect 7515 18785 7527 18819
rect 7469 18779 7527 18785
rect 9493 18819 9551 18825
rect 9493 18785 9505 18819
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 5721 18751 5779 18757
rect 5721 18748 5733 18751
rect 4341 18711 4399 18717
rect 4599 18721 4657 18727
rect 4356 18612 4384 18711
rect 4599 18687 4611 18721
rect 4645 18718 4657 18721
rect 5644 18720 5733 18748
rect 4645 18687 4660 18718
rect 5721 18717 5733 18720
rect 5767 18717 5779 18751
rect 5721 18711 5779 18717
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 5902 18720 6101 18748
rect 4599 18681 4660 18687
rect 4632 18680 4660 18681
rect 4798 18680 4804 18692
rect 4632 18652 4804 18680
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 5902 18680 5930 18720
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6347 18751 6405 18757
rect 6347 18748 6359 18751
rect 6089 18711 6147 18717
rect 6288 18720 6359 18748
rect 6178 18680 6184 18692
rect 5644 18652 6184 18680
rect 5644 18624 5672 18652
rect 6178 18640 6184 18652
rect 6236 18640 6242 18692
rect 5626 18612 5632 18624
rect 4356 18584 5632 18612
rect 5626 18572 5632 18584
rect 5684 18572 5690 18624
rect 5994 18572 6000 18624
rect 6052 18572 6058 18624
rect 6086 18572 6092 18624
rect 6144 18612 6150 18624
rect 6288 18612 6316 18720
rect 6347 18717 6359 18720
rect 6393 18717 6405 18751
rect 6347 18711 6405 18717
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 7374 18748 7380 18760
rect 6880 18720 7380 18748
rect 6880 18708 6886 18720
rect 7374 18708 7380 18720
rect 7432 18748 7438 18760
rect 7484 18748 7512 18779
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 9953 18819 10011 18825
rect 9953 18816 9965 18819
rect 9916 18788 9965 18816
rect 9916 18776 9922 18788
rect 9953 18785 9965 18788
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 11422 18776 11428 18828
rect 11480 18816 11486 18828
rect 12345 18819 12403 18825
rect 12345 18816 12357 18819
rect 11480 18788 12357 18816
rect 11480 18776 11486 18788
rect 12345 18785 12357 18788
rect 12391 18785 12403 18819
rect 12345 18779 12403 18785
rect 7432 18720 7512 18748
rect 7432 18708 7438 18720
rect 7650 18708 7656 18760
rect 7708 18748 7714 18760
rect 7743 18751 7801 18757
rect 7743 18748 7755 18751
rect 7708 18720 7755 18748
rect 7708 18708 7714 18720
rect 7743 18717 7755 18720
rect 7789 18717 7801 18751
rect 7743 18711 7801 18717
rect 8941 18751 8999 18757
rect 8941 18717 8953 18751
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 8956 18680 8984 18711
rect 9030 18708 9036 18760
rect 9088 18748 9094 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 9088 18720 9137 18748
rect 9088 18708 9094 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9232 18680 9260 18711
rect 9306 18708 9312 18760
rect 9364 18708 9370 18760
rect 10134 18708 10140 18760
rect 10192 18748 10198 18760
rect 10227 18751 10285 18757
rect 10227 18748 10239 18751
rect 10192 18720 10239 18748
rect 10192 18708 10198 18720
rect 10227 18717 10239 18720
rect 10273 18717 10285 18751
rect 11517 18751 11575 18757
rect 10227 18711 10285 18717
rect 10704 18720 11100 18748
rect 7116 18652 9260 18680
rect 7116 18621 7144 18652
rect 6144 18584 6316 18612
rect 7101 18615 7159 18621
rect 6144 18572 6150 18584
rect 7101 18581 7113 18615
rect 7147 18581 7159 18615
rect 7101 18575 7159 18581
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 7742 18612 7748 18624
rect 7432 18584 7748 18612
rect 7432 18572 7438 18584
rect 7742 18572 7748 18584
rect 7800 18572 7806 18624
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 8938 18612 8944 18624
rect 8527 18584 8944 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9493 18615 9551 18621
rect 9493 18581 9505 18615
rect 9539 18612 9551 18615
rect 10042 18612 10048 18624
rect 9539 18584 10048 18612
rect 9539 18581 9551 18584
rect 9493 18575 9551 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10594 18572 10600 18624
rect 10652 18612 10658 18624
rect 10704 18612 10732 18720
rect 11072 18680 11100 18720
rect 11517 18717 11529 18751
rect 11563 18748 11575 18751
rect 12066 18748 12072 18760
rect 11563 18720 12072 18748
rect 11563 18717 11575 18720
rect 11517 18711 11575 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12587 18751 12645 18757
rect 12587 18717 12599 18751
rect 12633 18748 12645 18751
rect 12710 18748 12716 18760
rect 12633 18720 12716 18748
rect 12633 18717 12645 18720
rect 12587 18711 12645 18717
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 13906 18708 13912 18760
rect 13964 18708 13970 18760
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 11072 18652 11897 18680
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 14200 18680 14228 18856
rect 14292 18757 14320 18924
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18717 14335 18751
rect 14277 18711 14335 18717
rect 14458 18680 14464 18692
rect 14200 18652 14464 18680
rect 11885 18643 11943 18649
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 15102 18640 15108 18692
rect 15160 18640 15166 18692
rect 10652 18584 10732 18612
rect 10652 18572 10658 18584
rect 10778 18572 10784 18624
rect 10836 18612 10842 18624
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 10836 18584 11345 18612
rect 10836 18572 10842 18584
rect 11333 18581 11345 18584
rect 11379 18581 11391 18615
rect 11333 18575 11391 18581
rect 13262 18572 13268 18624
rect 13320 18612 13326 18624
rect 13357 18615 13415 18621
rect 13357 18612 13369 18615
rect 13320 18584 13369 18612
rect 13320 18572 13326 18584
rect 13357 18581 13369 18584
rect 13403 18581 13415 18615
rect 13357 18575 13415 18581
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 1104 18522 14971 18544
rect 1104 18470 4376 18522
rect 4428 18470 4440 18522
rect 4492 18470 4504 18522
rect 4556 18470 4568 18522
rect 4620 18470 4632 18522
rect 4684 18470 7803 18522
rect 7855 18470 7867 18522
rect 7919 18470 7931 18522
rect 7983 18470 7995 18522
rect 8047 18470 8059 18522
rect 8111 18470 11230 18522
rect 11282 18470 11294 18522
rect 11346 18470 11358 18522
rect 11410 18470 11422 18522
rect 11474 18470 11486 18522
rect 11538 18470 14657 18522
rect 14709 18470 14721 18522
rect 14773 18470 14785 18522
rect 14837 18470 14849 18522
rect 14901 18470 14913 18522
rect 14965 18470 14971 18522
rect 1104 18448 14971 18470
rect 5534 18368 5540 18420
rect 5592 18368 5598 18420
rect 5810 18368 5816 18420
rect 5868 18368 5874 18420
rect 5994 18368 6000 18420
rect 6052 18368 6058 18420
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 8754 18408 8760 18420
rect 6880 18380 8760 18408
rect 6880 18368 6886 18380
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 10321 18411 10379 18417
rect 10321 18408 10333 18411
rect 9364 18380 10333 18408
rect 9364 18368 9370 18380
rect 10321 18377 10333 18380
rect 10367 18377 10379 18411
rect 10321 18371 10379 18377
rect 11333 18411 11391 18417
rect 11333 18377 11345 18411
rect 11379 18377 11391 18411
rect 13354 18408 13360 18420
rect 11333 18371 11391 18377
rect 12084 18380 13360 18408
rect 6012 18340 6040 18368
rect 6012 18312 6592 18340
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 4154 18232 4160 18284
rect 4212 18232 4218 18284
rect 4430 18281 4436 18284
rect 4424 18272 4436 18281
rect 4391 18244 4436 18272
rect 4424 18235 4436 18244
rect 4430 18232 4436 18235
rect 4488 18232 4494 18284
rect 6564 18281 6592 18312
rect 6730 18300 6736 18352
rect 6788 18340 6794 18352
rect 7650 18340 7656 18352
rect 6788 18312 7656 18340
rect 6788 18300 6794 18312
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 10686 18340 10692 18352
rect 9600 18312 10692 18340
rect 5721 18275 5779 18281
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6181 18275 6239 18281
rect 5767 18244 6040 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 566 18164 572 18216
rect 624 18204 630 18216
rect 4172 18204 4200 18232
rect 624 18176 4200 18204
rect 624 18164 630 18176
rect 1673 18139 1731 18145
rect 1673 18105 1685 18139
rect 1719 18136 1731 18139
rect 2498 18136 2504 18148
rect 1719 18108 2504 18136
rect 1719 18105 1731 18108
rect 1673 18099 1731 18105
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 6012 18145 6040 18244
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6181 18235 6239 18241
rect 6549 18275 6607 18281
rect 6549 18241 6561 18275
rect 6595 18241 6607 18275
rect 6549 18235 6607 18241
rect 6196 18204 6224 18235
rect 8754 18232 8760 18284
rect 8812 18232 8818 18284
rect 9030 18232 9036 18284
rect 9088 18232 9094 18284
rect 6196 18176 7052 18204
rect 7024 18148 7052 18176
rect 7374 18164 7380 18216
rect 7432 18204 7438 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7432 18176 7849 18204
rect 7432 18164 7438 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7837 18167 7895 18173
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18173 8079 18207
rect 8021 18167 8079 18173
rect 5997 18139 6055 18145
rect 5997 18105 6009 18139
rect 6043 18105 6055 18139
rect 5997 18099 6055 18105
rect 7006 18096 7012 18148
rect 7064 18136 7070 18148
rect 8036 18136 8064 18167
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8260 18176 8493 18204
rect 8260 18164 8266 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 8895 18207 8953 18213
rect 8895 18173 8907 18207
rect 8941 18204 8953 18207
rect 9600 18204 9628 18312
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 10778 18300 10784 18352
rect 10836 18300 10842 18352
rect 10870 18300 10876 18352
rect 10928 18300 10934 18352
rect 11348 18340 11376 18371
rect 12084 18340 12112 18380
rect 13354 18368 13360 18380
rect 13412 18368 13418 18420
rect 13633 18411 13691 18417
rect 13633 18377 13645 18411
rect 13679 18408 13691 18411
rect 14366 18408 14372 18420
rect 13679 18380 14372 18408
rect 13679 18377 13691 18380
rect 13633 18371 13691 18377
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 15120 18408 15148 18640
rect 14700 18380 15148 18408
rect 14700 18368 14706 18380
rect 15286 18368 15292 18420
rect 15344 18368 15350 18420
rect 11348 18312 12112 18340
rect 12158 18300 12164 18352
rect 12216 18340 12222 18352
rect 13446 18340 13452 18352
rect 12216 18312 13452 18340
rect 12216 18300 12222 18312
rect 13446 18300 13452 18312
rect 13504 18300 13510 18352
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 13872 18312 14105 18340
rect 13872 18300 13878 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 14093 18303 14151 18309
rect 14461 18343 14519 18349
rect 14461 18309 14473 18343
rect 14507 18309 14519 18343
rect 14461 18303 14519 18309
rect 9674 18232 9680 18284
rect 9732 18232 9738 18284
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18272 10287 18275
rect 10796 18272 10824 18300
rect 10275 18244 10824 18272
rect 10888 18272 10916 18300
rect 11057 18275 11115 18281
rect 11057 18272 11069 18275
rect 10888 18244 11069 18272
rect 10275 18241 10287 18244
rect 10229 18235 10287 18241
rect 11057 18241 11069 18244
rect 11103 18241 11115 18275
rect 11057 18235 11115 18241
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11238 18272 11244 18284
rect 11195 18244 11244 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11238 18232 11244 18244
rect 11296 18232 11302 18284
rect 11790 18272 11796 18284
rect 11751 18244 11796 18272
rect 11790 18232 11796 18244
rect 11848 18232 11854 18284
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18272 13415 18275
rect 14366 18272 14372 18284
rect 13403 18244 14372 18272
rect 13403 18241 13415 18244
rect 13357 18235 13415 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14476 18272 14504 18303
rect 15304 18272 15332 18368
rect 14476 18244 15332 18272
rect 8941 18176 9628 18204
rect 8941 18173 8953 18176
rect 8895 18167 8953 18173
rect 10778 18164 10784 18216
rect 10836 18204 10842 18216
rect 11517 18207 11575 18213
rect 11517 18204 11529 18207
rect 10836 18176 11529 18204
rect 10836 18164 10842 18176
rect 11517 18173 11529 18176
rect 11563 18173 11575 18207
rect 11517 18167 11575 18173
rect 10962 18136 10968 18148
rect 7064 18108 8064 18136
rect 10520 18108 10968 18136
rect 7064 18096 7070 18108
rect 10520 18080 10548 18108
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 6365 18071 6423 18077
rect 6365 18037 6377 18071
rect 6411 18068 6423 18071
rect 8202 18068 8208 18080
rect 6411 18040 8208 18068
rect 6411 18037 6423 18040
rect 6365 18031 6423 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 10502 18028 10508 18080
rect 10560 18028 10566 18080
rect 10873 18071 10931 18077
rect 10873 18037 10885 18071
rect 10919 18068 10931 18071
rect 12434 18068 12440 18080
rect 10919 18040 12440 18068
rect 10919 18037 10931 18040
rect 10873 18031 10931 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12529 18071 12587 18077
rect 12529 18037 12541 18071
rect 12575 18068 12587 18071
rect 12710 18068 12716 18080
rect 12575 18040 12716 18068
rect 12575 18037 12587 18040
rect 12529 18031 12587 18037
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 12989 18071 13047 18077
rect 12989 18068 13001 18071
rect 12860 18040 13001 18068
rect 12860 18028 12866 18040
rect 12989 18037 13001 18040
rect 13035 18037 13047 18071
rect 12989 18031 13047 18037
rect 13446 18028 13452 18080
rect 13504 18068 13510 18080
rect 14182 18068 14188 18080
rect 13504 18040 14188 18068
rect 13504 18028 13510 18040
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 1104 17978 14812 18000
rect 1104 17926 2663 17978
rect 2715 17926 2727 17978
rect 2779 17926 2791 17978
rect 2843 17926 2855 17978
rect 2907 17926 2919 17978
rect 2971 17926 6090 17978
rect 6142 17926 6154 17978
rect 6206 17926 6218 17978
rect 6270 17926 6282 17978
rect 6334 17926 6346 17978
rect 6398 17926 9517 17978
rect 9569 17926 9581 17978
rect 9633 17926 9645 17978
rect 9697 17926 9709 17978
rect 9761 17926 9773 17978
rect 9825 17926 12944 17978
rect 12996 17926 13008 17978
rect 13060 17926 13072 17978
rect 13124 17926 13136 17978
rect 13188 17926 13200 17978
rect 13252 17926 14812 17978
rect 1104 17904 14812 17926
rect 10229 17867 10287 17873
rect 10229 17833 10241 17867
rect 10275 17864 10287 17867
rect 10594 17864 10600 17876
rect 10275 17836 10600 17864
rect 10275 17833 10287 17836
rect 10229 17827 10287 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 10686 17824 10692 17876
rect 10744 17824 10750 17876
rect 12526 17824 12532 17876
rect 12584 17824 12590 17876
rect 13265 17867 13323 17873
rect 13265 17833 13277 17867
rect 13311 17864 13323 17867
rect 13354 17864 13360 17876
rect 13311 17836 13360 17864
rect 13311 17833 13323 17836
rect 13265 17827 13323 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 14369 17867 14427 17873
rect 14369 17833 14381 17867
rect 14415 17864 14427 17867
rect 15102 17864 15108 17876
rect 14415 17836 15108 17864
rect 14415 17833 14427 17836
rect 14369 17827 14427 17833
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 15562 17824 15568 17876
rect 15620 17824 15626 17876
rect 7193 17799 7251 17805
rect 7193 17796 7205 17799
rect 7024 17768 7205 17796
rect 4890 17688 4896 17740
rect 4948 17728 4954 17740
rect 5442 17728 5448 17740
rect 4948 17700 5448 17728
rect 4948 17688 4954 17700
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 6178 17688 6184 17740
rect 6236 17688 6242 17740
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 7024 17660 7052 17768
rect 7193 17765 7205 17768
rect 7239 17765 7251 17799
rect 13722 17796 13728 17808
rect 7193 17759 7251 17765
rect 12544 17768 13728 17796
rect 9766 17728 9772 17740
rect 9324 17700 9772 17728
rect 9324 17672 9352 17700
rect 9766 17688 9772 17700
rect 9824 17728 9830 17740
rect 10778 17728 10784 17740
rect 9824 17700 10784 17728
rect 9824 17688 9830 17700
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 12434 17728 12440 17740
rect 12124 17700 12440 17728
rect 12124 17688 12130 17700
rect 12434 17688 12440 17700
rect 12492 17688 12498 17740
rect 4028 17632 7052 17660
rect 4028 17620 4034 17632
rect 9306 17620 9312 17672
rect 9364 17620 9370 17672
rect 9858 17620 9864 17672
rect 9916 17660 9922 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 9916 17632 10425 17660
rect 9916 17620 9922 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10505 17663 10563 17669
rect 10505 17629 10517 17663
rect 10551 17629 10563 17663
rect 11054 17660 11060 17672
rect 11015 17632 11060 17660
rect 10505 17623 10563 17629
rect 4154 17552 4160 17604
rect 4212 17592 4218 17604
rect 4430 17592 4436 17604
rect 4212 17564 4436 17592
rect 4212 17552 4218 17564
rect 4430 17552 4436 17564
rect 4488 17592 4494 17604
rect 5077 17595 5135 17601
rect 5077 17592 5089 17595
rect 4488 17564 5089 17592
rect 4488 17552 4494 17564
rect 5077 17561 5089 17564
rect 5123 17561 5135 17595
rect 5077 17555 5135 17561
rect 5902 17552 5908 17604
rect 5960 17552 5966 17604
rect 6181 17595 6239 17601
rect 6181 17561 6193 17595
rect 6227 17561 6239 17595
rect 6181 17555 6239 17561
rect 6273 17595 6331 17601
rect 6273 17561 6285 17595
rect 6319 17592 6331 17595
rect 6546 17592 6552 17604
rect 6319 17564 6552 17592
rect 6319 17561 6331 17564
rect 6273 17555 6331 17561
rect 5169 17527 5227 17533
rect 5169 17493 5181 17527
rect 5215 17524 5227 17527
rect 6196 17524 6224 17555
rect 6546 17552 6552 17564
rect 6604 17552 6610 17604
rect 6638 17552 6644 17604
rect 6696 17552 6702 17604
rect 6822 17552 6828 17604
rect 6880 17552 6886 17604
rect 10520 17592 10548 17623
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12544 17660 12572 17768
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 13817 17799 13875 17805
rect 13817 17765 13829 17799
rect 13863 17796 13875 17799
rect 15580 17796 15608 17824
rect 13863 17768 15608 17796
rect 13863 17765 13875 17768
rect 13817 17759 13875 17765
rect 14274 17728 14280 17740
rect 12636 17700 14280 17728
rect 12636 17669 12664 17700
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 12391 17632 12572 17660
rect 12621 17663 12679 17669
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12621 17629 12633 17663
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12802 17620 12808 17672
rect 12860 17660 12866 17672
rect 12989 17663 13047 17669
rect 12989 17660 13001 17663
rect 12860 17632 13001 17660
rect 12860 17620 12866 17632
rect 12989 17629 13001 17632
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 13078 17620 13084 17672
rect 13136 17660 13142 17672
rect 13136 17632 13676 17660
rect 13136 17620 13142 17632
rect 11422 17592 11428 17604
rect 10520 17564 11428 17592
rect 11422 17552 11428 17564
rect 11480 17552 11486 17604
rect 11882 17592 11888 17604
rect 11716 17564 11888 17592
rect 6840 17524 6868 17552
rect 5215 17496 6868 17524
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 7006 17484 7012 17536
rect 7064 17484 7070 17536
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 11054 17524 11060 17536
rect 9088 17496 11060 17524
rect 9088 17484 9094 17496
rect 11054 17484 11060 17496
rect 11112 17524 11118 17536
rect 11716 17524 11744 17564
rect 11882 17552 11888 17564
rect 11940 17552 11946 17604
rect 12066 17552 12072 17604
rect 12124 17592 12130 17604
rect 13541 17595 13599 17601
rect 13541 17592 13553 17595
rect 12124 17564 13553 17592
rect 12124 17552 12130 17564
rect 13541 17561 13553 17564
rect 13587 17561 13599 17595
rect 13648 17592 13676 17632
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 14148 17632 14197 17660
rect 14148 17620 14154 17632
rect 14185 17629 14197 17632
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 14642 17592 14648 17604
rect 13648 17564 14648 17592
rect 13541 17555 13599 17561
rect 14642 17552 14648 17564
rect 14700 17552 14706 17604
rect 11112 17496 11744 17524
rect 11793 17527 11851 17533
rect 11112 17484 11118 17496
rect 11793 17493 11805 17527
rect 11839 17524 11851 17527
rect 12158 17524 12164 17536
rect 11839 17496 12164 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12805 17527 12863 17533
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 15856 17524 15884 17620
rect 12851 17496 15884 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 1104 17434 14971 17456
rect 1104 17382 4376 17434
rect 4428 17382 4440 17434
rect 4492 17382 4504 17434
rect 4556 17382 4568 17434
rect 4620 17382 4632 17434
rect 4684 17382 7803 17434
rect 7855 17382 7867 17434
rect 7919 17382 7931 17434
rect 7983 17382 7995 17434
rect 8047 17382 8059 17434
rect 8111 17382 11230 17434
rect 11282 17382 11294 17434
rect 11346 17382 11358 17434
rect 11410 17382 11422 17434
rect 11474 17382 11486 17434
rect 11538 17382 14657 17434
rect 14709 17382 14721 17434
rect 14773 17382 14785 17434
rect 14837 17382 14849 17434
rect 14901 17382 14913 17434
rect 14965 17382 14971 17434
rect 1104 17360 14971 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1627 17292 5178 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 750 17144 756 17196
rect 808 17184 814 17196
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 808 17156 1501 17184
rect 808 17144 814 17156
rect 1489 17153 1501 17156
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 4890 17144 4896 17196
rect 4948 17144 4954 17196
rect 5150 17193 5178 17292
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 7558 17320 7564 17332
rect 5960 17292 7564 17320
rect 5960 17280 5966 17292
rect 7558 17280 7564 17292
rect 7616 17320 7622 17332
rect 7742 17320 7748 17332
rect 7616 17292 7748 17320
rect 7616 17280 7622 17292
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8720 17292 11744 17320
rect 8720 17280 8726 17292
rect 5150 17187 5225 17193
rect 5150 17156 5179 17187
rect 5167 17153 5179 17156
rect 5213 17184 5225 17187
rect 5258 17184 5264 17196
rect 5213 17156 5264 17184
rect 5213 17153 5225 17156
rect 5167 17147 5225 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 6457 17187 6515 17193
rect 6457 17184 6469 17187
rect 5644 17156 6469 17184
rect 5644 17128 5672 17156
rect 6457 17153 6469 17156
rect 6503 17153 6515 17187
rect 6457 17147 6515 17153
rect 6731 17187 6789 17193
rect 6731 17153 6743 17187
rect 6777 17184 6789 17187
rect 9030 17184 9036 17196
rect 6777 17156 9036 17184
rect 6777 17153 6789 17156
rect 6731 17147 6789 17153
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 9214 17144 9220 17196
rect 9272 17184 9278 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9272 17156 9413 17184
rect 9272 17144 9278 17156
rect 9401 17153 9413 17156
rect 9447 17153 9459 17187
rect 11716 17184 11744 17292
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 13357 17323 13415 17329
rect 13357 17320 13369 17323
rect 12032 17292 13369 17320
rect 12032 17280 12038 17292
rect 13357 17289 13369 17292
rect 13403 17289 13415 17323
rect 13357 17283 13415 17289
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 15194 17320 15200 17332
rect 14231 17292 15200 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 15286 17212 15292 17264
rect 15344 17252 15350 17264
rect 15562 17252 15568 17264
rect 15344 17224 15568 17252
rect 15344 17212 15350 17224
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 11716 17156 11928 17184
rect 9401 17147 9459 17153
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 6178 17076 6184 17128
rect 6236 17076 6242 17128
rect 8846 17076 8852 17128
rect 8904 17116 8910 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 8904 17088 9597 17116
rect 8904 17076 8910 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17048 5963 17051
rect 6196 17048 6224 17076
rect 8294 17048 8300 17060
rect 5951 17020 6224 17048
rect 7392 17020 8300 17048
rect 5951 17017 5963 17020
rect 5905 17011 5963 17017
rect 4890 16940 4896 16992
rect 4948 16980 4954 16992
rect 7392 16980 7420 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 4948 16952 7420 16980
rect 7469 16983 7527 16989
rect 4948 16940 4954 16952
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 7558 16980 7564 16992
rect 7515 16952 7564 16980
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 9600 16980 9628 17079
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 10502 17125 10508 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10192 17088 10333 17116
rect 10192 17076 10198 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 10321 17079 10379 17085
rect 10459 17119 10508 17125
rect 10459 17085 10471 17119
rect 10505 17085 10508 17119
rect 10459 17079 10508 17085
rect 10502 17076 10508 17079
rect 10560 17076 10566 17128
rect 10594 17076 10600 17128
rect 10652 17076 10658 17128
rect 11517 17119 11575 17125
rect 11517 17085 11529 17119
rect 11563 17116 11575 17119
rect 11606 17116 11612 17128
rect 11563 17088 11612 17116
rect 11563 17085 11575 17088
rect 11517 17079 11575 17085
rect 11606 17076 11612 17088
rect 11664 17076 11670 17128
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 10042 17008 10048 17060
rect 10100 17008 10106 17060
rect 10778 16980 10784 16992
rect 9600 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11238 16940 11244 16992
rect 11296 16940 11302 16992
rect 11716 16980 11744 17079
rect 11900 17048 11928 17156
rect 12434 17144 12440 17196
rect 12492 17144 12498 17196
rect 12710 17144 12716 17196
rect 12768 17144 12774 17196
rect 13538 17144 13544 17196
rect 13596 17144 13602 17196
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 13909 17187 13967 17193
rect 13909 17184 13921 17187
rect 13688 17156 13921 17184
rect 13688 17144 13694 17156
rect 13909 17153 13921 17156
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 12158 17076 12164 17128
rect 12216 17076 12222 17128
rect 12526 17076 12532 17128
rect 12584 17125 12590 17128
rect 12584 17119 12633 17125
rect 12584 17085 12587 17119
rect 12621 17116 12633 17119
rect 13078 17116 13084 17128
rect 12621 17088 13084 17116
rect 12621 17085 12633 17088
rect 12584 17079 12633 17085
rect 12584 17076 12590 17079
rect 13078 17076 13084 17088
rect 13136 17076 13142 17128
rect 11900 17020 12296 17048
rect 11882 16980 11888 16992
rect 11716 16952 11888 16980
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12268 16980 12296 17020
rect 13096 17020 13676 17048
rect 13096 16980 13124 17020
rect 13648 16989 13676 17020
rect 12268 16952 13124 16980
rect 13633 16983 13691 16989
rect 13633 16949 13645 16983
rect 13679 16949 13691 16983
rect 13633 16943 13691 16949
rect 1104 16890 14812 16912
rect 1104 16838 2663 16890
rect 2715 16838 2727 16890
rect 2779 16838 2791 16890
rect 2843 16838 2855 16890
rect 2907 16838 2919 16890
rect 2971 16838 6090 16890
rect 6142 16838 6154 16890
rect 6206 16838 6218 16890
rect 6270 16838 6282 16890
rect 6334 16838 6346 16890
rect 6398 16838 9517 16890
rect 9569 16838 9581 16890
rect 9633 16838 9645 16890
rect 9697 16838 9709 16890
rect 9761 16838 9773 16890
rect 9825 16838 12944 16890
rect 12996 16838 13008 16890
rect 13060 16838 13072 16890
rect 13124 16838 13136 16890
rect 13188 16838 13200 16890
rect 13252 16838 14812 16890
rect 1104 16816 14812 16838
rect 4890 16776 4896 16788
rect 1688 16748 4896 16776
rect 1688 16717 1716 16748
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 6546 16736 6552 16788
rect 6604 16736 6610 16788
rect 8294 16736 8300 16788
rect 8352 16776 8358 16788
rect 9674 16776 9680 16788
rect 8352 16748 9680 16776
rect 8352 16736 8358 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10413 16779 10471 16785
rect 10413 16745 10425 16779
rect 10459 16776 10471 16779
rect 10594 16776 10600 16788
rect 10459 16748 10600 16776
rect 10459 16745 10471 16748
rect 10413 16739 10471 16745
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 11793 16779 11851 16785
rect 11793 16745 11805 16779
rect 11839 16776 11851 16779
rect 12066 16776 12072 16788
rect 11839 16748 12072 16776
rect 11839 16745 11851 16748
rect 11793 16739 11851 16745
rect 12066 16736 12072 16748
rect 12124 16736 12130 16788
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 14369 16779 14427 16785
rect 14369 16776 14381 16779
rect 12768 16748 14381 16776
rect 12768 16736 12774 16748
rect 14369 16745 14381 16748
rect 14415 16745 14427 16779
rect 14369 16739 14427 16745
rect 1673 16711 1731 16717
rect 1673 16677 1685 16711
rect 1719 16677 1731 16711
rect 1673 16671 1731 16677
rect 8113 16711 8171 16717
rect 8113 16677 8125 16711
rect 8159 16708 8171 16711
rect 8662 16708 8668 16720
rect 8159 16680 8668 16708
rect 8159 16677 8171 16680
rect 8113 16671 8171 16677
rect 8662 16668 8668 16680
rect 8720 16668 8726 16720
rect 13909 16711 13967 16717
rect 13909 16677 13921 16711
rect 13955 16708 13967 16711
rect 14182 16708 14188 16720
rect 13955 16680 14188 16708
rect 13955 16677 13967 16680
rect 13909 16671 13967 16677
rect 14182 16668 14188 16680
rect 14240 16668 14246 16720
rect 5442 16600 5448 16652
rect 5500 16640 5506 16652
rect 5537 16643 5595 16649
rect 5537 16640 5549 16643
rect 5500 16612 5549 16640
rect 5500 16600 5506 16612
rect 5537 16609 5549 16612
rect 5583 16609 5595 16643
rect 7101 16643 7159 16649
rect 7101 16640 7113 16643
rect 5537 16603 5595 16609
rect 6196 16612 7113 16640
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 5166 16572 5172 16584
rect 2556 16544 5172 16572
rect 2556 16532 2562 16544
rect 5166 16532 5172 16544
rect 5224 16572 5230 16584
rect 5779 16575 5837 16581
rect 5779 16572 5791 16575
rect 5224 16544 5791 16572
rect 5224 16532 5230 16544
rect 5779 16541 5791 16544
rect 5825 16541 5837 16575
rect 6196 16572 6224 16612
rect 7101 16609 7113 16612
rect 7147 16609 7159 16643
rect 7101 16603 7159 16609
rect 11882 16600 11888 16652
rect 11940 16640 11946 16652
rect 12253 16643 12311 16649
rect 12253 16640 12265 16643
rect 11940 16612 12265 16640
rect 11940 16600 11946 16612
rect 12253 16609 12265 16612
rect 12299 16609 12311 16643
rect 12253 16603 12311 16609
rect 12618 16600 12624 16652
rect 12676 16640 12682 16652
rect 12713 16643 12771 16649
rect 12713 16640 12725 16643
rect 12676 16612 12725 16640
rect 12676 16600 12682 16612
rect 12713 16609 12725 16612
rect 12759 16609 12771 16643
rect 12713 16603 12771 16609
rect 13078 16600 13084 16652
rect 13136 16649 13142 16652
rect 13136 16643 13164 16649
rect 13152 16609 13164 16643
rect 13136 16603 13164 16609
rect 13136 16600 13142 16603
rect 13262 16600 13268 16652
rect 13320 16600 13326 16652
rect 5779 16535 5837 16541
rect 5902 16544 6224 16572
rect 750 16464 756 16516
rect 808 16504 814 16516
rect 1489 16507 1547 16513
rect 1489 16504 1501 16507
rect 808 16476 1501 16504
rect 808 16464 814 16476
rect 1489 16473 1501 16476
rect 1535 16473 1547 16507
rect 1489 16467 1547 16473
rect 5626 16464 5632 16516
rect 5684 16504 5690 16516
rect 5902 16504 5930 16544
rect 6546 16532 6552 16584
rect 6604 16572 6610 16584
rect 7343 16575 7401 16581
rect 7098 16572 7104 16574
rect 6604 16544 7104 16572
rect 6604 16532 6610 16544
rect 7098 16522 7104 16544
rect 7156 16572 7162 16574
rect 7343 16572 7355 16575
rect 7156 16544 7355 16572
rect 7156 16522 7162 16544
rect 7343 16541 7355 16544
rect 7389 16541 7401 16575
rect 7343 16535 7401 16541
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 9364 16544 9413 16572
rect 9364 16532 9370 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9674 16572 9680 16584
rect 9635 16544 9680 16572
rect 9401 16535 9459 16541
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 11238 16532 11244 16584
rect 11296 16572 11302 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11296 16544 11989 16572
rect 11296 16532 11302 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 11977 16535 12035 16541
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 5684 16476 5930 16504
rect 5684 16464 5690 16476
rect 7742 16464 7748 16516
rect 7800 16504 7806 16516
rect 10134 16504 10140 16516
rect 7800 16476 10140 16504
rect 7800 16464 7806 16476
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 9582 16436 9588 16448
rect 7156 16408 9588 16436
rect 7156 16396 7162 16408
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 12084 16436 12112 16535
rect 12986 16532 12992 16584
rect 13044 16532 13050 16584
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 12802 16436 12808 16448
rect 12084 16408 12808 16436
rect 12802 16396 12808 16408
rect 12860 16436 12866 16448
rect 13814 16436 13820 16448
rect 12860 16408 13820 16436
rect 12860 16396 12866 16408
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 1104 16346 14971 16368
rect 1104 16294 4376 16346
rect 4428 16294 4440 16346
rect 4492 16294 4504 16346
rect 4556 16294 4568 16346
rect 4620 16294 4632 16346
rect 4684 16294 7803 16346
rect 7855 16294 7867 16346
rect 7919 16294 7931 16346
rect 7983 16294 7995 16346
rect 8047 16294 8059 16346
rect 8111 16294 11230 16346
rect 11282 16294 11294 16346
rect 11346 16294 11358 16346
rect 11410 16294 11422 16346
rect 11474 16294 11486 16346
rect 11538 16294 14657 16346
rect 14709 16294 14721 16346
rect 14773 16294 14785 16346
rect 14837 16294 14849 16346
rect 14901 16294 14913 16346
rect 14965 16294 14971 16346
rect 1104 16272 14971 16294
rect 7834 16192 7840 16244
rect 7892 16232 7898 16244
rect 7892 16204 9996 16232
rect 7892 16192 7898 16204
rect 1673 16167 1731 16173
rect 1673 16133 1685 16167
rect 1719 16164 1731 16167
rect 7098 16164 7104 16176
rect 1719 16136 7104 16164
rect 1719 16133 1731 16136
rect 1673 16127 1731 16133
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 9309 16167 9367 16173
rect 9309 16133 9321 16167
rect 9355 16164 9367 16167
rect 9858 16164 9864 16176
rect 9355 16136 9864 16164
rect 9355 16133 9367 16136
rect 9309 16127 9367 16133
rect 9858 16124 9864 16136
rect 9916 16124 9922 16176
rect 9968 16164 9996 16204
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10413 16235 10471 16241
rect 10413 16232 10425 16235
rect 10100 16204 10425 16232
rect 10100 16192 10106 16204
rect 10413 16201 10425 16204
rect 10459 16201 10471 16235
rect 10413 16195 10471 16201
rect 12342 16192 12348 16244
rect 12400 16192 12406 16244
rect 14461 16235 14519 16241
rect 14461 16232 14473 16235
rect 12544 16204 14473 16232
rect 9968 16136 10088 16164
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1489 16099 1547 16105
rect 1489 16096 1501 16099
rect 900 16068 1501 16096
rect 900 16056 906 16068
rect 1489 16065 1501 16068
rect 1535 16065 1547 16099
rect 1489 16059 1547 16065
rect 7282 16056 7288 16108
rect 7340 16096 7346 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7340 16068 7481 16096
rect 7340 16056 7346 16068
rect 7469 16065 7481 16068
rect 7515 16096 7527 16099
rect 7515 16068 7880 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 15988 7564 16040
rect 7616 15988 7622 16040
rect 7653 16031 7711 16037
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 7742 16028 7748 16040
rect 7699 16000 7748 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 7852 16028 7880 16068
rect 8386 16056 8392 16108
rect 8444 16056 8450 16108
rect 8570 16105 8576 16108
rect 8527 16099 8576 16105
rect 8527 16065 8539 16099
rect 8573 16065 8576 16099
rect 8527 16059 8576 16065
rect 8570 16056 8576 16059
rect 8628 16056 8634 16108
rect 8662 16056 8668 16108
rect 8720 16056 8726 16108
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 9675 16099 9733 16105
rect 9675 16096 9687 16099
rect 9640 16068 9687 16096
rect 9640 16056 9646 16068
rect 9675 16065 9687 16068
rect 9721 16065 9733 16099
rect 9675 16059 9733 16065
rect 8202 16028 8208 16040
rect 7852 16000 8208 16028
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 9306 15988 9312 16040
rect 9364 16028 9370 16040
rect 9401 16031 9459 16037
rect 9401 16028 9413 16031
rect 9364 16000 9413 16028
rect 9364 15988 9370 16000
rect 9401 15997 9413 16000
rect 9447 15997 9459 16031
rect 10060 16028 10088 16136
rect 12544 16105 12572 16204
rect 14461 16201 14473 16204
rect 14507 16201 14519 16235
rect 14461 16195 14519 16201
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 12710 16096 12716 16108
rect 12667 16068 12716 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12710 16056 12716 16068
rect 12768 16056 12774 16108
rect 12802 16056 12808 16108
rect 12860 16056 12866 16108
rect 13814 16056 13820 16108
rect 13872 16056 13878 16108
rect 10060 16000 12848 16028
rect 9401 15991 9459 15997
rect 7576 15960 7604 15988
rect 12820 15972 12848 16000
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 13372 16000 13553 16028
rect 8113 15963 8171 15969
rect 8113 15960 8125 15963
rect 7576 15932 8125 15960
rect 8113 15929 8125 15932
rect 8159 15929 8171 15963
rect 8113 15923 8171 15929
rect 9048 15932 9444 15960
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 9048 15892 9076 15932
rect 2556 15864 9076 15892
rect 9416 15892 9444 15932
rect 12802 15920 12808 15972
rect 12860 15920 12866 15972
rect 13372 15960 13400 16000
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 13541 15991 13599 15997
rect 13630 15988 13636 16040
rect 13688 16037 13694 16040
rect 13688 16031 13716 16037
rect 13704 15997 13716 16031
rect 13688 15991 13716 15997
rect 13688 15988 13694 15991
rect 13188 15932 13400 15960
rect 9858 15892 9864 15904
rect 9416 15864 9864 15892
rect 2556 15852 2562 15864
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 13078 15892 13084 15904
rect 11664 15864 13084 15892
rect 11664 15852 11670 15864
rect 13078 15852 13084 15864
rect 13136 15892 13142 15904
rect 13188 15892 13216 15932
rect 13136 15864 13216 15892
rect 13136 15852 13142 15864
rect 1104 15802 14812 15824
rect 1104 15750 2663 15802
rect 2715 15750 2727 15802
rect 2779 15750 2791 15802
rect 2843 15750 2855 15802
rect 2907 15750 2919 15802
rect 2971 15750 6090 15802
rect 6142 15750 6154 15802
rect 6206 15750 6218 15802
rect 6270 15750 6282 15802
rect 6334 15750 6346 15802
rect 6398 15750 9517 15802
rect 9569 15750 9581 15802
rect 9633 15750 9645 15802
rect 9697 15750 9709 15802
rect 9761 15750 9773 15802
rect 9825 15750 12944 15802
rect 12996 15750 13008 15802
rect 13060 15750 13072 15802
rect 13124 15750 13136 15802
rect 13188 15750 13200 15802
rect 13252 15750 14812 15802
rect 1104 15728 14812 15750
rect 5626 15688 5632 15700
rect 5552 15660 5632 15688
rect 1302 15444 1308 15496
rect 1360 15484 1366 15496
rect 1397 15487 1455 15493
rect 1397 15484 1409 15487
rect 1360 15456 1409 15484
rect 1360 15444 1366 15456
rect 1397 15453 1409 15456
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 1671 15487 1729 15493
rect 1671 15453 1683 15487
rect 1717 15484 1729 15487
rect 2038 15484 2044 15496
rect 1717 15456 2044 15484
rect 1717 15453 1729 15456
rect 1671 15447 1729 15453
rect 2038 15444 2044 15456
rect 2096 15484 2102 15496
rect 2498 15484 2504 15496
rect 2096 15456 2504 15484
rect 2096 15444 2102 15456
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5552 15493 5580 15660
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 8386 15648 8392 15700
rect 8444 15688 8450 15700
rect 8444 15660 13216 15688
rect 8444 15648 8450 15660
rect 11606 15580 11612 15632
rect 11664 15620 11670 15632
rect 12161 15623 12219 15629
rect 12161 15620 12173 15623
rect 11664 15592 12173 15620
rect 11664 15580 11670 15592
rect 12161 15589 12173 15592
rect 12207 15589 12219 15623
rect 13188 15620 13216 15660
rect 13262 15648 13268 15700
rect 13320 15648 13326 15700
rect 14369 15691 14427 15697
rect 14369 15657 14381 15691
rect 14415 15657 14427 15691
rect 14369 15651 14427 15657
rect 14384 15620 14412 15651
rect 13188 15592 14412 15620
rect 12161 15583 12219 15589
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 11848 15524 11928 15552
rect 11848 15512 11854 15524
rect 5537 15487 5595 15493
rect 5537 15484 5549 15487
rect 5500 15456 5549 15484
rect 5500 15444 5506 15456
rect 5537 15453 5549 15456
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5811 15487 5869 15493
rect 5811 15453 5823 15487
rect 5857 15484 5869 15487
rect 6914 15484 6920 15496
rect 5857 15456 6920 15484
rect 5857 15453 5869 15456
rect 5811 15447 5869 15453
rect 6914 15444 6920 15456
rect 6972 15484 6978 15496
rect 7282 15484 7288 15496
rect 6972 15456 7288 15484
rect 6972 15444 6978 15456
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9306 15484 9312 15496
rect 8996 15456 9312 15484
rect 8996 15444 9002 15456
rect 9306 15444 9312 15456
rect 9364 15484 9370 15496
rect 9493 15487 9551 15493
rect 9493 15484 9505 15487
rect 9364 15456 9505 15484
rect 9364 15444 9370 15456
rect 9493 15453 9505 15456
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9735 15487 9793 15493
rect 9735 15453 9747 15487
rect 9781 15484 9793 15487
rect 9858 15484 9864 15496
rect 9781 15456 9864 15484
rect 9781 15453 9793 15456
rect 9735 15447 9793 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 11900 15484 11928 15524
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 12253 15555 12311 15561
rect 12253 15552 12265 15555
rect 12032 15524 12265 15552
rect 12032 15512 12038 15524
rect 12253 15521 12265 15524
rect 12299 15521 12311 15555
rect 12253 15515 12311 15521
rect 12495 15487 12553 15493
rect 12495 15484 12507 15487
rect 11900 15456 12507 15484
rect 5184 15416 5212 15444
rect 5184 15388 8524 15416
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15348 2467 15351
rect 2498 15348 2504 15360
rect 2455 15320 2504 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 2498 15308 2504 15320
rect 2556 15308 2562 15360
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 7190 15348 7196 15360
rect 6595 15320 7196 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 7190 15308 7196 15320
rect 7248 15308 7254 15360
rect 8496 15348 8524 15388
rect 8570 15376 8576 15428
rect 8628 15416 8634 15428
rect 11790 15416 11796 15428
rect 8628 15388 11796 15416
rect 8628 15376 8634 15388
rect 11790 15376 11796 15388
rect 11848 15376 11854 15428
rect 10410 15348 10416 15360
rect 8496 15320 10416 15348
rect 10410 15308 10416 15320
rect 10468 15308 10474 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 10686 15348 10692 15360
rect 10551 15320 10692 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 11900 15348 11928 15456
rect 12495 15453 12507 15456
rect 12541 15453 12553 15487
rect 12495 15447 12553 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14826 15484 14832 15496
rect 13771 15456 14832 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12342 15416 12348 15428
rect 12023 15388 12348 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12342 15376 12348 15388
rect 12400 15376 12406 15428
rect 14277 15419 14335 15425
rect 14277 15385 14289 15419
rect 14323 15416 14335 15419
rect 15102 15416 15108 15428
rect 14323 15388 15108 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 10928 15320 11928 15348
rect 10928 15308 10934 15320
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13817 15351 13875 15357
rect 13817 15348 13829 15351
rect 13228 15320 13829 15348
rect 13228 15308 13234 15320
rect 13817 15317 13829 15320
rect 13863 15317 13875 15351
rect 13817 15311 13875 15317
rect 1104 15258 14971 15280
rect 1104 15206 4376 15258
rect 4428 15206 4440 15258
rect 4492 15206 4504 15258
rect 4556 15206 4568 15258
rect 4620 15206 4632 15258
rect 4684 15206 7803 15258
rect 7855 15206 7867 15258
rect 7919 15206 7931 15258
rect 7983 15206 7995 15258
rect 8047 15206 8059 15258
rect 8111 15206 11230 15258
rect 11282 15206 11294 15258
rect 11346 15206 11358 15258
rect 11410 15206 11422 15258
rect 11474 15206 11486 15258
rect 11538 15206 14657 15258
rect 14709 15206 14721 15258
rect 14773 15206 14785 15258
rect 14837 15206 14849 15258
rect 14901 15206 14913 15258
rect 14965 15206 14971 15258
rect 1104 15184 14971 15206
rect 8570 15144 8576 15156
rect 7116 15116 8576 15144
rect 1671 15011 1729 15017
rect 1671 14977 1683 15011
rect 1717 15008 1729 15011
rect 2038 15008 2044 15020
rect 1717 14980 2044 15008
rect 1717 14977 1729 14980
rect 1671 14971 1729 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 1397 14943 1455 14949
rect 1397 14940 1409 14943
rect 1360 14912 1409 14940
rect 1360 14900 1366 14912
rect 1397 14909 1409 14912
rect 1443 14909 1455 14943
rect 1397 14903 1455 14909
rect 2056 14872 2084 14968
rect 7116 14949 7144 15116
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 13354 15144 13360 15156
rect 9416 15116 11284 15144
rect 7834 14968 7840 15020
rect 7892 14968 7898 15020
rect 7975 15011 8033 15017
rect 7975 14977 7987 15011
rect 8021 14977 8033 15011
rect 7975 14971 8033 14977
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 6932 14872 6960 14903
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7248 14912 7573 14940
rect 7248 14900 7254 14912
rect 7561 14909 7573 14912
rect 7607 14909 7619 14943
rect 7990 14940 8018 14971
rect 8110 14968 8116 15020
rect 8168 14968 8174 15020
rect 9416 14940 9444 15116
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 7990 14912 9444 14940
rect 9493 14943 9551 14949
rect 7561 14903 7619 14909
rect 9493 14909 9505 14943
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 7466 14872 7472 14884
rect 2056 14844 2774 14872
rect 6932 14844 7472 14872
rect 2406 14764 2412 14816
rect 2464 14764 2470 14816
rect 2746 14804 2774 14844
rect 7466 14832 7472 14844
rect 7524 14832 7530 14884
rect 8496 14844 9260 14872
rect 8496 14804 8524 14844
rect 9232 14816 9260 14844
rect 9306 14832 9312 14884
rect 9364 14872 9370 14884
rect 9508 14872 9536 14903
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 10428 14940 10456 14971
rect 10686 14968 10692 15020
rect 10744 14968 10750 15020
rect 11256 15008 11284 15116
rect 12452 15116 13360 15144
rect 11333 15079 11391 15085
rect 11333 15045 11345 15079
rect 11379 15076 11391 15079
rect 12452 15076 12480 15116
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 13814 15104 13820 15156
rect 13872 15104 13878 15156
rect 11379 15048 12480 15076
rect 12544 15048 13676 15076
rect 11379 15045 11391 15048
rect 11333 15039 11391 15045
rect 11698 15008 11704 15020
rect 11256 14980 11704 15008
rect 11698 14968 11704 14980
rect 11756 15008 11762 15020
rect 12342 15008 12348 15020
rect 11756 14980 12348 15008
rect 11756 14968 11762 14980
rect 12342 14968 12348 14980
rect 12400 14968 12406 15020
rect 12544 15017 12572 15048
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 13047 15011 13105 15017
rect 13047 15008 13059 15011
rect 12768 14980 13059 15008
rect 12768 14968 12774 14980
rect 13047 14977 13059 14980
rect 13093 14977 13105 15011
rect 13648 15008 13676 15048
rect 13722 15036 13728 15088
rect 13780 15076 13786 15088
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 13780 15048 14289 15076
rect 13780 15036 13786 15048
rect 14277 15045 14289 15048
rect 14323 15045 14335 15079
rect 14277 15039 14335 15045
rect 14182 15008 14188 15020
rect 13648 14980 14188 15008
rect 13047 14971 13105 14977
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 10284 14912 10456 14940
rect 10284 14900 10290 14912
rect 10502 14900 10508 14952
rect 10560 14949 10566 14952
rect 10560 14943 10588 14949
rect 10576 14909 10588 14943
rect 10560 14903 10588 14909
rect 10560 14900 10566 14903
rect 11974 14900 11980 14952
rect 12032 14940 12038 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12032 14912 12817 14940
rect 12032 14900 12038 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 9364 14844 9536 14872
rect 9364 14832 9370 14844
rect 10134 14832 10140 14884
rect 10192 14832 10198 14884
rect 2746 14776 8524 14804
rect 8754 14764 8760 14816
rect 8812 14764 8818 14816
rect 9214 14764 9220 14816
rect 9272 14764 9278 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12713 14807 12771 14813
rect 12713 14804 12725 14807
rect 12400 14776 12725 14804
rect 12400 14764 12406 14776
rect 12713 14773 12725 14776
rect 12759 14773 12771 14807
rect 12713 14767 12771 14773
rect 12894 14764 12900 14816
rect 12952 14804 12958 14816
rect 14369 14807 14427 14813
rect 14369 14804 14381 14807
rect 12952 14776 14381 14804
rect 12952 14764 12958 14776
rect 14369 14773 14381 14776
rect 14415 14773 14427 14807
rect 14369 14767 14427 14773
rect 1104 14714 14812 14736
rect 1104 14662 2663 14714
rect 2715 14662 2727 14714
rect 2779 14662 2791 14714
rect 2843 14662 2855 14714
rect 2907 14662 2919 14714
rect 2971 14662 6090 14714
rect 6142 14662 6154 14714
rect 6206 14662 6218 14714
rect 6270 14662 6282 14714
rect 6334 14662 6346 14714
rect 6398 14662 9517 14714
rect 9569 14662 9581 14714
rect 9633 14662 9645 14714
rect 9697 14662 9709 14714
rect 9761 14662 9773 14714
rect 9825 14662 12944 14714
rect 12996 14662 13008 14714
rect 13060 14662 13072 14714
rect 13124 14662 13136 14714
rect 13188 14662 13200 14714
rect 13252 14662 14812 14714
rect 1104 14640 14812 14662
rect 842 14560 848 14612
rect 900 14600 906 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 900 14572 1593 14600
rect 900 14560 906 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 2406 14560 2412 14612
rect 2464 14560 2470 14612
rect 3602 14560 3608 14612
rect 3660 14600 3666 14612
rect 7469 14603 7527 14609
rect 3660 14572 7144 14600
rect 3660 14560 3666 14572
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2424 14396 2452 14560
rect 7116 14532 7144 14572
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 8110 14600 8116 14612
rect 7515 14572 8116 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 8110 14560 8116 14572
rect 8168 14560 8174 14612
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8570 14600 8576 14612
rect 8352 14572 8576 14600
rect 8352 14560 8358 14572
rect 8570 14560 8576 14572
rect 8628 14600 8634 14612
rect 9953 14603 10011 14609
rect 8628 14572 9904 14600
rect 8628 14560 8634 14572
rect 8662 14532 8668 14544
rect 7116 14504 8668 14532
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 9876 14532 9904 14572
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10134 14600 10140 14612
rect 9999 14572 10140 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 12250 14600 12256 14612
rect 10520 14572 12256 14600
rect 10520 14532 10548 14572
rect 12250 14560 12256 14572
rect 12308 14560 12314 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13998 14600 14004 14612
rect 13219 14572 14004 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 9876 14504 10548 14532
rect 13538 14492 13544 14544
rect 13596 14532 13602 14544
rect 14461 14535 14519 14541
rect 14461 14532 14473 14535
rect 13596 14504 14473 14532
rect 13596 14492 13602 14504
rect 14461 14501 14473 14504
rect 14507 14501 14519 14535
rect 14461 14495 14519 14501
rect 7834 14424 7840 14476
rect 7892 14424 7898 14476
rect 13170 14424 13176 14476
rect 13228 14464 13234 14476
rect 13630 14464 13636 14476
rect 13228 14436 13636 14464
rect 13228 14424 13234 14436
rect 13630 14424 13636 14436
rect 13688 14464 13694 14476
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 13688 14436 13921 14464
rect 13688 14424 13694 14436
rect 13909 14433 13921 14436
rect 13955 14433 13967 14467
rect 13909 14427 13967 14433
rect 2271 14368 2452 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2498 14356 2504 14408
rect 2556 14356 2562 14408
rect 6362 14356 6368 14408
rect 6420 14396 6426 14408
rect 6457 14399 6515 14405
rect 6457 14396 6469 14399
rect 6420 14368 6469 14396
rect 6420 14356 6426 14368
rect 6457 14365 6469 14368
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6715 14369 6773 14375
rect 1489 14331 1547 14337
rect 1489 14297 1501 14331
rect 1535 14328 1547 14331
rect 6715 14335 6727 14369
rect 6761 14366 6773 14369
rect 6761 14335 6776 14366
rect 6715 14329 6776 14335
rect 6748 14328 6776 14329
rect 7190 14328 7196 14340
rect 1535 14300 2360 14328
rect 6748 14300 7196 14328
rect 1535 14297 1547 14300
rect 1489 14291 1547 14297
rect 2038 14220 2044 14272
rect 2096 14220 2102 14272
rect 2332 14269 2360 14300
rect 7190 14288 7196 14300
rect 7248 14328 7254 14340
rect 7650 14328 7656 14340
rect 7248 14300 7656 14328
rect 7248 14288 7254 14300
rect 7650 14288 7656 14300
rect 7708 14288 7714 14340
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14229 2375 14263
rect 7852 14260 7880 14424
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8938 14396 8944 14408
rect 8444 14368 8944 14396
rect 8444 14356 8450 14368
rect 8938 14356 8944 14368
rect 8996 14396 9002 14408
rect 9214 14405 9220 14408
rect 9183 14399 9220 14405
rect 8996 14368 9150 14396
rect 8996 14356 9002 14368
rect 8570 14288 8576 14340
rect 8628 14328 8634 14340
rect 9030 14328 9036 14340
rect 8628 14300 9036 14328
rect 8628 14288 8634 14300
rect 9030 14288 9036 14300
rect 9088 14288 9094 14340
rect 9122 14328 9150 14368
rect 9183 14365 9195 14399
rect 9183 14359 9220 14365
rect 9214 14356 9220 14359
rect 9272 14356 9278 14408
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 12066 14405 12072 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10284 14368 10425 14396
rect 10284 14356 10290 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10687 14399 10745 14405
rect 10687 14365 10699 14399
rect 10733 14392 10745 14399
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 10796 14392 11008 14396
rect 10733 14368 11008 14392
rect 10733 14365 10824 14368
rect 10687 14364 10824 14365
rect 10687 14359 10745 14364
rect 10042 14328 10048 14340
rect 9122 14300 10048 14328
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10428 14328 10456 14359
rect 10980 14340 11008 14368
rect 11070 14368 11805 14396
rect 10428 14300 10916 14328
rect 10778 14260 10784 14272
rect 7852 14232 10784 14260
rect 2317 14223 2375 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10888 14260 10916 14300
rect 10962 14288 10968 14340
rect 11020 14288 11026 14340
rect 11070 14260 11098 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 12035 14399 12072 14405
rect 12035 14365 12047 14399
rect 12035 14359 12072 14365
rect 12066 14356 12072 14359
rect 12124 14356 12130 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 12406 14368 13369 14396
rect 11146 14288 11152 14340
rect 11204 14328 11210 14340
rect 12406 14328 12434 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 14826 14396 14832 14408
rect 13771 14368 14832 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 11204 14300 12434 14328
rect 11204 14288 11210 14300
rect 14274 14288 14280 14340
rect 14332 14288 14338 14340
rect 10888 14232 11098 14260
rect 11425 14263 11483 14269
rect 11425 14229 11437 14263
rect 11471 14260 11483 14263
rect 11698 14260 11704 14272
rect 11471 14232 11704 14260
rect 11471 14229 11483 14232
rect 11425 14223 11483 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 12805 14263 12863 14269
rect 12805 14260 12817 14263
rect 12768 14232 12817 14260
rect 12768 14220 12774 14232
rect 12805 14229 12817 14232
rect 12851 14229 12863 14263
rect 12805 14223 12863 14229
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13630 14260 13636 14272
rect 13504 14232 13636 14260
rect 13504 14220 13510 14232
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 1104 14170 14971 14192
rect 1104 14118 4376 14170
rect 4428 14118 4440 14170
rect 4492 14118 4504 14170
rect 4556 14118 4568 14170
rect 4620 14118 4632 14170
rect 4684 14118 7803 14170
rect 7855 14118 7867 14170
rect 7919 14118 7931 14170
rect 7983 14118 7995 14170
rect 8047 14118 8059 14170
rect 8111 14118 11230 14170
rect 11282 14118 11294 14170
rect 11346 14118 11358 14170
rect 11410 14118 11422 14170
rect 11474 14118 11486 14170
rect 11538 14118 14657 14170
rect 14709 14118 14721 14170
rect 14773 14118 14785 14170
rect 14837 14118 14849 14170
rect 14901 14118 14913 14170
rect 14965 14118 14971 14170
rect 1104 14096 14971 14118
rect 2038 14016 2044 14068
rect 2096 14016 2102 14068
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14025 7435 14059
rect 7377 14019 7435 14025
rect 2056 13988 2084 14016
rect 2409 13991 2467 13997
rect 2409 13988 2421 13991
rect 2056 13960 2421 13988
rect 2409 13957 2421 13960
rect 2455 13957 2467 13991
rect 2409 13951 2467 13957
rect 6454 13948 6460 14000
rect 6512 13948 6518 14000
rect 1854 13880 1860 13932
rect 1912 13880 1918 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6362 13920 6368 13932
rect 5500 13892 6368 13920
rect 5500 13880 5506 13892
rect 6362 13880 6368 13892
rect 6420 13880 6426 13932
rect 6472 13920 6500 13948
rect 6638 13920 6644 13932
rect 6472 13892 6644 13920
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 7392 13920 7420 14019
rect 7466 14016 7472 14068
rect 7524 14056 7530 14068
rect 9214 14056 9220 14068
rect 7524 14028 9220 14056
rect 7524 14016 7530 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9861 14059 9919 14065
rect 9861 14025 9873 14059
rect 9907 14056 9919 14059
rect 11146 14056 11152 14068
rect 9907 14028 11152 14056
rect 9907 14025 9919 14028
rect 9861 14019 9919 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11698 14016 11704 14068
rect 11756 14016 11762 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12216 14028 13768 14056
rect 12216 14016 12222 14028
rect 9950 13948 9956 14000
rect 10008 13988 10014 14000
rect 10008 13960 11652 13988
rect 10008 13948 10014 13960
rect 7392 13892 8432 13920
rect 7116 13852 7144 13880
rect 7650 13852 7656 13864
rect 7116 13824 7656 13852
rect 7650 13812 7656 13824
rect 7708 13852 7714 13864
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7708 13824 8033 13852
rect 7708 13812 7714 13824
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8294 13852 8300 13864
rect 8260 13812 8300 13852
rect 8352 13812 8358 13864
rect 8404 13852 8432 13892
rect 9030 13880 9036 13932
rect 9088 13929 9094 13932
rect 9088 13923 9116 13929
rect 9104 13889 9116 13923
rect 9088 13883 9116 13889
rect 9088 13880 9094 13883
rect 9214 13880 9220 13932
rect 9272 13880 9278 13932
rect 10319 13923 10377 13929
rect 10319 13889 10331 13923
rect 10365 13920 10377 13923
rect 10410 13920 10416 13932
rect 10365 13892 10416 13920
rect 10365 13889 10377 13892
rect 10319 13883 10377 13889
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 8404 13824 8677 13852
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 8938 13812 8944 13864
rect 8996 13812 9002 13864
rect 10042 13812 10048 13864
rect 10100 13812 10106 13864
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 11624 13852 11652 13960
rect 11716 13920 11744 14016
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 13630 13988 13636 14000
rect 13403 13960 13636 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 11716 13892 11836 13920
rect 11698 13852 11704 13864
rect 11624 13824 11704 13852
rect 11698 13812 11704 13824
rect 11756 13812 11762 13864
rect 11808 13852 11836 13892
rect 12710 13880 12716 13932
rect 12768 13880 12774 13932
rect 13740 13864 13768 14028
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11808 13824 12173 13852
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 12437 13855 12495 13861
rect 12437 13852 12449 13855
rect 12308 13824 12449 13852
rect 12308 13812 12314 13824
rect 12437 13821 12449 13824
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 12526 13812 12532 13864
rect 12584 13861 12590 13864
rect 12584 13855 12612 13861
rect 12600 13821 12612 13855
rect 12584 13815 12612 13821
rect 12584 13812 12590 13815
rect 13630 13812 13636 13864
rect 13688 13812 13694 13864
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13780 13824 13921 13852
rect 13780 13812 13786 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 13909 13815 13967 13821
rect 1946 13676 1952 13728
rect 2004 13676 2010 13728
rect 2498 13676 2504 13728
rect 2556 13676 2562 13728
rect 8266 13716 8294 13812
rect 9030 13716 9036 13728
rect 8266 13688 9036 13716
rect 9030 13676 9036 13688
rect 9088 13676 9094 13728
rect 10060 13716 10088 13812
rect 11974 13784 11980 13796
rect 10702 13756 11980 13784
rect 10702 13716 10730 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 10060 13688 10730 13716
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13716 11115 13719
rect 11422 13716 11428 13728
rect 11103 13688 11428 13716
rect 11103 13685 11115 13688
rect 11057 13679 11115 13685
rect 11422 13676 11428 13688
rect 11480 13676 11486 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 13354 13716 13360 13728
rect 13228 13688 13360 13716
rect 13228 13676 13234 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 1104 13626 14812 13648
rect 1104 13574 2663 13626
rect 2715 13574 2727 13626
rect 2779 13574 2791 13626
rect 2843 13574 2855 13626
rect 2907 13574 2919 13626
rect 2971 13574 6090 13626
rect 6142 13574 6154 13626
rect 6206 13574 6218 13626
rect 6270 13574 6282 13626
rect 6334 13574 6346 13626
rect 6398 13574 9517 13626
rect 9569 13574 9581 13626
rect 9633 13574 9645 13626
rect 9697 13574 9709 13626
rect 9761 13574 9773 13626
rect 9825 13574 12944 13626
rect 12996 13574 13008 13626
rect 13060 13574 13072 13626
rect 13124 13574 13136 13626
rect 13188 13574 13200 13626
rect 13252 13574 14812 13626
rect 1104 13552 14812 13574
rect 5442 13512 5448 13524
rect 1412 13484 5448 13512
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 1412 13317 1440 13484
rect 4724 13385 4752 13484
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 7466 13512 7472 13524
rect 5767 13484 7472 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 8386 13512 8392 13524
rect 7576 13484 8392 13512
rect 7576 13444 7604 13484
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8754 13472 8760 13524
rect 8812 13512 8818 13524
rect 8812 13484 13860 13512
rect 8812 13472 8818 13484
rect 13832 13444 13860 13484
rect 13906 13472 13912 13524
rect 13964 13472 13970 13524
rect 14093 13515 14151 13521
rect 14093 13481 14105 13515
rect 14139 13512 14151 13515
rect 14366 13512 14372 13524
rect 14139 13484 14372 13512
rect 14139 13481 14151 13484
rect 14093 13475 14151 13481
rect 14366 13472 14372 13484
rect 14424 13472 14430 13524
rect 7484 13416 7604 13444
rect 10612 13416 12848 13444
rect 13832 13416 14320 13444
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13345 4767 13379
rect 4709 13339 4767 13345
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 1360 13280 1409 13308
rect 1360 13268 1366 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1397 13271 1455 13277
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 4246 13308 4252 13320
rect 2188 13280 4252 13308
rect 2188 13268 2194 13280
rect 4246 13268 4252 13280
rect 4304 13308 4310 13320
rect 4951 13311 5009 13317
rect 4951 13308 4963 13311
rect 4304 13280 4963 13308
rect 4304 13268 4310 13280
rect 4951 13277 4963 13280
rect 4997 13277 5009 13311
rect 4951 13271 5009 13277
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 6086 13308 6092 13320
rect 5684 13280 6092 13308
rect 5684 13268 5690 13280
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 6347 13281 6405 13287
rect 1688 13240 1716 13268
rect 6347 13247 6359 13281
rect 6393 13278 6405 13281
rect 6393 13247 6408 13278
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 7484 13317 7512 13416
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 6512 13280 7481 13308
rect 6512 13268 6518 13280
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7711 13311 7769 13317
rect 7711 13308 7723 13311
rect 7469 13271 7527 13277
rect 7576 13280 7723 13308
rect 6347 13241 6408 13247
rect 6380 13240 6408 13241
rect 6730 13240 6736 13252
rect 1688 13212 6316 13240
rect 6380 13212 6736 13240
rect 2409 13175 2467 13181
rect 2409 13141 2421 13175
rect 2455 13172 2467 13175
rect 2498 13172 2504 13184
rect 2455 13144 2504 13172
rect 2455 13141 2467 13144
rect 2409 13135 2467 13141
rect 2498 13132 2504 13144
rect 2556 13132 2562 13184
rect 6288 13172 6316 13212
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 7576 13240 7604 13280
rect 7711 13277 7723 13280
rect 7757 13277 7769 13311
rect 7711 13271 7769 13277
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 9548 13280 9689 13308
rect 9548 13268 9554 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 9951 13311 10009 13317
rect 9951 13277 9963 13311
rect 9997 13308 10009 13311
rect 10410 13308 10416 13320
rect 9997 13280 10416 13308
rect 9997 13277 10009 13280
rect 9951 13271 10009 13277
rect 7024 13212 7604 13240
rect 9692 13240 9720 13271
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10226 13240 10232 13252
rect 9692 13212 10232 13240
rect 7024 13172 7052 13212
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 6288 13144 7052 13172
rect 7098 13132 7104 13184
rect 7156 13132 7162 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8754 13172 8760 13184
rect 8527 13144 8760 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8754 13132 8760 13144
rect 8812 13132 8818 13184
rect 10134 13132 10140 13184
rect 10192 13172 10198 13184
rect 10612 13172 10640 13416
rect 11514 13336 11520 13388
rect 11572 13376 11578 13388
rect 11572 13348 12204 13376
rect 11572 13336 11578 13348
rect 12176 13320 12204 13348
rect 12710 13336 12716 13388
rect 12768 13336 12774 13388
rect 12820 13376 12848 13416
rect 12986 13376 12992 13388
rect 12820 13348 12992 13376
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 13078 13336 13084 13388
rect 13136 13385 13142 13388
rect 13136 13379 13164 13385
rect 13152 13345 13164 13379
rect 13136 13339 13164 13345
rect 13136 13336 13142 13339
rect 11790 13268 11796 13320
rect 11848 13268 11854 13320
rect 12066 13268 12072 13320
rect 12124 13268 12130 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 12216 13280 12265 13308
rect 12216 13268 12222 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 13262 13268 13268 13320
rect 13320 13268 13326 13320
rect 14292 13317 14320 13416
rect 15286 13336 15292 13388
rect 15344 13376 15350 13388
rect 15838 13376 15844 13388
rect 15344 13348 15844 13376
rect 15344 13336 15350 13348
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 10192 13144 10640 13172
rect 10192 13132 10198 13144
rect 10686 13132 10692 13184
rect 10744 13132 10750 13184
rect 11808 13172 11836 13268
rect 14458 13240 14464 13252
rect 14016 13212 14464 13240
rect 14016 13172 14044 13212
rect 14458 13200 14464 13212
rect 14516 13200 14522 13252
rect 11808 13144 14044 13172
rect 1104 13082 14971 13104
rect 1104 13030 4376 13082
rect 4428 13030 4440 13082
rect 4492 13030 4504 13082
rect 4556 13030 4568 13082
rect 4620 13030 4632 13082
rect 4684 13030 7803 13082
rect 7855 13030 7867 13082
rect 7919 13030 7931 13082
rect 7983 13030 7995 13082
rect 8047 13030 8059 13082
rect 8111 13030 11230 13082
rect 11282 13030 11294 13082
rect 11346 13030 11358 13082
rect 11410 13030 11422 13082
rect 11474 13030 11486 13082
rect 11538 13030 14657 13082
rect 14709 13030 14721 13082
rect 14773 13030 14785 13082
rect 14837 13030 14849 13082
rect 14901 13030 14913 13082
rect 14965 13030 14971 13082
rect 1104 13008 14971 13030
rect 1762 12928 1768 12980
rect 1820 12968 1826 12980
rect 6730 12968 6736 12980
rect 1820 12940 6736 12968
rect 1820 12928 1826 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7098 12928 7104 12980
rect 7156 12928 7162 12980
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 7616 12940 9260 12968
rect 7616 12928 7622 12940
rect 1780 12900 1808 12928
rect 1686 12872 1808 12900
rect 1686 12871 1714 12872
rect 1655 12865 1714 12871
rect 1655 12831 1667 12865
rect 1701 12834 1714 12865
rect 1701 12831 1713 12834
rect 1655 12825 1713 12831
rect 7116 12832 7144 12928
rect 9232 12900 9260 12940
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 9508 12940 11989 12968
rect 9508 12900 9536 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 12253 12971 12311 12977
rect 11977 12931 12035 12937
rect 12082 12940 12204 12968
rect 9232 12872 9536 12900
rect 7116 12804 7880 12832
rect 1302 12724 1308 12776
rect 1360 12764 1366 12776
rect 1397 12767 1455 12773
rect 1397 12764 1409 12767
rect 1360 12736 1409 12764
rect 1360 12724 1366 12736
rect 1397 12733 1409 12736
rect 1443 12733 1455 12767
rect 1397 12727 1455 12733
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 7650 12764 7656 12776
rect 7607 12736 7656 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 7650 12724 7656 12736
rect 7708 12724 7714 12776
rect 7745 12767 7803 12773
rect 7745 12733 7757 12767
rect 7791 12733 7803 12767
rect 7852 12764 7880 12804
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 8570 12792 8576 12844
rect 8628 12841 8634 12844
rect 8628 12835 8656 12841
rect 8644 12801 8656 12835
rect 8628 12795 8656 12801
rect 8628 12792 8634 12795
rect 8754 12792 8760 12844
rect 8812 12792 8818 12844
rect 9766 12832 9772 12844
rect 9727 12804 9772 12832
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 11790 12792 11796 12844
rect 11848 12792 11854 12844
rect 12082 12842 12110 12940
rect 12176 12900 12204 12940
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12434 12968 12440 12980
rect 12299 12940 12440 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13357 12971 13415 12977
rect 13357 12968 13369 12971
rect 12768 12940 13369 12968
rect 12768 12928 12774 12940
rect 13357 12937 13369 12940
rect 13403 12937 13415 12971
rect 13357 12931 13415 12937
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 12342 12900 12348 12912
rect 12176 12872 12348 12900
rect 12342 12860 12348 12872
rect 12400 12860 12406 12912
rect 12634 12872 13032 12900
rect 12634 12871 12662 12872
rect 12603 12865 12662 12871
rect 12082 12841 12112 12842
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12603 12831 12615 12865
rect 12649 12834 12662 12865
rect 12649 12831 12661 12834
rect 12603 12825 12661 12831
rect 13004 12832 13032 12872
rect 13170 12860 13176 12912
rect 13228 12900 13234 12912
rect 13924 12900 13952 12931
rect 14458 12928 14464 12980
rect 14516 12928 14522 12980
rect 13228 12872 13952 12900
rect 13228 12860 13234 12872
rect 13725 12835 13783 12841
rect 13004 12804 13584 12832
rect 12069 12795 12127 12801
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 7852 12736 8217 12764
rect 7745 12727 7803 12733
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 7466 12656 7472 12708
rect 7524 12696 7530 12708
rect 7760 12696 7788 12727
rect 9398 12724 9404 12776
rect 9456 12764 9462 12776
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9456 12736 9505 12764
rect 9456 12724 9462 12736
rect 9493 12733 9505 12736
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12345 12767 12403 12773
rect 12345 12764 12357 12767
rect 12032 12736 12357 12764
rect 12032 12724 12038 12736
rect 12345 12733 12357 12736
rect 12391 12733 12403 12767
rect 13556 12764 13584 12804
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 13906 12832 13912 12844
rect 13771 12804 13912 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 13998 12792 14004 12844
rect 14056 12792 14062 12844
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 15102 12832 15108 12844
rect 14323 12804 15108 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 14182 12764 14188 12776
rect 13556 12736 14188 12764
rect 12345 12727 12403 12733
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 7524 12668 7788 12696
rect 7524 12656 7530 12668
rect 13538 12656 13544 12708
rect 13596 12696 13602 12708
rect 13814 12696 13820 12708
rect 13596 12668 13820 12696
rect 13596 12656 13602 12668
rect 13814 12656 13820 12668
rect 13872 12656 13878 12708
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 7006 12588 7012 12640
rect 7064 12628 7070 12640
rect 7650 12628 7656 12640
rect 7064 12600 7656 12628
rect 7064 12588 7070 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 9950 12628 9956 12640
rect 7984 12600 9956 12628
rect 7984 12588 7990 12600
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 10502 12588 10508 12640
rect 10560 12588 10566 12640
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 10652 12600 14197 12628
rect 10652 12588 10658 12600
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14185 12591 14243 12597
rect 1104 12538 14812 12560
rect 1104 12486 2663 12538
rect 2715 12486 2727 12538
rect 2779 12486 2791 12538
rect 2843 12486 2855 12538
rect 2907 12486 2919 12538
rect 2971 12486 6090 12538
rect 6142 12486 6154 12538
rect 6206 12486 6218 12538
rect 6270 12486 6282 12538
rect 6334 12486 6346 12538
rect 6398 12486 9517 12538
rect 9569 12486 9581 12538
rect 9633 12486 9645 12538
rect 9697 12486 9709 12538
rect 9761 12486 9773 12538
rect 9825 12486 12944 12538
rect 12996 12486 13008 12538
rect 13060 12486 13072 12538
rect 13124 12486 13136 12538
rect 13188 12486 13200 12538
rect 13252 12486 14812 12538
rect 1104 12464 14812 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2317 12427 2375 12433
rect 2317 12424 2329 12427
rect 1912 12396 2329 12424
rect 1912 12384 1918 12396
rect 2317 12393 2329 12396
rect 2363 12393 2375 12427
rect 2317 12387 2375 12393
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 9674 12424 9680 12436
rect 5040 12396 9680 12424
rect 5040 12384 5046 12396
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 13449 12427 13507 12433
rect 11664 12396 13216 12424
rect 11664 12384 11670 12396
rect 7374 12316 7380 12368
rect 7432 12356 7438 12368
rect 13188 12356 13216 12396
rect 13449 12393 13461 12427
rect 13495 12424 13507 12427
rect 14090 12424 14096 12436
rect 13495 12396 14096 12424
rect 13495 12393 13507 12396
rect 13449 12387 13507 12393
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 15930 12384 15936 12436
rect 15988 12384 15994 12436
rect 13909 12359 13967 12365
rect 7432 12328 7696 12356
rect 13188 12328 13492 12356
rect 7432 12316 7438 12328
rect 7558 12248 7564 12300
rect 7616 12248 7622 12300
rect 7668 12288 7696 12328
rect 13464 12300 13492 12328
rect 13909 12325 13921 12359
rect 13955 12356 13967 12359
rect 15948 12356 15976 12384
rect 13955 12328 15976 12356
rect 13955 12325 13967 12328
rect 13909 12319 13967 12325
rect 7926 12288 7932 12300
rect 7984 12297 7990 12300
rect 7984 12291 8012 12297
rect 7668 12260 7932 12288
rect 7926 12248 7932 12260
rect 8000 12257 8012 12291
rect 7984 12251 8012 12257
rect 7984 12248 7990 12251
rect 10318 12248 10324 12300
rect 10376 12248 10382 12300
rect 10870 12248 10876 12300
rect 10928 12288 10934 12300
rect 10928 12260 11282 12288
rect 10928 12248 10934 12260
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2406 12220 2412 12232
rect 2271 12192 2412 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2498 12180 2504 12232
rect 2556 12180 2562 12232
rect 6730 12180 6736 12232
rect 6788 12220 6794 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6788 12192 6929 12220
rect 6788 12180 6794 12192
rect 6917 12189 6929 12192
rect 6963 12189 6975 12223
rect 6917 12183 6975 12189
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 7101 12223 7159 12229
rect 7101 12220 7113 12223
rect 7064 12192 7113 12220
rect 7064 12180 7070 12192
rect 7101 12189 7113 12192
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7834 12180 7840 12232
rect 7892 12180 7898 12232
rect 8110 12180 8116 12232
rect 8168 12180 8174 12232
rect 11254 12220 11282 12260
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 13354 12288 13360 12300
rect 12544 12260 13360 12288
rect 12544 12229 12572 12260
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 13446 12248 13452 12300
rect 13504 12248 13510 12300
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 9968 12192 11192 12220
rect 11254 12192 11805 12220
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12152 1547 12155
rect 9968 12152 9996 12192
rect 1535 12124 2084 12152
rect 1535 12121 1547 12124
rect 1489 12115 1547 12121
rect 842 12044 848 12096
rect 900 12084 906 12096
rect 2056 12093 2084 12124
rect 8772 12124 9996 12152
rect 10045 12155 10103 12161
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 900 12056 1593 12084
rect 900 12044 906 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12053 2099 12087
rect 2041 12047 2099 12053
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 8386 12084 8392 12096
rect 7892 12056 8392 12084
rect 7892 12044 7898 12056
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 8772 12093 8800 12124
rect 10045 12121 10057 12155
rect 10091 12121 10103 12155
rect 10045 12115 10103 12121
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10410 12152 10416 12164
rect 10183 12124 10416 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 8757 12087 8815 12093
rect 8757 12053 8769 12087
rect 8803 12053 8815 12087
rect 8757 12047 8815 12053
rect 9766 12044 9772 12096
rect 9824 12044 9830 12096
rect 9950 12044 9956 12096
rect 10008 12084 10014 12096
rect 10060 12084 10088 12115
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 10505 12155 10563 12161
rect 10505 12121 10517 12155
rect 10551 12121 10563 12155
rect 10505 12115 10563 12121
rect 10008 12056 10088 12084
rect 10520 12084 10548 12115
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 10836 12124 11100 12152
rect 10836 12112 10842 12124
rect 10686 12084 10692 12096
rect 10520 12056 10692 12084
rect 10008 12044 10014 12056
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 10870 12044 10876 12096
rect 10928 12044 10934 12096
rect 11072 12093 11100 12124
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12053 11115 12087
rect 11164 12084 11192 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12616 12180 12622 12232
rect 12674 12229 12680 12232
rect 12674 12223 12704 12229
rect 12692 12189 12704 12223
rect 12674 12183 12704 12189
rect 12674 12180 12680 12183
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 13740 12152 13768 12183
rect 14274 12180 14280 12232
rect 14332 12180 14338 12232
rect 13280 12124 13768 12152
rect 13280 12084 13308 12124
rect 11164 12056 13308 12084
rect 11057 12047 11115 12053
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 13872 12056 14473 12084
rect 13872 12044 13878 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 1104 11994 14971 12016
rect 1104 11942 4376 11994
rect 4428 11942 4440 11994
rect 4492 11942 4504 11994
rect 4556 11942 4568 11994
rect 4620 11942 4632 11994
rect 4684 11942 7803 11994
rect 7855 11942 7867 11994
rect 7919 11942 7931 11994
rect 7983 11942 7995 11994
rect 8047 11942 8059 11994
rect 8111 11942 11230 11994
rect 11282 11942 11294 11994
rect 11346 11942 11358 11994
rect 11410 11942 11422 11994
rect 11474 11942 11486 11994
rect 11538 11942 14657 11994
rect 14709 11942 14721 11994
rect 14773 11942 14785 11994
rect 14837 11942 14849 11994
rect 14901 11942 14913 11994
rect 14965 11942 14971 11994
rect 1104 11920 14971 11942
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 7745 11883 7803 11889
rect 5592 11852 7144 11880
rect 5592 11840 5598 11852
rect 3786 11772 3792 11824
rect 3844 11812 3850 11824
rect 3844 11784 6960 11812
rect 3844 11772 3850 11784
rect 6932 11756 6960 11784
rect 1486 11704 1492 11756
rect 1544 11704 1550 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 5644 11716 6745 11744
rect 5644 11688 5672 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7007 11747 7065 11753
rect 7007 11744 7019 11747
rect 6972 11716 7019 11744
rect 6972 11704 6978 11716
rect 7007 11713 7019 11716
rect 7053 11713 7065 11747
rect 7116 11744 7144 11852
rect 7745 11849 7757 11883
rect 7791 11880 7803 11883
rect 8202 11880 8208 11892
rect 7791 11852 8208 11880
rect 7791 11849 7803 11852
rect 7745 11843 7803 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 10134 11880 10140 11892
rect 8444 11852 10140 11880
rect 8444 11840 8450 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 10778 11840 10784 11892
rect 10836 11880 10842 11892
rect 11146 11880 11152 11892
rect 10836 11852 11152 11880
rect 10836 11840 10842 11852
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11606 11840 11612 11892
rect 11664 11880 11670 11892
rect 13354 11880 13360 11892
rect 11664 11852 13360 11880
rect 11664 11840 11670 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 15562 11880 15568 11892
rect 14415 11852 15568 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 7282 11772 7288 11824
rect 7340 11812 7346 11824
rect 10870 11812 10876 11824
rect 7340 11784 8984 11812
rect 7340 11772 7346 11784
rect 8846 11744 8852 11756
rect 7116 11716 8852 11744
rect 7007 11707 7065 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 8956 11744 8984 11784
rect 9876 11784 10876 11812
rect 9876 11756 9904 11784
rect 10870 11772 10876 11784
rect 10928 11772 10934 11824
rect 9091 11747 9149 11753
rect 9091 11744 9103 11747
rect 8956 11716 9103 11744
rect 9091 11713 9103 11716
rect 9137 11713 9149 11747
rect 9091 11707 9149 11713
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 10686 11704 10692 11756
rect 10744 11744 10750 11756
rect 12253 11747 12311 11753
rect 10744 11716 11192 11744
rect 10744 11704 10750 11716
rect 11164 11688 11192 11716
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12342 11744 12348 11756
rect 12299 11716 12348 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 12713 11747 12771 11753
rect 12713 11744 12725 11747
rect 12452 11716 12725 11744
rect 5626 11636 5632 11688
rect 5684 11636 5690 11688
rect 9766 11636 9772 11688
rect 9824 11676 9830 11688
rect 10870 11676 10876 11688
rect 9824 11648 10876 11676
rect 9824 11636 9830 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 12452 11676 12480 11716
rect 12713 11713 12725 11716
rect 12759 11713 12771 11747
rect 12713 11707 12771 11713
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 11204 11648 12480 11676
rect 12529 11679 12587 11685
rect 11204 11636 11210 11648
rect 12529 11645 12541 11679
rect 12575 11645 12587 11679
rect 12529 11639 12587 11645
rect 6730 11568 6736 11620
rect 6788 11568 6794 11620
rect 12544 11608 12572 11639
rect 13538 11636 13544 11688
rect 13596 11685 13602 11688
rect 13596 11679 13624 11685
rect 13612 11645 13624 11679
rect 13596 11639 13624 11645
rect 13596 11636 13602 11639
rect 13722 11636 13728 11688
rect 13780 11636 13786 11688
rect 12710 11608 12716 11620
rect 9508 11580 12112 11608
rect 12544 11580 12716 11608
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 900 11512 1593 11540
rect 900 11500 906 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 6748 11540 6776 11568
rect 9508 11540 9536 11580
rect 12084 11552 12112 11580
rect 12710 11568 12716 11580
rect 12768 11568 12774 11620
rect 13173 11611 13231 11617
rect 13173 11577 13185 11611
rect 13219 11608 13231 11611
rect 13262 11608 13268 11620
rect 13219 11580 13268 11608
rect 13219 11577 13231 11580
rect 13173 11571 13231 11577
rect 13262 11568 13268 11580
rect 13320 11568 13326 11620
rect 6748 11512 9536 11540
rect 9861 11543 9919 11549
rect 1581 11503 1639 11509
rect 9861 11509 9873 11543
rect 9907 11540 9919 11543
rect 10594 11540 10600 11552
rect 9907 11512 10600 11540
rect 9907 11509 9919 11512
rect 9861 11503 9919 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12437 11543 12495 11549
rect 12437 11540 12449 11543
rect 12124 11512 12449 11540
rect 12124 11500 12130 11512
rect 12437 11509 12449 11512
rect 12483 11509 12495 11543
rect 12437 11503 12495 11509
rect 12894 11500 12900 11552
rect 12952 11540 12958 11552
rect 13446 11540 13452 11552
rect 12952 11512 13452 11540
rect 12952 11500 12958 11512
rect 13446 11500 13452 11512
rect 13504 11500 13510 11552
rect 1104 11450 14812 11472
rect 1104 11398 2663 11450
rect 2715 11398 2727 11450
rect 2779 11398 2791 11450
rect 2843 11398 2855 11450
rect 2907 11398 2919 11450
rect 2971 11398 6090 11450
rect 6142 11398 6154 11450
rect 6206 11398 6218 11450
rect 6270 11398 6282 11450
rect 6334 11398 6346 11450
rect 6398 11398 9517 11450
rect 9569 11398 9581 11450
rect 9633 11398 9645 11450
rect 9697 11398 9709 11450
rect 9761 11398 9773 11450
rect 9825 11398 12944 11450
rect 12996 11398 13008 11450
rect 13060 11398 13072 11450
rect 13124 11398 13136 11450
rect 13188 11398 13200 11450
rect 13252 11398 14812 11450
rect 1104 11376 14812 11398
rect 5718 11296 5724 11348
rect 5776 11336 5782 11348
rect 6641 11339 6699 11345
rect 5776 11308 6500 11336
rect 5776 11296 5782 11308
rect 6472 11212 6500 11308
rect 6641 11305 6653 11339
rect 6687 11336 6699 11339
rect 7558 11336 7564 11348
rect 6687 11308 7564 11336
rect 6687 11305 6699 11308
rect 6641 11299 6699 11305
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 9674 11336 9680 11348
rect 8904 11308 9680 11336
rect 8904 11296 8910 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10686 11336 10692 11348
rect 9784 11308 10692 11336
rect 5626 11160 5632 11212
rect 5684 11160 5690 11212
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 9784 11200 9812 11308
rect 10686 11296 10692 11308
rect 10744 11336 10750 11348
rect 11238 11336 11244 11348
rect 10744 11308 11244 11336
rect 10744 11296 10750 11308
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12250 11336 12256 11348
rect 12023 11308 12256 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 13357 11339 13415 11345
rect 13357 11336 13369 11339
rect 12860 11308 13369 11336
rect 12860 11296 12866 11308
rect 13357 11305 13369 11308
rect 13403 11305 13415 11339
rect 13357 11299 13415 11305
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 13538 11228 13544 11280
rect 13596 11268 13602 11280
rect 14461 11271 14519 11277
rect 14461 11268 14473 11271
rect 13596 11240 14473 11268
rect 13596 11228 13602 11240
rect 14461 11237 14473 11240
rect 14507 11237 14519 11271
rect 14461 11231 14519 11237
rect 13814 11200 13820 11212
rect 6512 11172 9812 11200
rect 13648 11172 13820 11200
rect 6512 11160 6518 11172
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 5810 11132 5816 11144
rect 3936 11104 5816 11132
rect 3936 11092 3942 11104
rect 5810 11092 5816 11104
rect 5868 11141 5874 11144
rect 5868 11135 5929 11141
rect 5868 11101 5883 11135
rect 5917 11101 5929 11135
rect 5868 11095 5929 11101
rect 5868 11092 5874 11095
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 10965 11135 11023 11141
rect 10965 11132 10977 11135
rect 10468 11104 10977 11132
rect 10468 11092 10474 11104
rect 10965 11101 10977 11104
rect 11011 11101 11023 11135
rect 11238 11132 11244 11144
rect 11199 11104 11244 11132
rect 10965 11095 11023 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 12066 11092 12072 11144
rect 12124 11132 12130 11144
rect 12618 11141 12624 11144
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 12124 11104 12357 11132
rect 12124 11092 12130 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12587 11135 12624 11141
rect 12587 11101 12599 11135
rect 12587 11095 12624 11101
rect 12618 11092 12624 11095
rect 12676 11092 12682 11144
rect 8570 11024 8576 11076
rect 8628 11064 8634 11076
rect 13648 11064 13676 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14090 11132 14096 11144
rect 13771 11104 14096 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14090 11092 14096 11104
rect 14148 11092 14154 11144
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11132 14335 11135
rect 15194 11132 15200 11144
rect 14323 11104 15200 11132
rect 14323 11101 14335 11104
rect 14277 11095 14335 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 8628 11036 13676 11064
rect 8628 11024 8634 11036
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12342 10996 12348 11008
rect 11756 10968 12348 10996
rect 11756 10956 11762 10968
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13906 10996 13912 11008
rect 12768 10968 13912 10996
rect 12768 10956 12774 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 1104 10906 14971 10928
rect 1104 10854 4376 10906
rect 4428 10854 4440 10906
rect 4492 10854 4504 10906
rect 4556 10854 4568 10906
rect 4620 10854 4632 10906
rect 4684 10854 7803 10906
rect 7855 10854 7867 10906
rect 7919 10854 7931 10906
rect 7983 10854 7995 10906
rect 8047 10854 8059 10906
rect 8111 10854 11230 10906
rect 11282 10854 11294 10906
rect 11346 10854 11358 10906
rect 11410 10854 11422 10906
rect 11474 10854 11486 10906
rect 11538 10854 14657 10906
rect 14709 10854 14721 10906
rect 14773 10854 14785 10906
rect 14837 10854 14849 10906
rect 14901 10854 14913 10906
rect 14965 10854 14971 10906
rect 1104 10832 14971 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1544 10764 1961 10792
rect 1544 10752 1550 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 12618 10792 12624 10804
rect 1949 10755 2007 10761
rect 2148 10764 12624 10792
rect 1486 10616 1492 10668
rect 1544 10616 1550 10668
rect 2148 10665 2176 10764
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 13722 10752 13728 10804
rect 13780 10792 13786 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 13780 10764 13829 10792
rect 13780 10752 13786 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 14461 10795 14519 10801
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 15838 10792 15844 10804
rect 14507 10764 15844 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 15838 10752 15844 10764
rect 15896 10752 15902 10804
rect 4246 10684 4252 10736
rect 4304 10684 4310 10736
rect 5350 10684 5356 10736
rect 5408 10724 5414 10736
rect 14182 10724 14188 10736
rect 5408 10696 11744 10724
rect 5408 10684 5414 10696
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 4264 10656 4292 10684
rect 6822 10665 6828 10668
rect 4491 10659 4549 10665
rect 4491 10656 4503 10659
rect 4264 10628 4503 10656
rect 2133 10619 2191 10625
rect 4491 10625 4503 10628
rect 4537 10625 4549 10659
rect 4491 10619 4549 10625
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6791 10659 6828 10665
rect 6791 10625 6803 10659
rect 6791 10619 6828 10625
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10557 4307 10591
rect 5920 10588 5948 10619
rect 6822 10616 6828 10619
rect 6880 10616 6886 10668
rect 10287 10659 10345 10665
rect 10287 10656 10299 10659
rect 8496 10628 10299 10656
rect 6362 10588 6368 10600
rect 5920 10560 6368 10588
rect 4249 10551 4307 10557
rect 4264 10520 4292 10551
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 5534 10520 5540 10532
rect 4264 10492 4384 10520
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 900 10424 1593 10452
rect 900 10412 906 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 4356 10452 4384 10492
rect 4908 10492 5540 10520
rect 4908 10452 4936 10492
rect 5534 10480 5540 10492
rect 5592 10520 5598 10532
rect 6564 10520 6592 10551
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7892 10560 8217 10588
rect 7892 10548 7898 10560
rect 8205 10557 8217 10560
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 5592 10492 5864 10520
rect 5592 10480 5598 10492
rect 4356 10424 4936 10452
rect 1581 10415 1639 10421
rect 5258 10412 5264 10464
rect 5316 10412 5322 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5721 10455 5779 10461
rect 5721 10452 5733 10455
rect 5500 10424 5733 10452
rect 5500 10412 5506 10424
rect 5721 10421 5733 10424
rect 5767 10421 5779 10455
rect 5836 10452 5864 10492
rect 6288 10492 6592 10520
rect 6288 10452 6316 10492
rect 8496 10464 8524 10628
rect 10287 10625 10299 10628
rect 10333 10656 10345 10659
rect 10333 10628 11652 10656
rect 10333 10625 10345 10628
rect 10287 10619 10345 10625
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9732 10560 10057 10588
rect 9732 10548 9738 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 11624 10520 11652 10628
rect 11716 10588 11744 10696
rect 12406 10696 14188 10724
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10656 11943 10659
rect 12406 10656 12434 10696
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 11931 10628 12434 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12526 10616 12532 10668
rect 12584 10656 12590 10668
rect 13047 10659 13105 10665
rect 13047 10656 13059 10659
rect 12584 10628 13059 10656
rect 12584 10616 12590 10628
rect 13047 10625 13059 10628
rect 13093 10625 13105 10659
rect 13047 10619 13105 10625
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 15102 10656 15108 10668
rect 14323 10628 15108 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 11974 10588 11980 10600
rect 11716 10560 11980 10588
rect 11974 10548 11980 10560
rect 12032 10588 12038 10600
rect 12161 10591 12219 10597
rect 12161 10588 12173 10591
rect 12032 10560 12173 10588
rect 12032 10548 12038 10560
rect 12161 10557 12173 10560
rect 12207 10557 12219 10591
rect 12161 10551 12219 10557
rect 12805 10591 12863 10597
rect 12805 10557 12817 10591
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12250 10520 12256 10532
rect 11624 10492 12256 10520
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 5836 10424 6316 10452
rect 5721 10415 5779 10421
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 7374 10452 7380 10464
rect 6420 10424 7380 10452
rect 6420 10412 6426 10424
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 8110 10452 8116 10464
rect 7607 10424 8116 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8478 10412 8484 10464
rect 8536 10412 8542 10464
rect 11057 10455 11115 10461
rect 11057 10421 11069 10455
rect 11103 10452 11115 10455
rect 11606 10452 11612 10464
rect 11103 10424 11612 10452
rect 11103 10421 11115 10424
rect 11057 10415 11115 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 12066 10412 12072 10464
rect 12124 10452 12130 10464
rect 12820 10452 12848 10551
rect 12124 10424 12848 10452
rect 12124 10412 12130 10424
rect 1104 10362 14812 10384
rect 1104 10310 2663 10362
rect 2715 10310 2727 10362
rect 2779 10310 2791 10362
rect 2843 10310 2855 10362
rect 2907 10310 2919 10362
rect 2971 10310 6090 10362
rect 6142 10310 6154 10362
rect 6206 10310 6218 10362
rect 6270 10310 6282 10362
rect 6334 10310 6346 10362
rect 6398 10310 9517 10362
rect 9569 10310 9581 10362
rect 9633 10310 9645 10362
rect 9697 10310 9709 10362
rect 9761 10310 9773 10362
rect 9825 10310 12944 10362
rect 12996 10310 13008 10362
rect 13060 10310 13072 10362
rect 13124 10310 13136 10362
rect 13188 10310 13200 10362
rect 13252 10310 14812 10362
rect 1104 10288 14812 10310
rect 8478 10248 8484 10260
rect 2746 10220 8484 10248
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1397 10047 1455 10053
rect 1397 10044 1409 10047
rect 1360 10016 1409 10044
rect 1360 10004 1366 10016
rect 1397 10013 1409 10016
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1412 9976 1440 10007
rect 1578 10004 1584 10056
rect 1636 10044 1642 10056
rect 1671 10047 1729 10053
rect 1671 10044 1683 10047
rect 1636 10016 1683 10044
rect 1636 10004 1642 10016
rect 1671 10013 1683 10016
rect 1717 10013 1729 10047
rect 1671 10007 1729 10013
rect 1686 9976 1714 10007
rect 2746 9976 2774 10220
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 12066 10248 12072 10260
rect 9456 10220 9996 10248
rect 9456 10208 9462 10220
rect 5258 10140 5264 10192
rect 5316 10140 5322 10192
rect 5442 10140 5448 10192
rect 5500 10140 5506 10192
rect 6549 10183 6607 10189
rect 6549 10149 6561 10183
rect 6595 10180 6607 10183
rect 7561 10183 7619 10189
rect 7561 10180 7573 10183
rect 6595 10152 7573 10180
rect 6595 10149 6607 10152
rect 6549 10143 6607 10149
rect 7561 10149 7573 10152
rect 7607 10180 7619 10183
rect 7650 10180 7656 10192
rect 7607 10152 7656 10180
rect 7607 10149 7619 10152
rect 7561 10143 7619 10149
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 9416 10180 9444 10208
rect 9324 10152 9444 10180
rect 5074 10112 5080 10124
rect 5000 10084 5080 10112
rect 5000 10053 5028 10084
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 5276 10112 5304 10140
rect 5132 10084 5304 10112
rect 5132 10072 5138 10084
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10013 5227 10047
rect 5169 10007 5227 10013
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5460 10044 5488 10140
rect 5534 10072 5540 10124
rect 5592 10072 5598 10124
rect 7101 10115 7159 10121
rect 7101 10081 7113 10115
rect 7147 10112 7159 10115
rect 7466 10112 7472 10124
rect 7147 10084 7472 10112
rect 7147 10081 7159 10084
rect 7101 10075 7159 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7834 10072 7840 10124
rect 7892 10072 7898 10124
rect 9324 10121 9352 10152
rect 7975 10115 8033 10121
rect 7975 10081 7987 10115
rect 8021 10112 8033 10115
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8021 10084 9137 10112
rect 8021 10081 8033 10084
rect 7975 10075 8033 10081
rect 9125 10081 9137 10084
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10081 9367 10115
rect 9968 10112 9996 10220
rect 10428 10220 12072 10248
rect 10428 10192 10456 10220
rect 12066 10208 12072 10220
rect 12124 10208 12130 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13262 10248 13268 10260
rect 13127 10220 13268 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13262 10208 13268 10220
rect 13320 10208 13326 10260
rect 13354 10208 13360 10260
rect 13412 10248 13418 10260
rect 13633 10251 13691 10257
rect 13633 10248 13645 10251
rect 13412 10220 13645 10248
rect 13412 10208 13418 10220
rect 13633 10217 13645 10220
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 13906 10208 13912 10260
rect 13964 10208 13970 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14369 10251 14427 10257
rect 14369 10248 14381 10251
rect 14148 10220 14381 10248
rect 14148 10208 14154 10220
rect 14369 10217 14381 10220
rect 14415 10217 14427 10251
rect 14369 10211 14427 10217
rect 10410 10140 10416 10192
rect 10468 10140 10474 10192
rect 12084 10121 12112 10208
rect 13814 10180 13820 10192
rect 12728 10152 13820 10180
rect 12069 10115 12127 10121
rect 9968 10084 10548 10112
rect 9309 10075 9367 10081
rect 10520 10056 10548 10084
rect 12069 10081 12081 10115
rect 12115 10081 12127 10115
rect 12069 10075 12127 10081
rect 5307 10016 5488 10044
rect 5811 10047 5869 10053
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5811 10013 5823 10047
rect 5857 10044 5869 10047
rect 6546 10044 6552 10056
rect 5857 10016 6552 10044
rect 5857 10013 5869 10016
rect 5811 10007 5869 10013
rect 1412 9948 1624 9976
rect 1686 9948 2774 9976
rect 5184 9976 5212 10007
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 5626 9976 5632 9988
rect 5184 9948 5632 9976
rect 1596 9920 1624 9948
rect 5626 9936 5632 9948
rect 5684 9936 5690 9988
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6932 9976 6960 10007
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9583 10047 9641 10053
rect 9583 10044 9595 10047
rect 9272 10016 9595 10044
rect 9272 10004 9278 10016
rect 9583 10013 9595 10016
rect 9629 10013 9641 10047
rect 9583 10007 9641 10013
rect 10502 10004 10508 10056
rect 10560 10044 10566 10056
rect 10689 10047 10747 10053
rect 10689 10044 10701 10047
rect 10560 10016 10701 10044
rect 10560 10004 10566 10016
rect 10689 10013 10701 10016
rect 10735 10013 10747 10047
rect 10689 10007 10747 10013
rect 10963 10047 11021 10053
rect 10963 10013 10975 10047
rect 11009 10044 11021 10047
rect 11054 10044 11060 10056
rect 11009 10016 11060 10044
rect 11009 10013 11021 10016
rect 10963 10007 11021 10013
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 12343 10047 12401 10053
rect 12343 10044 12355 10047
rect 12308 10016 12355 10044
rect 12308 10004 12314 10016
rect 12343 10013 12355 10016
rect 12389 10013 12401 10047
rect 12343 10007 12401 10013
rect 12728 9976 12756 10152
rect 13814 10140 13820 10152
rect 13872 10140 13878 10192
rect 14642 10112 14648 10124
rect 13464 10084 14648 10112
rect 13464 10053 13492 10084
rect 14642 10072 14648 10084
rect 14700 10072 14706 10124
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 15194 10044 15200 10056
rect 13771 10016 15200 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 15194 10004 15200 10016
rect 15252 10004 15258 10056
rect 5960 9948 6960 9976
rect 10336 9948 12756 9976
rect 14277 9979 14335 9985
rect 5960 9936 5966 9948
rect 1578 9868 1584 9920
rect 1636 9868 1642 9920
rect 2406 9868 2412 9920
rect 2464 9868 2470 9920
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5258 9908 5264 9920
rect 5215 9880 5264 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5350 9868 5356 9920
rect 5408 9868 5414 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 10336 9917 10364 9948
rect 14277 9945 14289 9979
rect 14323 9976 14335 9979
rect 15102 9976 15108 9988
rect 14323 9948 15108 9976
rect 14323 9945 14335 9948
rect 14277 9939 14335 9945
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 7524 9880 8769 9908
rect 7524 9868 7530 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 10321 9911 10379 9917
rect 10321 9877 10333 9911
rect 10367 9877 10379 9911
rect 10321 9871 10379 9877
rect 11701 9911 11759 9917
rect 11701 9877 11713 9911
rect 11747 9908 11759 9911
rect 13262 9908 13268 9920
rect 11747 9880 13268 9908
rect 11747 9877 11759 9880
rect 11701 9871 11759 9877
rect 13262 9868 13268 9880
rect 13320 9868 13326 9920
rect 1104 9818 14971 9840
rect 1104 9766 4376 9818
rect 4428 9766 4440 9818
rect 4492 9766 4504 9818
rect 4556 9766 4568 9818
rect 4620 9766 4632 9818
rect 4684 9766 7803 9818
rect 7855 9766 7867 9818
rect 7919 9766 7931 9818
rect 7983 9766 7995 9818
rect 8047 9766 8059 9818
rect 8111 9766 11230 9818
rect 11282 9766 11294 9818
rect 11346 9766 11358 9818
rect 11410 9766 11422 9818
rect 11474 9766 11486 9818
rect 11538 9766 14657 9818
rect 14709 9766 14721 9818
rect 14773 9766 14785 9818
rect 14837 9766 14849 9818
rect 14901 9766 14913 9818
rect 14965 9766 14971 9818
rect 1104 9744 14971 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 1673 9707 1731 9713
rect 1673 9704 1685 9707
rect 1544 9676 1685 9704
rect 1544 9664 1550 9676
rect 1673 9673 1685 9676
rect 1719 9673 1731 9707
rect 1673 9667 1731 9673
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9673 2099 9707
rect 2041 9667 2099 9673
rect 934 9596 940 9648
rect 992 9636 998 9648
rect 2056 9636 2084 9667
rect 5074 9664 5080 9716
rect 5132 9664 5138 9716
rect 5626 9664 5632 9716
rect 5684 9704 5690 9716
rect 5905 9707 5963 9713
rect 5905 9704 5917 9707
rect 5684 9676 5917 9704
rect 5684 9664 5690 9676
rect 5905 9673 5917 9676
rect 5951 9673 5963 9707
rect 7466 9704 7472 9716
rect 5905 9667 5963 9673
rect 7208 9676 7472 9704
rect 4154 9636 4160 9648
rect 992 9608 1900 9636
rect 2056 9608 4160 9636
rect 992 9596 998 9608
rect 1872 9577 1900 9608
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9537 1639 9571
rect 1581 9531 1639 9537
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2406 9568 2412 9580
rect 2363 9540 2412 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 1596 9432 1624 9531
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 5092 9577 5120 9664
rect 5350 9596 5356 9648
rect 5408 9596 5414 9648
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5368 9568 5396 9596
rect 5215 9540 5396 9568
rect 6089 9571 6147 9577
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 7208 9568 7236 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10410 9704 10416 9716
rect 10008 9676 10416 9704
rect 10008 9664 10014 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 11514 9704 11520 9716
rect 10744 9676 11520 9704
rect 10744 9664 10750 9676
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 13538 9704 13544 9716
rect 12492 9676 13544 9704
rect 12492 9664 12498 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 14090 9664 14096 9716
rect 14148 9704 14154 9716
rect 15378 9704 15384 9716
rect 14148 9676 15384 9704
rect 14148 9664 14154 9676
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 12710 9636 12716 9648
rect 12360 9608 12716 9636
rect 6135 9540 7236 9568
rect 7300 9540 7512 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 5258 9460 5264 9512
rect 5316 9500 5322 9512
rect 7300 9509 7328 9540
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 5316 9472 5365 9500
rect 5316 9460 5322 9472
rect 5353 9469 5365 9472
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 7101 9503 7159 9509
rect 7101 9469 7113 9503
rect 7147 9469 7159 9503
rect 7101 9463 7159 9469
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7285 9463 7343 9469
rect 6546 9432 6552 9444
rect 1596 9404 6552 9432
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 5261 9367 5319 9373
rect 5261 9364 5273 9367
rect 4028 9336 5273 9364
rect 4028 9324 4034 9336
rect 5261 9333 5273 9336
rect 5307 9333 5319 9367
rect 7116 9364 7144 9463
rect 7374 9460 7380 9512
rect 7432 9460 7438 9512
rect 7282 9364 7288 9376
rect 7116 9336 7288 9364
rect 5261 9327 5319 9333
rect 7282 9324 7288 9336
rect 7340 9324 7346 9376
rect 7392 9364 7420 9460
rect 7484 9432 7512 9540
rect 8294 9528 8300 9580
rect 8352 9528 8358 9580
rect 9677 9571 9735 9577
rect 9677 9568 9689 9571
rect 9140 9540 9689 9568
rect 9140 9512 9168 9540
rect 9677 9537 9689 9540
rect 9723 9568 9735 9571
rect 9858 9568 9864 9580
rect 9723 9540 9864 9568
rect 9723 9537 9735 9540
rect 9677 9531 9735 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10686 9528 10692 9580
rect 10744 9528 10750 9580
rect 11330 9528 11336 9580
rect 11388 9528 11394 9580
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 7708 9472 7757 9500
rect 7708 9460 7714 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8018 9460 8024 9512
rect 8076 9460 8082 9512
rect 8202 9509 8208 9512
rect 8159 9503 8208 9509
rect 8159 9469 8171 9503
rect 8205 9469 8208 9503
rect 8159 9463 8208 9469
rect 8202 9460 8208 9463
rect 8260 9500 8266 9512
rect 9122 9500 9128 9512
rect 8260 9472 9128 9500
rect 8260 9460 8266 9472
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 9493 9503 9551 9509
rect 9493 9500 9505 9503
rect 9456 9472 9505 9500
rect 9456 9460 9462 9472
rect 9493 9469 9505 9472
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 10226 9460 10232 9512
rect 10284 9500 10290 9512
rect 10413 9503 10471 9509
rect 10413 9500 10425 9503
rect 10284 9472 10425 9500
rect 10284 9460 10290 9472
rect 10413 9469 10425 9472
rect 10459 9469 10471 9503
rect 10413 9463 10471 9469
rect 10502 9460 10508 9512
rect 10560 9509 10566 9512
rect 10560 9503 10588 9509
rect 10576 9469 10588 9503
rect 10560 9463 10588 9469
rect 10560 9460 10566 9463
rect 7834 9432 7840 9444
rect 7484 9404 7840 9432
rect 7834 9392 7840 9404
rect 7892 9392 7898 9444
rect 10134 9392 10140 9444
rect 10192 9392 10198 9444
rect 11146 9392 11152 9444
rect 11204 9392 11210 9444
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 11808 9432 11836 9531
rect 11974 9528 11980 9580
rect 12032 9528 12038 9580
rect 12360 9577 12388 9608
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 14461 9639 14519 9645
rect 14461 9636 14473 9639
rect 14424 9608 14473 9636
rect 14424 9596 14430 9608
rect 14461 9605 14473 9608
rect 14507 9605 14519 9639
rect 14461 9599 14519 9605
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12360 9571 12429 9577
rect 12360 9540 12383 9571
rect 12069 9531 12127 9537
rect 12371 9537 12383 9540
rect 12417 9537 12429 9571
rect 12371 9531 12429 9537
rect 11992 9441 12020 9528
rect 12084 9444 12112 9531
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12621 9571 12679 9577
rect 12621 9568 12633 9571
rect 12584 9540 12633 9568
rect 12584 9528 12590 9540
rect 12621 9537 12633 9540
rect 12667 9537 12679 9571
rect 12621 9531 12679 9537
rect 13538 9528 13544 9580
rect 13596 9528 13602 9580
rect 13814 9528 13820 9580
rect 13872 9528 13878 9580
rect 12802 9509 12808 9512
rect 12759 9503 12808 9509
rect 12759 9469 12771 9503
rect 12805 9469 12808 9503
rect 12759 9463 12808 9469
rect 12802 9460 12808 9463
rect 12860 9460 12866 9512
rect 13658 9503 13716 9509
rect 13658 9500 13670 9503
rect 12894 9472 13670 9500
rect 11756 9404 11836 9432
rect 11977 9435 12035 9441
rect 11756 9392 11762 9404
rect 11977 9401 11989 9435
rect 12023 9401 12035 9435
rect 11977 9395 12035 9401
rect 12066 9392 12072 9444
rect 12124 9392 12130 9444
rect 12894 9432 12922 9472
rect 13658 9469 13670 9472
rect 13704 9469 13716 9503
rect 13658 9463 13716 9469
rect 12544 9404 12922 9432
rect 13265 9435 13323 9441
rect 8941 9367 8999 9373
rect 8941 9364 8953 9367
rect 7392 9336 8953 9364
rect 8941 9333 8953 9336
rect 8987 9333 8999 9367
rect 8941 9327 8999 9333
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 11164 9364 11192 9392
rect 12253 9367 12311 9373
rect 12253 9364 12265 9367
rect 10560 9336 12265 9364
rect 10560 9324 10566 9336
rect 12253 9333 12265 9336
rect 12299 9333 12311 9367
rect 12253 9327 12311 9333
rect 12434 9324 12440 9376
rect 12492 9364 12498 9376
rect 12544 9373 12572 9404
rect 13265 9401 13277 9435
rect 13311 9401 13323 9435
rect 13265 9395 13323 9401
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12492 9336 12541 9364
rect 12492 9324 12498 9336
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 13280 9364 13308 9395
rect 13814 9364 13820 9376
rect 13280 9336 13820 9364
rect 12529 9327 12587 9333
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 1104 9274 14812 9296
rect 1104 9222 2663 9274
rect 2715 9222 2727 9274
rect 2779 9222 2791 9274
rect 2843 9222 2855 9274
rect 2907 9222 2919 9274
rect 2971 9222 6090 9274
rect 6142 9222 6154 9274
rect 6206 9222 6218 9274
rect 6270 9222 6282 9274
rect 6334 9222 6346 9274
rect 6398 9222 9517 9274
rect 9569 9222 9581 9274
rect 9633 9222 9645 9274
rect 9697 9222 9709 9274
rect 9761 9222 9773 9274
rect 9825 9222 12944 9274
rect 12996 9222 13008 9274
rect 13060 9222 13072 9274
rect 13124 9222 13136 9274
rect 13188 9222 13200 9274
rect 13252 9222 14812 9274
rect 1104 9200 14812 9222
rect 1486 9120 1492 9172
rect 1544 9120 1550 9172
rect 10134 9160 10140 9172
rect 9600 9132 10140 9160
rect 1504 9092 1532 9120
rect 9600 9101 9628 9132
rect 10134 9120 10140 9132
rect 10192 9160 10198 9172
rect 10192 9132 11560 9160
rect 10192 9120 10198 9132
rect 11532 9101 11560 9132
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 15102 9160 15108 9172
rect 12124 9132 15108 9160
rect 12124 9120 12130 9132
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 1412 9064 1532 9092
rect 9585 9095 9643 9101
rect 1412 9033 1440 9064
rect 9585 9061 9597 9095
rect 9631 9061 9643 9095
rect 9585 9055 9643 9061
rect 11517 9095 11575 9101
rect 11517 9061 11529 9095
rect 11563 9061 11575 9095
rect 12986 9092 12992 9104
rect 11517 9055 11575 9061
rect 12452 9064 12992 9092
rect 12452 9036 12480 9064
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 7282 8984 7288 9036
rect 7340 9024 7346 9036
rect 8386 9024 8392 9036
rect 7340 8996 8392 9024
rect 7340 8984 7346 8996
rect 8386 8984 8392 8996
rect 8444 9024 8450 9036
rect 9858 9024 9864 9036
rect 8444 8996 9864 9024
rect 8444 8984 8450 8996
rect 9858 8984 9864 8996
rect 9916 8984 9922 9036
rect 10137 9027 10195 9033
rect 10137 8993 10149 9027
rect 10183 9024 10195 9027
rect 10318 9024 10324 9036
rect 10183 8996 10324 9024
rect 10183 8993 10195 8996
rect 10137 8987 10195 8993
rect 10318 8984 10324 8996
rect 10376 9024 10382 9036
rect 10686 9024 10692 9036
rect 10376 8996 10692 9024
rect 10376 8984 10382 8996
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 10873 9027 10931 9033
rect 10873 8993 10885 9027
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 1655 8929 1713 8935
rect 1655 8926 1667 8929
rect 1394 8848 1400 8900
rect 1452 8888 1458 8900
rect 1596 8898 1667 8926
rect 1596 8888 1624 8898
rect 1655 8895 1667 8898
rect 1701 8895 1713 8929
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 8018 8956 8024 8968
rect 7524 8928 8024 8956
rect 7524 8916 7530 8928
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8904 8928 8953 8956
rect 8904 8916 8910 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 1655 8889 1713 8895
rect 1452 8860 1624 8888
rect 1452 8848 1458 8860
rect 7834 8848 7840 8900
rect 7892 8848 7898 8900
rect 9030 8848 9036 8900
rect 9088 8888 9094 8900
rect 9140 8888 9168 8919
rect 9950 8916 9956 8968
rect 10008 8965 10014 8968
rect 10008 8959 10036 8965
rect 10024 8925 10036 8959
rect 10888 8956 10916 8987
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 11793 9027 11851 9033
rect 11793 9024 11805 9027
rect 11020 8996 11805 9024
rect 11020 8984 11026 8996
rect 11793 8993 11805 8996
rect 11839 8993 11851 9027
rect 11793 8987 11851 8993
rect 12434 8984 12440 9036
rect 12492 8984 12498 9036
rect 14366 9024 14372 9036
rect 12820 8996 14372 9024
rect 10008 8919 10036 8925
rect 10704 8928 10916 8956
rect 11057 8959 11115 8965
rect 10008 8916 10014 8919
rect 10704 8900 10732 8928
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11238 8956 11244 8968
rect 11103 8928 11244 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11974 8965 11980 8968
rect 11931 8959 11980 8965
rect 11931 8925 11943 8959
rect 11977 8925 11980 8959
rect 11931 8919 11980 8925
rect 11974 8916 11980 8919
rect 12032 8916 12038 8968
rect 12066 8916 12072 8968
rect 12124 8916 12130 8968
rect 12820 8965 12848 8996
rect 14366 8984 14372 8996
rect 14424 8984 14430 9036
rect 14458 8984 14464 9036
rect 14516 8984 14522 9036
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13081 8959 13139 8965
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 9088 8860 9168 8888
rect 9088 8848 9094 8860
rect 10686 8848 10692 8900
rect 10744 8848 10750 8900
rect 10781 8891 10839 8897
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 10870 8888 10876 8900
rect 10827 8860 10876 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8888 12771 8891
rect 12894 8888 12900 8900
rect 12759 8860 12900 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 13096 8888 13124 8919
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 14274 8916 14280 8968
rect 14332 8916 14338 8968
rect 14476 8888 14504 8984
rect 13096 8860 14504 8888
rect 2406 8780 2412 8832
rect 2464 8780 2470 8832
rect 7852 8820 7880 8848
rect 9306 8820 9312 8832
rect 7852 8792 9312 8820
rect 9306 8780 9312 8792
rect 9364 8820 9370 8832
rect 9950 8820 9956 8832
rect 9364 8792 9956 8820
rect 9364 8780 9370 8792
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 10226 8780 10232 8832
rect 10284 8820 10290 8832
rect 12526 8820 12532 8832
rect 10284 8792 12532 8820
rect 10284 8780 10290 8792
rect 12526 8780 12532 8792
rect 12584 8820 12590 8832
rect 12989 8823 13047 8829
rect 12989 8820 13001 8823
rect 12584 8792 13001 8820
rect 12584 8780 12590 8792
rect 12989 8789 13001 8792
rect 13035 8789 13047 8823
rect 12989 8783 13047 8789
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 13504 8792 14473 8820
rect 13504 8780 13510 8792
rect 14461 8789 14473 8792
rect 14507 8789 14519 8823
rect 14461 8783 14519 8789
rect 1104 8730 14971 8752
rect 1104 8678 4376 8730
rect 4428 8678 4440 8730
rect 4492 8678 4504 8730
rect 4556 8678 4568 8730
rect 4620 8678 4632 8730
rect 4684 8678 7803 8730
rect 7855 8678 7867 8730
rect 7919 8678 7931 8730
rect 7983 8678 7995 8730
rect 8047 8678 8059 8730
rect 8111 8678 11230 8730
rect 11282 8678 11294 8730
rect 11346 8678 11358 8730
rect 11410 8678 11422 8730
rect 11474 8678 11486 8730
rect 11538 8678 14657 8730
rect 14709 8678 14721 8730
rect 14773 8678 14785 8730
rect 14837 8678 14849 8730
rect 14901 8678 14913 8730
rect 14965 8678 14971 8730
rect 1104 8656 14971 8678
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 6454 8616 6460 8628
rect 5184 8588 6460 8616
rect 1673 8551 1731 8557
rect 1673 8517 1685 8551
rect 1719 8548 1731 8551
rect 2148 8548 2176 8576
rect 1719 8520 2176 8548
rect 1719 8517 1731 8520
rect 1673 8511 1731 8517
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8480 2375 8483
rect 2424 8480 2452 8576
rect 4982 8508 4988 8560
rect 5040 8508 5046 8560
rect 5184 8519 5212 8588
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6546 8576 6552 8628
rect 6604 8616 6610 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 6604 8588 6653 8616
rect 6604 8576 6610 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10226 8616 10232 8628
rect 10008 8588 10232 8616
rect 10008 8576 10014 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 10928 8588 11468 8616
rect 10928 8576 10934 8588
rect 11440 8548 11468 8588
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 12768 8588 13369 8616
rect 12768 8576 12774 8588
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 14093 8619 14151 8625
rect 14093 8616 14105 8619
rect 13596 8588 14105 8616
rect 13596 8576 13602 8588
rect 14093 8585 14105 8588
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 5151 8513 5212 8519
rect 2363 8452 2452 8480
rect 4893 8483 4951 8489
rect 2363 8449 2375 8452
rect 2317 8443 2375 8449
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5000 8480 5028 8508
rect 4939 8452 5028 8480
rect 5151 8479 5163 8513
rect 5197 8482 5212 8513
rect 6380 8520 7052 8548
rect 11440 8520 11560 8548
rect 6380 8489 6408 8520
rect 6365 8483 6423 8489
rect 5197 8479 5209 8482
rect 6365 8480 6377 8483
rect 5151 8473 5209 8479
rect 5920 8452 6377 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 1854 8304 1860 8356
rect 1912 8304 1918 8356
rect 5920 8353 5948 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 7024 8489 7052 8520
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7558 8440 7564 8492
rect 7616 8480 7622 8492
rect 9401 8483 9459 8489
rect 9401 8480 9413 8483
rect 7616 8452 9413 8480
rect 7616 8440 7622 8452
rect 9401 8449 9413 8452
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 10410 8440 10416 8492
rect 10468 8489 10474 8492
rect 10468 8483 10496 8489
rect 10484 8449 10496 8483
rect 10468 8443 10496 8449
rect 10468 8440 10474 8443
rect 10594 8440 10600 8492
rect 10652 8440 10658 8492
rect 11241 8483 11299 8489
rect 11241 8449 11253 8483
rect 11287 8480 11299 8483
rect 11422 8480 11428 8492
rect 11287 8452 11428 8480
rect 11287 8449 11299 8452
rect 11241 8443 11299 8449
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11532 8489 11560 8520
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 12437 8483 12495 8489
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6687 8384 7113 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 8570 8372 8576 8424
rect 8628 8372 8634 8424
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9674 8412 9680 8424
rect 9631 8384 9680 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6503 8316 6837 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 9600 8344 9628 8375
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9784 8412 9812 8440
rect 10321 8415 10379 8421
rect 10321 8412 10333 8415
rect 9784 8384 10333 8412
rect 10321 8381 10333 8384
rect 10367 8381 10379 8415
rect 10321 8375 10379 8381
rect 11606 8372 11612 8424
rect 11664 8372 11670 8424
rect 11698 8372 11704 8424
rect 11756 8372 11762 8424
rect 12161 8415 12219 8421
rect 12161 8381 12173 8415
rect 12207 8381 12219 8415
rect 12452 8412 12480 8443
rect 12526 8440 12532 8492
rect 12584 8489 12590 8492
rect 12584 8483 12612 8489
rect 12600 8449 12612 8483
rect 12584 8443 12612 8449
rect 12584 8440 12590 8443
rect 13722 8440 13728 8492
rect 13780 8480 13786 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13780 8452 13921 8480
rect 13780 8440 13786 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14274 8440 14280 8492
rect 14332 8440 14338 8492
rect 12161 8375 12219 8381
rect 12268 8384 12480 8412
rect 7524 8316 9628 8344
rect 7524 8304 7530 8316
rect 10042 8304 10048 8356
rect 10100 8353 10106 8356
rect 10100 8344 10109 8353
rect 10100 8316 10145 8344
rect 10100 8307 10109 8316
rect 10100 8304 10106 8307
rect 11422 8304 11428 8356
rect 11480 8344 11486 8356
rect 11624 8344 11652 8372
rect 12176 8344 12204 8375
rect 11480 8316 11560 8344
rect 11624 8316 12204 8344
rect 11480 8304 11486 8316
rect 2130 8236 2136 8288
rect 2188 8236 2194 8288
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8481 8279 8539 8285
rect 8481 8276 8493 8279
rect 7984 8248 8493 8276
rect 7984 8236 7990 8248
rect 8481 8245 8493 8248
rect 8527 8245 8539 8279
rect 8481 8239 8539 8245
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 11146 8276 11152 8288
rect 10468 8248 11152 8276
rect 10468 8236 10474 8248
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 11532 8276 11560 8316
rect 11606 8276 11612 8288
rect 11532 8248 11612 8276
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 12268 8276 12296 8384
rect 12710 8372 12716 8424
rect 12768 8372 12774 8424
rect 13538 8372 13544 8424
rect 13596 8412 13602 8424
rect 14090 8412 14096 8424
rect 13596 8384 14096 8412
rect 13596 8372 13602 8384
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 12894 8276 12900 8288
rect 12268 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 13354 8236 13360 8288
rect 13412 8276 13418 8288
rect 14369 8279 14427 8285
rect 14369 8276 14381 8279
rect 13412 8248 14381 8276
rect 13412 8236 13418 8248
rect 14369 8245 14381 8248
rect 14415 8245 14427 8279
rect 14369 8239 14427 8245
rect 1104 8186 14812 8208
rect 1104 8134 2663 8186
rect 2715 8134 2727 8186
rect 2779 8134 2791 8186
rect 2843 8134 2855 8186
rect 2907 8134 2919 8186
rect 2971 8134 6090 8186
rect 6142 8134 6154 8186
rect 6206 8134 6218 8186
rect 6270 8134 6282 8186
rect 6334 8134 6346 8186
rect 6398 8134 9517 8186
rect 9569 8134 9581 8186
rect 9633 8134 9645 8186
rect 9697 8134 9709 8186
rect 9761 8134 9773 8186
rect 9825 8134 12944 8186
rect 12996 8134 13008 8186
rect 13060 8134 13072 8186
rect 13124 8134 13136 8186
rect 13188 8134 13200 8186
rect 13252 8134 14812 8186
rect 1104 8112 14812 8134
rect 1578 8032 1584 8084
rect 1636 8032 1642 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6730 8072 6736 8084
rect 6411 8044 6736 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 8570 8072 8576 8084
rect 7668 8044 8576 8072
rect 6641 8007 6699 8013
rect 6641 7973 6653 8007
rect 6687 8004 6699 8007
rect 7208 8004 7236 8032
rect 6687 7976 7236 8004
rect 6687 7973 6699 7976
rect 6641 7967 6699 7973
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 7064 7908 7113 7936
rect 7064 7896 7070 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 7466 7936 7472 7948
rect 7101 7899 7159 7905
rect 7300 7908 7472 7936
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 2130 7868 2136 7880
rect 1535 7840 2136 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 6546 7828 6552 7880
rect 6604 7828 6610 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7868 6975 7871
rect 7300 7868 7328 7908
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7558 7896 7564 7948
rect 7616 7896 7622 7948
rect 7668 7936 7696 8044
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9180 8044 11284 8072
rect 9180 8032 9186 8044
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7668 7908 7849 7936
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 7926 7896 7932 7948
rect 7984 7945 7990 7948
rect 9600 7945 9628 8044
rect 11256 8016 11284 8044
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 12345 8075 12403 8081
rect 11848 8044 12020 8072
rect 11848 8032 11854 8044
rect 9950 8004 9956 8016
rect 9784 7976 9956 8004
rect 9784 7948 9812 7976
rect 9950 7964 9956 7976
rect 10008 8004 10014 8016
rect 10008 7976 10180 8004
rect 10008 7964 10014 7976
rect 7984 7939 8012 7945
rect 8000 7905 8012 7939
rect 9585 7939 9643 7945
rect 7984 7899 8012 7905
rect 8128 7908 8708 7936
rect 7984 7896 7990 7899
rect 8128 7877 8156 7908
rect 6963 7840 7328 7868
rect 8113 7871 8171 7877
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 8113 7837 8125 7871
rect 8159 7837 8171 7871
rect 8680 7868 8708 7908
rect 9585 7905 9597 7939
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 9766 7896 9772 7948
rect 9824 7896 9830 7948
rect 10042 7896 10048 7948
rect 10100 7896 10106 7948
rect 10152 7936 10180 7976
rect 11238 7964 11244 8016
rect 11296 7964 11302 8016
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 10152 7908 10333 7936
rect 10321 7905 10333 7908
rect 10367 7905 10379 7939
rect 10321 7899 10379 7905
rect 10594 7896 10600 7948
rect 10652 7896 10658 7948
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11333 7939 11391 7945
rect 11333 7936 11345 7939
rect 11204 7908 11345 7936
rect 11204 7896 11210 7908
rect 11333 7905 11345 7908
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 9122 7868 9128 7880
rect 8680 7840 9128 7868
rect 8113 7831 8171 7837
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 6730 7732 6736 7744
rect 4856 7704 6736 7732
rect 4856 7692 4862 7704
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6840 7732 6868 7831
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 9398 7828 9404 7880
rect 9456 7828 9462 7880
rect 10410 7828 10416 7880
rect 10468 7877 10474 7880
rect 10468 7871 10496 7877
rect 10484 7837 10496 7871
rect 10468 7831 10496 7837
rect 11607 7871 11665 7877
rect 11607 7837 11619 7871
rect 11653 7868 11665 7871
rect 11992 7868 12020 8044
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12710 8072 12716 8084
rect 12391 8044 12716 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 14461 8007 14519 8013
rect 14461 8004 14473 8007
rect 12952 7976 14473 8004
rect 12952 7964 12958 7976
rect 14461 7973 14473 7976
rect 14507 7973 14519 8007
rect 14461 7967 14519 7973
rect 12710 7936 12716 7948
rect 12084 7908 12716 7936
rect 12084 7880 12112 7908
rect 12710 7896 12716 7908
rect 12768 7936 12774 7948
rect 13909 7939 13967 7945
rect 13909 7936 13921 7939
rect 12768 7908 13921 7936
rect 12768 7896 12774 7908
rect 13909 7905 13921 7908
rect 13955 7905 13967 7939
rect 13909 7899 13967 7905
rect 11653 7840 12020 7868
rect 11653 7837 11665 7840
rect 11607 7831 11665 7837
rect 10468 7828 10474 7831
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 14182 7868 14188 7880
rect 12820 7840 14188 7868
rect 9030 7760 9036 7812
rect 9088 7800 9094 7812
rect 9416 7800 9444 7828
rect 12820 7809 12848 7840
rect 14182 7828 14188 7840
rect 14240 7828 14246 7880
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 12805 7803 12863 7809
rect 9088 7772 9444 7800
rect 11256 7772 12434 7800
rect 9088 7760 9094 7772
rect 11256 7741 11284 7772
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 6840 7704 8769 7732
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 8757 7695 8815 7701
rect 11241 7735 11299 7741
rect 11241 7701 11253 7735
rect 11287 7701 11299 7735
rect 12406 7732 12434 7772
rect 12805 7769 12817 7803
rect 12851 7769 12863 7803
rect 12805 7763 12863 7769
rect 13725 7803 13783 7809
rect 13725 7769 13737 7803
rect 13771 7800 13783 7803
rect 14550 7800 14556 7812
rect 13771 7772 14556 7800
rect 13771 7769 13783 7772
rect 13725 7763 13783 7769
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 12618 7732 12624 7744
rect 12406 7704 12624 7732
rect 11241 7695 11299 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12894 7692 12900 7744
rect 12952 7692 12958 7744
rect 1104 7642 14971 7664
rect 1104 7590 4376 7642
rect 4428 7590 4440 7642
rect 4492 7590 4504 7642
rect 4556 7590 4568 7642
rect 4620 7590 4632 7642
rect 4684 7590 7803 7642
rect 7855 7590 7867 7642
rect 7919 7590 7931 7642
rect 7983 7590 7995 7642
rect 8047 7590 8059 7642
rect 8111 7590 11230 7642
rect 11282 7590 11294 7642
rect 11346 7590 11358 7642
rect 11410 7590 11422 7642
rect 11474 7590 11486 7642
rect 11538 7590 14657 7642
rect 14709 7590 14721 7642
rect 14773 7590 14785 7642
rect 14837 7590 14849 7642
rect 14901 7590 14913 7642
rect 14965 7590 14971 7642
rect 1104 7568 14971 7590
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1504 7500 1961 7528
rect 1504 7469 1532 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6822 7528 6828 7540
rect 6052 7500 6828 7528
rect 6052 7488 6058 7500
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7558 7488 7564 7540
rect 7616 7488 7622 7540
rect 9582 7488 9588 7540
rect 9640 7528 9646 7540
rect 9769 7531 9827 7537
rect 9769 7528 9781 7531
rect 9640 7500 9781 7528
rect 9640 7488 9646 7500
rect 9769 7497 9781 7500
rect 9815 7497 9827 7531
rect 9769 7491 9827 7497
rect 9876 7500 10640 7528
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7429 1547 7463
rect 7190 7460 7196 7472
rect 1489 7423 1547 7429
rect 6564 7432 7196 7460
rect 2130 7352 2136 7404
rect 2188 7352 2194 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 6564 7401 6592 7432
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 5776 7364 6561 7392
rect 5776 7352 5782 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6822 7392 6828 7404
rect 6783 7364 6828 7392
rect 6549 7355 6607 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7576 7392 7604 7488
rect 9030 7401 9036 7404
rect 8987 7395 9036 7401
rect 7576 7364 8248 7392
rect 7929 7327 7987 7333
rect 7929 7293 7941 7327
rect 7975 7293 7987 7327
rect 7929 7287 7987 7293
rect 7944 7256 7972 7287
rect 8110 7284 8116 7336
rect 8168 7284 8174 7336
rect 8220 7324 8248 7364
rect 8987 7361 8999 7395
rect 9033 7361 9036 7395
rect 8987 7355 9036 7361
rect 9030 7352 9036 7355
rect 9088 7352 9094 7404
rect 9876 7392 9904 7500
rect 10612 7472 10640 7500
rect 11882 7488 11888 7540
rect 11940 7488 11946 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 13262 7528 13268 7540
rect 12400 7500 13268 7528
rect 12400 7488 12406 7500
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 14461 7531 14519 7537
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 15654 7528 15660 7540
rect 14507 7500 15660 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 9950 7420 9956 7472
rect 10008 7460 10014 7472
rect 10008 7432 10180 7460
rect 10008 7420 10014 7432
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9876 7364 10057 7392
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10152 7392 10180 7432
rect 10594 7420 10600 7472
rect 10652 7420 10658 7472
rect 10319 7395 10377 7401
rect 10319 7392 10331 7395
rect 10152 7364 10331 7392
rect 10045 7355 10103 7361
rect 10319 7361 10331 7364
rect 10365 7392 10377 7395
rect 10778 7392 10784 7404
rect 10365 7364 10784 7392
rect 10365 7361 10377 7364
rect 10319 7355 10377 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 11900 7392 11928 7488
rect 11977 7395 12035 7401
rect 11977 7392 11989 7395
rect 11900 7364 11989 7392
rect 11977 7361 11989 7364
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 8573 7327 8631 7333
rect 8573 7324 8585 7327
rect 8220 7296 8585 7324
rect 8573 7293 8585 7296
rect 8619 7293 8631 7327
rect 8849 7327 8907 7333
rect 8849 7324 8861 7327
rect 8573 7287 8631 7293
rect 8680 7296 8861 7324
rect 8202 7256 8208 7268
rect 7944 7228 8208 7256
rect 8202 7216 8208 7228
rect 8260 7216 8266 7268
rect 842 7148 848 7200
rect 900 7188 906 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 900 7160 1593 7188
rect 900 7148 906 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 8680 7188 8708 7296
rect 8849 7293 8861 7296
rect 8895 7293 8907 7327
rect 8849 7287 8907 7293
rect 9122 7284 9128 7336
rect 9180 7284 9186 7336
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7324 11759 7327
rect 11882 7324 11888 7336
rect 11747 7296 11888 7324
rect 11747 7293 11759 7296
rect 11701 7287 11759 7293
rect 11882 7284 11888 7296
rect 11940 7284 11946 7336
rect 11992 7324 12020 7355
rect 12250 7352 12256 7404
rect 12308 7392 12314 7404
rect 12621 7395 12679 7401
rect 12621 7392 12633 7395
rect 12308 7364 12633 7392
rect 12308 7352 12314 7364
rect 12621 7361 12633 7364
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 12802 7352 12808 7404
rect 12860 7352 12866 7404
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 13722 7401 13728 7404
rect 13679 7395 13728 7401
rect 13679 7361 13691 7395
rect 13725 7361 13728 7395
rect 13679 7355 13728 7361
rect 13722 7352 13728 7355
rect 13780 7352 13786 7404
rect 12710 7324 12716 7336
rect 11992 7296 12716 7324
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13814 7284 13820 7336
rect 13872 7284 13878 7336
rect 11057 7259 11115 7265
rect 11057 7225 11069 7259
rect 11103 7256 11115 7259
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 11103 7228 13277 7256
rect 11103 7225 11115 7228
rect 11057 7219 11115 7225
rect 13265 7225 13277 7228
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 10410 7188 10416 7200
rect 8680 7160 10416 7188
rect 1581 7151 1639 7157
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 14366 7188 14372 7200
rect 12584 7160 14372 7188
rect 12584 7148 12590 7160
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 1104 7098 14812 7120
rect 1104 7046 2663 7098
rect 2715 7046 2727 7098
rect 2779 7046 2791 7098
rect 2843 7046 2855 7098
rect 2907 7046 2919 7098
rect 2971 7046 6090 7098
rect 6142 7046 6154 7098
rect 6206 7046 6218 7098
rect 6270 7046 6282 7098
rect 6334 7046 6346 7098
rect 6398 7046 9517 7098
rect 9569 7046 9581 7098
rect 9633 7046 9645 7098
rect 9697 7046 9709 7098
rect 9761 7046 9773 7098
rect 9825 7046 12944 7098
rect 12996 7046 13008 7098
rect 13060 7046 13072 7098
rect 13124 7046 13136 7098
rect 13188 7046 13200 7098
rect 13252 7046 14812 7098
rect 1104 7024 14812 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2188 6956 2421 6984
rect 2188 6944 2194 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 9950 6984 9956 6996
rect 6880 6956 9956 6984
rect 6880 6944 6886 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10870 6984 10876 6996
rect 10545 6956 10876 6984
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 10042 6916 10048 6928
rect 8168 6888 8432 6916
rect 8168 6876 8174 6888
rect 1394 6740 1400 6792
rect 1452 6740 1458 6792
rect 1671 6783 1729 6789
rect 1671 6749 1683 6783
rect 1717 6780 1729 6783
rect 6914 6780 6920 6792
rect 1717 6752 6920 6780
rect 1717 6749 1729 6752
rect 1671 6743 1729 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 8404 6780 8432 6888
rect 9646 6888 10048 6916
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 9646 6848 9674 6888
rect 10042 6876 10048 6888
rect 10100 6916 10106 6928
rect 10100 6888 10456 6916
rect 10100 6876 10106 6888
rect 10428 6857 10456 6888
rect 9456 6820 9674 6848
rect 9953 6851 10011 6857
rect 9456 6808 9462 6820
rect 9953 6817 9965 6851
rect 9999 6817 10011 6851
rect 9953 6811 10011 6817
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6817 10471 6851
rect 10545 6848 10573 6956
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 14366 6944 14372 6996
rect 14424 6944 14430 6996
rect 10806 6851 10864 6857
rect 10806 6848 10818 6851
rect 10545 6820 10818 6848
rect 10413 6811 10471 6817
rect 10806 6817 10818 6820
rect 10852 6817 10864 6851
rect 10806 6811 10864 6817
rect 8404 6752 9674 6780
rect 9646 6724 9674 6752
rect 9766 6740 9772 6792
rect 9824 6740 9830 6792
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 9646 6684 9680 6724
rect 9674 6672 9680 6684
rect 9732 6712 9738 6724
rect 9876 6712 9904 6740
rect 9732 6684 9904 6712
rect 9732 6672 9738 6684
rect 9968 6656 9996 6811
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 12250 6848 12256 6860
rect 11664 6820 12256 6848
rect 11664 6808 11670 6820
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 13354 6808 13360 6860
rect 13412 6808 13418 6860
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 12802 6780 12808 6792
rect 11848 6752 12808 6780
rect 11848 6740 11854 6752
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13998 6780 14004 6792
rect 13311 6752 14004 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 11440 6684 12204 6712
rect 9950 6604 9956 6656
rect 10008 6644 10014 6656
rect 11440 6644 11468 6684
rect 10008 6616 11468 6644
rect 11609 6647 11667 6653
rect 10008 6604 10014 6616
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 12066 6644 12072 6656
rect 11655 6616 12072 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 12066 6604 12072 6616
rect 12124 6604 12130 6656
rect 12176 6644 12204 6684
rect 12526 6672 12532 6724
rect 12584 6672 12590 6724
rect 12710 6672 12716 6724
rect 12768 6672 12774 6724
rect 12728 6644 12756 6672
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 12176 6616 13645 6644
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 13906 6644 13912 6656
rect 13863 6616 13912 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 1104 6554 14971 6576
rect 1104 6502 4376 6554
rect 4428 6502 4440 6554
rect 4492 6502 4504 6554
rect 4556 6502 4568 6554
rect 4620 6502 4632 6554
rect 4684 6502 7803 6554
rect 7855 6502 7867 6554
rect 7919 6502 7931 6554
rect 7983 6502 7995 6554
rect 8047 6502 8059 6554
rect 8111 6502 11230 6554
rect 11282 6502 11294 6554
rect 11346 6502 11358 6554
rect 11410 6502 11422 6554
rect 11474 6502 11486 6554
rect 11538 6502 14657 6554
rect 14709 6502 14721 6554
rect 14773 6502 14785 6554
rect 14837 6502 14849 6554
rect 14901 6502 14913 6554
rect 14965 6502 14971 6554
rect 1104 6480 14971 6502
rect 842 6400 848 6452
rect 900 6440 906 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 900 6412 1593 6440
rect 900 6400 906 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 2317 6443 2375 6449
rect 2317 6440 2329 6443
rect 1581 6403 1639 6409
rect 1872 6412 2329 6440
rect 1489 6375 1547 6381
rect 1489 6341 1501 6375
rect 1535 6372 1547 6375
rect 1872 6372 1900 6412
rect 2317 6409 2329 6412
rect 2363 6409 2375 6443
rect 11974 6440 11980 6452
rect 2317 6403 2375 6409
rect 8864 6412 11980 6440
rect 8294 6372 8300 6384
rect 1535 6344 1900 6372
rect 2240 6344 8300 6372
rect 1535 6341 1547 6344
rect 1489 6335 1547 6341
rect 2240 6313 2268 6344
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 8864 6316 8892 6412
rect 11974 6400 11980 6412
rect 12032 6440 12038 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 12032 6412 12357 6440
rect 12032 6400 12038 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 12728 6412 12922 6440
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 12158 6372 12164 6384
rect 10744 6344 12164 6372
rect 10744 6332 10750 6344
rect 12158 6332 12164 6344
rect 12216 6332 12222 6384
rect 12728 6381 12756 6412
rect 12713 6375 12771 6381
rect 12713 6341 12725 6375
rect 12759 6341 12771 6375
rect 12894 6372 12922 6412
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 13633 6443 13691 6449
rect 13228 6412 13492 6440
rect 13228 6400 13234 6412
rect 13262 6372 13268 6384
rect 12894 6344 13268 6372
rect 12713 6335 12771 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13464 6381 13492 6412
rect 13633 6409 13645 6443
rect 13679 6440 13691 6443
rect 14458 6440 14464 6452
rect 13679 6412 14464 6440
rect 13679 6409 13691 6412
rect 13633 6403 13691 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 13449 6375 13507 6381
rect 13449 6341 13461 6375
rect 13495 6372 13507 6375
rect 13495 6344 13952 6372
rect 13495 6341 13507 6344
rect 13449 6335 13507 6341
rect 13924 6316 13952 6344
rect 2225 6307 2283 6313
rect 2225 6273 2237 6307
rect 2271 6273 2283 6307
rect 2225 6267 2283 6273
rect 2498 6264 2504 6316
rect 2556 6264 2562 6316
rect 6914 6264 6920 6316
rect 6972 6304 6978 6316
rect 7619 6307 7677 6313
rect 7619 6304 7631 6307
rect 6972 6276 7631 6304
rect 6972 6264 6978 6276
rect 7619 6273 7631 6276
rect 7665 6273 7677 6307
rect 8846 6304 8852 6316
rect 7619 6267 7677 6273
rect 8772 6276 8852 6304
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 8772 6245 8800 6276
rect 8846 6264 8852 6276
rect 8904 6264 8910 6316
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12802 6304 12808 6316
rect 12667 6276 12808 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13081 6307 13139 6313
rect 13081 6304 13093 6307
rect 13044 6276 13093 6304
rect 13044 6264 13050 6276
rect 13081 6273 13093 6276
rect 13127 6304 13139 6307
rect 13127 6276 13492 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7248 6208 7389 6236
rect 7248 6196 7254 6208
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 8757 6239 8815 6245
rect 8757 6205 8769 6239
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 9306 6196 9312 6248
rect 9364 6236 9370 6248
rect 9794 6239 9852 6245
rect 9794 6236 9806 6239
rect 9364 6208 9806 6236
rect 9364 6196 9370 6208
rect 9794 6205 9806 6208
rect 9840 6205 9852 6239
rect 9794 6199 9852 6205
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10980 6236 11008 6264
rect 9999 6208 11008 6236
rect 12348 6248 12400 6254
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 12348 6190 12400 6196
rect 9398 6128 9404 6180
rect 9456 6128 9462 6180
rect 10962 6168 10968 6180
rect 10520 6140 10968 6168
rect 2038 6060 2044 6112
rect 2096 6060 2102 6112
rect 8389 6103 8447 6109
rect 8389 6069 8401 6103
rect 8435 6100 8447 6103
rect 10318 6100 10324 6112
rect 8435 6072 10324 6100
rect 8435 6069 8447 6072
rect 8389 6063 8447 6069
rect 10318 6060 10324 6072
rect 10376 6100 10382 6112
rect 10520 6100 10548 6140
rect 10962 6128 10968 6140
rect 11020 6128 11026 6180
rect 13464 6168 13492 6276
rect 13906 6264 13912 6316
rect 13964 6264 13970 6316
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6304 14335 6307
rect 15102 6304 15108 6316
rect 14323 6276 15108 6304
rect 14323 6273 14335 6276
rect 14277 6267 14335 6273
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 14461 6171 14519 6177
rect 14461 6168 14473 6171
rect 13464 6140 14473 6168
rect 14461 6137 14473 6140
rect 14507 6137 14519 6171
rect 14461 6131 14519 6137
rect 10376 6072 10548 6100
rect 10597 6103 10655 6109
rect 10376 6060 10382 6072
rect 10597 6069 10609 6103
rect 10643 6100 10655 6103
rect 11146 6100 11152 6112
rect 10643 6072 11152 6100
rect 10643 6069 10655 6072
rect 10597 6063 10655 6069
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 1104 6010 14812 6032
rect 1104 5958 2663 6010
rect 2715 5958 2727 6010
rect 2779 5958 2791 6010
rect 2843 5958 2855 6010
rect 2907 5958 2919 6010
rect 2971 5958 6090 6010
rect 6142 5958 6154 6010
rect 6206 5958 6218 6010
rect 6270 5958 6282 6010
rect 6334 5958 6346 6010
rect 6398 5958 9517 6010
rect 9569 5958 9581 6010
rect 9633 5958 9645 6010
rect 9697 5958 9709 6010
rect 9761 5958 9773 6010
rect 9825 5958 12944 6010
rect 12996 5958 13008 6010
rect 13060 5958 13072 6010
rect 13124 5958 13136 6010
rect 13188 5958 13200 6010
rect 13252 5958 14812 6010
rect 1104 5936 14812 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 8389 5899 8447 5905
rect 8389 5865 8401 5899
rect 8435 5896 8447 5899
rect 9122 5896 9128 5908
rect 8435 5868 9128 5896
rect 8435 5865 8447 5868
rect 8389 5859 8447 5865
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 11146 5856 11152 5908
rect 11204 5896 11210 5908
rect 11204 5868 11376 5896
rect 11204 5856 11210 5868
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7248 5732 7389 5760
rect 7248 5720 7254 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7377 5723 7435 5729
rect 9766 5720 9772 5772
rect 9824 5720 9830 5772
rect 9950 5720 9956 5772
rect 10008 5720 10014 5772
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10192 5732 10425 5760
rect 10192 5720 10198 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10686 5720 10692 5772
rect 10744 5720 10750 5772
rect 10962 5720 10968 5772
rect 11020 5720 11026 5772
rect 11348 5760 11376 5868
rect 13538 5856 13544 5908
rect 13596 5856 13602 5908
rect 14366 5856 14372 5908
rect 14424 5856 14430 5908
rect 15286 5856 15292 5908
rect 15344 5856 15350 5908
rect 12066 5828 12072 5840
rect 11900 5800 12072 5828
rect 11900 5769 11928 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 12250 5788 12256 5840
rect 12308 5828 12314 5840
rect 13909 5831 13967 5837
rect 12308 5800 12480 5828
rect 12308 5788 12314 5800
rect 11885 5763 11943 5769
rect 11348 5732 11560 5760
rect 1394 5652 1400 5704
rect 1452 5692 1458 5704
rect 1452 5664 1624 5692
rect 1452 5652 1458 5664
rect 1596 5568 1624 5664
rect 1655 5665 1713 5671
rect 1655 5631 1667 5665
rect 1701 5662 1713 5665
rect 1701 5631 1716 5662
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7619 5695 7677 5701
rect 7619 5692 7631 5695
rect 6788 5664 7631 5692
rect 6788 5652 6794 5664
rect 7619 5661 7631 5664
rect 7665 5692 7677 5695
rect 8202 5692 8208 5704
rect 7665 5664 8208 5692
rect 7665 5661 7677 5664
rect 7619 5655 7677 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 10870 5701 10876 5704
rect 10827 5695 10876 5701
rect 10827 5661 10839 5695
rect 10873 5661 10876 5695
rect 10827 5655 10876 5661
rect 10870 5652 10876 5655
rect 10928 5652 10934 5704
rect 11532 5692 11560 5732
rect 11885 5729 11897 5763
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12345 5763 12403 5769
rect 12345 5760 12357 5763
rect 12032 5732 12357 5760
rect 12032 5720 12038 5732
rect 12345 5729 12357 5732
rect 12391 5729 12403 5763
rect 12452 5760 12480 5800
rect 13909 5797 13921 5831
rect 13955 5828 13967 5831
rect 15304 5828 15332 5856
rect 13955 5800 15332 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12452 5732 12633 5760
rect 12345 5723 12403 5729
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12710 5720 12716 5772
rect 12768 5769 12774 5772
rect 12768 5763 12796 5769
rect 12784 5729 12796 5763
rect 12768 5723 12796 5729
rect 12768 5720 12774 5723
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11532 5664 11713 5692
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 12894 5652 12900 5704
rect 12952 5652 12958 5704
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 14826 5692 14832 5704
rect 13771 5664 14832 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 1655 5625 1716 5631
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 1688 5556 1716 5625
rect 5810 5556 5816 5568
rect 1688 5528 5816 5556
rect 5810 5516 5816 5528
rect 5868 5556 5874 5568
rect 8294 5556 8300 5568
rect 5868 5528 8300 5556
rect 5868 5516 5874 5528
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 9324 5556 9352 5652
rect 11790 5624 11796 5636
rect 11532 5596 11796 5624
rect 11532 5556 11560 5596
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 14274 5584 14280 5636
rect 14332 5584 14338 5636
rect 9324 5528 11560 5556
rect 11609 5559 11667 5565
rect 11609 5525 11621 5559
rect 11655 5556 11667 5559
rect 11698 5556 11704 5568
rect 11655 5528 11704 5556
rect 11655 5525 11667 5528
rect 11609 5519 11667 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 1104 5466 14971 5488
rect 1104 5414 4376 5466
rect 4428 5414 4440 5466
rect 4492 5414 4504 5466
rect 4556 5414 4568 5466
rect 4620 5414 4632 5466
rect 4684 5414 7803 5466
rect 7855 5414 7867 5466
rect 7919 5414 7931 5466
rect 7983 5414 7995 5466
rect 8047 5414 8059 5466
rect 8111 5414 11230 5466
rect 11282 5414 11294 5466
rect 11346 5414 11358 5466
rect 11410 5414 11422 5466
rect 11474 5414 11486 5466
rect 11538 5414 14657 5466
rect 14709 5414 14721 5466
rect 14773 5414 14785 5466
rect 14837 5414 14849 5466
rect 14901 5414 14913 5466
rect 14965 5414 14971 5466
rect 1104 5392 14971 5414
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 9033 5355 9091 5361
rect 7708 5324 8984 5352
rect 7708 5312 7714 5324
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2225 5287 2283 5293
rect 2225 5284 2237 5287
rect 1719 5256 2237 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2225 5253 2237 5256
rect 2271 5253 2283 5287
rect 8294 5255 8300 5296
rect 2225 5247 2283 5253
rect 8279 5249 8300 5255
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 3970 5216 3976 5228
rect 2179 5188 3976 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7248 5188 8033 5216
rect 7248 5176 7254 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8279 5215 8291 5249
rect 8352 5244 8358 5296
rect 8956 5284 8984 5324
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 10134 5352 10140 5364
rect 9079 5324 10140 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 10244 5324 12173 5352
rect 10244 5284 10272 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 13265 5355 13323 5361
rect 13265 5321 13277 5355
rect 13311 5352 13323 5355
rect 13354 5352 13360 5364
rect 13311 5324 13360 5352
rect 13311 5321 13323 5324
rect 13265 5315 13323 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15102 5284 15108 5296
rect 8956 5256 10272 5284
rect 11992 5256 15108 5284
rect 8325 5218 8340 5244
rect 8325 5215 8337 5218
rect 8279 5209 8337 5215
rect 8021 5179 8079 5185
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 992 4984 1777 5012
rect 992 4972 998 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 8036 5012 8064 5179
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 11992 5225 12020 5256
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 11977 5219 12035 5225
rect 8996 5188 9674 5216
rect 8996 5176 9002 5188
rect 8294 5012 8300 5024
rect 8036 4984 8300 5012
rect 1765 4975 1823 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 9646 5012 9674 5188
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 12495 5219 12553 5225
rect 12495 5216 12507 5219
rect 11977 5179 12035 5185
rect 12084 5188 12507 5216
rect 10778 5108 10784 5160
rect 10836 5148 10842 5160
rect 12084 5148 12112 5188
rect 12495 5185 12507 5188
rect 12541 5185 12553 5219
rect 12495 5179 12553 5185
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 13722 5216 13728 5228
rect 13679 5188 13728 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 13722 5176 13728 5188
rect 13780 5176 13786 5228
rect 13909 5219 13967 5225
rect 13909 5185 13921 5219
rect 13955 5216 13967 5219
rect 13998 5216 14004 5228
rect 13955 5188 14004 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 13998 5176 14004 5188
rect 14056 5176 14062 5228
rect 12241 5151 12299 5157
rect 12241 5148 12253 5151
rect 10836 5120 12112 5148
rect 12176 5120 12253 5148
rect 10836 5108 10842 5120
rect 12066 5040 12072 5092
rect 12124 5080 12130 5092
rect 12176 5080 12204 5120
rect 12241 5117 12253 5120
rect 12287 5117 12299 5151
rect 12241 5111 12299 5117
rect 12124 5052 12204 5080
rect 12124 5040 12130 5052
rect 12526 5012 12532 5024
rect 9646 4984 12532 5012
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 1104 4922 14812 4944
rect 1104 4870 2663 4922
rect 2715 4870 2727 4922
rect 2779 4870 2791 4922
rect 2843 4870 2855 4922
rect 2907 4870 2919 4922
rect 2971 4870 6090 4922
rect 6142 4870 6154 4922
rect 6206 4870 6218 4922
rect 6270 4870 6282 4922
rect 6334 4870 6346 4922
rect 6398 4870 9517 4922
rect 9569 4870 9581 4922
rect 9633 4870 9645 4922
rect 9697 4870 9709 4922
rect 9761 4870 9773 4922
rect 9825 4870 12944 4922
rect 12996 4870 13008 4922
rect 13060 4870 13072 4922
rect 13124 4870 13136 4922
rect 13188 4870 13200 4922
rect 13252 4870 14812 4922
rect 1104 4848 14812 4870
rect 842 4768 848 4820
rect 900 4808 906 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 900 4780 1593 4808
rect 900 4768 906 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 10873 4811 10931 4817
rect 1581 4771 1639 4777
rect 9876 4780 10548 4808
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 9876 4681 9904 4780
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 8352 4644 9873 4672
rect 8352 4632 8358 4644
rect 9861 4641 9873 4644
rect 9907 4641 9919 4675
rect 10520 4672 10548 4780
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 11974 4808 11980 4820
rect 10919 4780 11980 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12710 4808 12716 4820
rect 12299 4780 12716 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 13906 4768 13912 4820
rect 13964 4808 13970 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13964 4780 14381 4808
rect 13964 4768 13970 4780
rect 14369 4777 14381 4780
rect 14415 4777 14427 4811
rect 14369 4771 14427 4777
rect 11146 4672 11152 4684
rect 10520 4644 11152 4672
rect 9861 4635 9919 4641
rect 11146 4632 11152 4644
rect 11204 4672 11210 4684
rect 11241 4675 11299 4681
rect 11241 4672 11253 4675
rect 11204 4644 11253 4672
rect 11204 4632 11210 4644
rect 11241 4641 11253 4644
rect 11287 4641 11299 4675
rect 12084 4672 12112 4768
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12084 4644 12633 4672
rect 11241 4635 11299 4641
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12621 4635 12679 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 2038 4604 2044 4616
rect 1535 4576 2044 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 10103 4607 10161 4613
rect 10103 4604 10115 4607
rect 9968 4576 10115 4604
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 9968 4536 9996 4576
rect 10103 4573 10115 4576
rect 10149 4573 10161 4607
rect 10103 4567 10161 4573
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11483 4607 11541 4613
rect 11483 4604 11495 4607
rect 11112 4576 11495 4604
rect 11112 4564 11118 4576
rect 11483 4573 11495 4576
rect 11529 4573 11541 4607
rect 14277 4607 14335 4613
rect 12879 4577 12937 4583
rect 12879 4574 12891 4577
rect 11483 4567 11541 4573
rect 7340 4508 9996 4536
rect 7340 4496 7346 4508
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 12820 4546 12891 4574
rect 12820 4536 12848 4546
rect 12879 4543 12891 4546
rect 12925 4543 12937 4577
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 15194 4604 15200 4616
rect 14323 4576 15200 4604
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 12879 4537 12937 4543
rect 12676 4508 12848 4536
rect 12676 4496 12682 4508
rect 1104 4378 14971 4400
rect 1104 4326 4376 4378
rect 4428 4326 4440 4378
rect 4492 4326 4504 4378
rect 4556 4326 4568 4378
rect 4620 4326 4632 4378
rect 4684 4326 7803 4378
rect 7855 4326 7867 4378
rect 7919 4326 7931 4378
rect 7983 4326 7995 4378
rect 8047 4326 8059 4378
rect 8111 4326 11230 4378
rect 11282 4326 11294 4378
rect 11346 4326 11358 4378
rect 11410 4326 11422 4378
rect 11474 4326 11486 4378
rect 11538 4326 14657 4378
rect 14709 4326 14721 4378
rect 14773 4326 14785 4378
rect 14837 4326 14849 4378
rect 14901 4326 14913 4378
rect 14965 4326 14971 4378
rect 1104 4304 14971 4326
rect 12618 4224 12624 4276
rect 12676 4224 12682 4276
rect 10594 4156 10600 4208
rect 10652 4196 10658 4208
rect 12636 4196 12664 4224
rect 10652 4168 12572 4196
rect 12636 4168 13216 4196
rect 10652 4156 10658 4168
rect 750 4088 756 4140
rect 808 4128 814 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 808 4100 1409 4128
rect 808 4088 814 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 1397 4091 1455 4097
rect 8754 4088 8760 4100
rect 8812 4128 8818 4140
rect 11146 4128 11152 4140
rect 8812 4100 11152 4128
rect 8812 4088 8818 4100
rect 11146 4088 11152 4100
rect 11204 4088 11210 4140
rect 11882 4137 11888 4140
rect 11851 4131 11888 4137
rect 11851 4097 11863 4131
rect 11851 4091 11888 4097
rect 11882 4088 11888 4091
rect 11940 4088 11946 4140
rect 12544 4072 12572 4168
rect 13188 4158 13216 4168
rect 13247 4161 13305 4167
rect 13247 4158 13259 4161
rect 13188 4130 13259 4158
rect 13247 4127 13259 4130
rect 13293 4127 13305 4161
rect 13247 4121 13305 4127
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8352 4032 8493 4060
rect 8352 4020 8358 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9493 3995 9551 4001
rect 9493 3992 9505 3995
rect 9456 3964 9505 3992
rect 9456 3952 9462 3964
rect 9493 3961 9505 3964
rect 9539 3961 9551 3995
rect 9493 3955 9551 3961
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 3418 3924 3424 3936
rect 1627 3896 3424 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 11624 3924 11652 4023
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 12989 4063 13047 4069
rect 12989 4060 13001 4063
rect 12584 4032 13001 4060
rect 12584 4020 12590 4032
rect 12989 4029 13001 4032
rect 13035 4029 13047 4063
rect 12989 4023 13047 4029
rect 12066 3924 12072 3936
rect 11624 3896 12072 3924
rect 12066 3884 12072 3896
rect 12124 3884 12130 3936
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 12400 3896 12633 3924
rect 12400 3884 12406 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14001 3927 14059 3933
rect 14001 3924 14013 3927
rect 13872 3896 14013 3924
rect 13872 3884 13878 3896
rect 14001 3893 14013 3896
rect 14047 3893 14059 3927
rect 14001 3887 14059 3893
rect 1104 3834 14812 3856
rect 1104 3782 2663 3834
rect 2715 3782 2727 3834
rect 2779 3782 2791 3834
rect 2843 3782 2855 3834
rect 2907 3782 2919 3834
rect 2971 3782 6090 3834
rect 6142 3782 6154 3834
rect 6206 3782 6218 3834
rect 6270 3782 6282 3834
rect 6334 3782 6346 3834
rect 6398 3782 9517 3834
rect 9569 3782 9581 3834
rect 9633 3782 9645 3834
rect 9697 3782 9709 3834
rect 9761 3782 9773 3834
rect 9825 3782 12944 3834
rect 12996 3782 13008 3834
rect 13060 3782 13072 3834
rect 13124 3782 13136 3834
rect 13188 3782 13200 3834
rect 13252 3782 14812 3834
rect 1104 3760 14812 3782
rect 13081 3723 13139 3729
rect 13081 3689 13093 3723
rect 13127 3720 13139 3723
rect 13262 3720 13268 3732
rect 13127 3692 13268 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 14366 3680 14372 3732
rect 14424 3680 14430 3732
rect 12066 3544 12072 3596
rect 12124 3544 12130 3596
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12311 3519 12369 3525
rect 12311 3516 12323 3519
rect 11204 3488 12323 3516
rect 11204 3476 11210 3488
rect 12311 3485 12323 3488
rect 12357 3485 12369 3519
rect 12311 3479 12369 3485
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 1104 3290 14971 3312
rect 1104 3238 4376 3290
rect 4428 3238 4440 3290
rect 4492 3238 4504 3290
rect 4556 3238 4568 3290
rect 4620 3238 4632 3290
rect 4684 3238 7803 3290
rect 7855 3238 7867 3290
rect 7919 3238 7931 3290
rect 7983 3238 7995 3290
rect 8047 3238 8059 3290
rect 8111 3238 11230 3290
rect 11282 3238 11294 3290
rect 11346 3238 11358 3290
rect 11410 3238 11422 3290
rect 11474 3238 11486 3290
rect 11538 3238 14657 3290
rect 14709 3238 14721 3290
rect 14773 3238 14785 3290
rect 14837 3238 14849 3290
rect 14901 3238 14913 3290
rect 14965 3238 14971 3290
rect 1104 3216 14971 3238
rect 1104 2746 14812 2768
rect 1104 2694 2663 2746
rect 2715 2694 2727 2746
rect 2779 2694 2791 2746
rect 2843 2694 2855 2746
rect 2907 2694 2919 2746
rect 2971 2694 6090 2746
rect 6142 2694 6154 2746
rect 6206 2694 6218 2746
rect 6270 2694 6282 2746
rect 6334 2694 6346 2746
rect 6398 2694 9517 2746
rect 9569 2694 9581 2746
rect 9633 2694 9645 2746
rect 9697 2694 9709 2746
rect 9761 2694 9773 2746
rect 9825 2694 12944 2746
rect 12996 2694 13008 2746
rect 13060 2694 13072 2746
rect 13124 2694 13136 2746
rect 13188 2694 13200 2746
rect 13252 2694 14812 2746
rect 1104 2672 14812 2694
rect 1210 2592 1216 2644
rect 1268 2632 1274 2644
rect 4433 2635 4491 2641
rect 4433 2632 4445 2635
rect 1268 2604 4445 2632
rect 1268 2592 1274 2604
rect 4433 2601 4445 2604
rect 4479 2601 4491 2635
rect 4433 2595 4491 2601
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 4341 2363 4399 2369
rect 4341 2360 4353 2363
rect 4120 2332 4353 2360
rect 4120 2320 4126 2332
rect 4341 2329 4353 2332
rect 4387 2329 4399 2363
rect 4341 2323 4399 2329
rect 1104 2202 14971 2224
rect 1104 2150 4376 2202
rect 4428 2150 4440 2202
rect 4492 2150 4504 2202
rect 4556 2150 4568 2202
rect 4620 2150 4632 2202
rect 4684 2150 7803 2202
rect 7855 2150 7867 2202
rect 7919 2150 7931 2202
rect 7983 2150 7995 2202
rect 8047 2150 8059 2202
rect 8111 2150 11230 2202
rect 11282 2150 11294 2202
rect 11346 2150 11358 2202
rect 11410 2150 11422 2202
rect 11474 2150 11486 2202
rect 11538 2150 14657 2202
rect 14709 2150 14721 2202
rect 14773 2150 14785 2202
rect 14837 2150 14849 2202
rect 14901 2150 14913 2202
rect 14965 2150 14971 2202
rect 1104 2128 14971 2150
rect 4062 2048 4068 2100
rect 4120 2048 4126 2100
rect 5077 2091 5135 2097
rect 5077 2057 5089 2091
rect 5123 2057 5135 2091
rect 5077 2051 5135 2057
rect 2222 1980 2228 2032
rect 2280 2020 2286 2032
rect 5092 2020 5120 2051
rect 5810 2048 5816 2100
rect 5868 2048 5874 2100
rect 6549 2091 6607 2097
rect 6549 2057 6561 2091
rect 6595 2088 6607 2091
rect 6638 2088 6644 2100
rect 6595 2060 6644 2088
rect 6595 2057 6607 2060
rect 6549 2051 6607 2057
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 7190 2048 7196 2100
rect 7248 2048 7254 2100
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 7929 2091 7987 2097
rect 7929 2088 7941 2091
rect 7708 2060 7941 2088
rect 7708 2048 7714 2060
rect 7929 2057 7941 2060
rect 7975 2057 7987 2091
rect 7929 2051 7987 2057
rect 8662 2048 8668 2100
rect 8720 2048 8726 2100
rect 10870 2048 10876 2100
rect 10928 2048 10934 2100
rect 12345 2091 12403 2097
rect 12345 2057 12357 2091
rect 12391 2088 12403 2091
rect 12434 2088 12440 2100
rect 12391 2060 12440 2088
rect 12391 2057 12403 2060
rect 12345 2051 12403 2057
rect 12434 2048 12440 2060
rect 12492 2048 12498 2100
rect 13081 2091 13139 2097
rect 13081 2057 13093 2091
rect 13127 2088 13139 2091
rect 13354 2088 13360 2100
rect 13127 2060 13360 2088
rect 13127 2057 13139 2060
rect 13081 2051 13139 2057
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 14185 2091 14243 2097
rect 14185 2057 14197 2091
rect 14231 2088 14243 2091
rect 15746 2088 15752 2100
rect 14231 2060 15752 2088
rect 14231 2057 14243 2060
rect 14185 2051 14243 2057
rect 15746 2048 15752 2060
rect 15804 2048 15810 2100
rect 12066 2020 12072 2032
rect 2280 1992 5120 2020
rect 6886 1992 12072 2020
rect 2280 1980 2286 1992
rect 2130 1912 2136 1964
rect 2188 1912 2194 1964
rect 4246 1912 4252 1964
rect 4304 1912 4310 1964
rect 4982 1912 4988 1964
rect 5040 1912 5046 1964
rect 5718 1912 5724 1964
rect 5776 1912 5782 1964
rect 6454 1912 6460 1964
rect 6512 1912 6518 1964
rect 2961 1887 3019 1893
rect 2961 1853 2973 1887
rect 3007 1884 3019 1887
rect 6886 1884 6914 1992
rect 12066 1980 12072 1992
rect 12124 1980 12130 2032
rect 13446 1980 13452 2032
rect 13504 2020 13510 2032
rect 14093 2023 14151 2029
rect 14093 2020 14105 2023
rect 13504 1992 14105 2020
rect 13504 1980 13510 1992
rect 14093 1989 14105 1992
rect 14139 1989 14151 2023
rect 14093 1983 14151 1989
rect 15010 1980 15016 2032
rect 15068 1980 15074 2032
rect 7098 1912 7104 1964
rect 7156 1912 7162 1964
rect 7834 1912 7840 1964
rect 7892 1912 7898 1964
rect 8570 1912 8576 1964
rect 8628 1912 8634 1964
rect 9306 1912 9312 1964
rect 9364 1912 9370 1964
rect 10042 1912 10048 1964
rect 10100 1912 10106 1964
rect 10778 1912 10784 1964
rect 10836 1912 10842 1964
rect 11606 1912 11612 1964
rect 11664 1912 11670 1964
rect 12250 1912 12256 1964
rect 12308 1912 12314 1964
rect 12989 1955 13047 1961
rect 12989 1921 13001 1955
rect 13035 1952 13047 1955
rect 13262 1952 13268 1964
rect 13035 1924 13268 1952
rect 13035 1921 13047 1924
rect 12989 1915 13047 1921
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 13722 1912 13728 1964
rect 13780 1912 13786 1964
rect 13909 1955 13967 1961
rect 13909 1921 13921 1955
rect 13955 1952 13967 1955
rect 15028 1952 15056 1980
rect 13955 1924 15056 1952
rect 13955 1921 13967 1924
rect 13909 1915 13967 1921
rect 3007 1856 6914 1884
rect 7760 1856 10272 1884
rect 3007 1853 3019 1856
rect 2961 1847 3019 1853
rect 3234 1776 3240 1828
rect 3292 1816 3298 1828
rect 7760 1816 7788 1856
rect 10244 1825 10272 1856
rect 10229 1819 10287 1825
rect 3292 1788 7788 1816
rect 7852 1788 9444 1816
rect 3292 1776 3298 1788
rect 2406 1708 2412 1760
rect 2464 1748 2470 1760
rect 7852 1748 7880 1788
rect 9416 1757 9444 1788
rect 10229 1785 10241 1819
rect 10275 1785 10287 1819
rect 10229 1779 10287 1785
rect 2464 1720 7880 1748
rect 9401 1751 9459 1757
rect 2464 1708 2470 1720
rect 9401 1717 9413 1751
rect 9447 1717 9459 1751
rect 9401 1711 9459 1717
rect 11698 1708 11704 1760
rect 11756 1708 11762 1760
rect 1104 1658 14812 1680
rect 1104 1606 2663 1658
rect 2715 1606 2727 1658
rect 2779 1606 2791 1658
rect 2843 1606 2855 1658
rect 2907 1606 2919 1658
rect 2971 1606 6090 1658
rect 6142 1606 6154 1658
rect 6206 1606 6218 1658
rect 6270 1606 6282 1658
rect 6334 1606 6346 1658
rect 6398 1606 9517 1658
rect 9569 1606 9581 1658
rect 9633 1606 9645 1658
rect 9697 1606 9709 1658
rect 9761 1606 9773 1658
rect 9825 1606 12944 1658
rect 12996 1606 13008 1658
rect 13060 1606 13072 1658
rect 13124 1606 13136 1658
rect 13188 1606 13200 1658
rect 13252 1606 14812 1658
rect 1104 1584 14812 1606
rect 4246 1504 4252 1556
rect 4304 1544 4310 1556
rect 4341 1547 4399 1553
rect 4341 1544 4353 1547
rect 4304 1516 4353 1544
rect 4304 1504 4310 1516
rect 4341 1513 4353 1516
rect 4387 1513 4399 1547
rect 4341 1507 4399 1513
rect 4982 1504 4988 1556
rect 5040 1544 5046 1556
rect 5077 1547 5135 1553
rect 5077 1544 5089 1547
rect 5040 1516 5089 1544
rect 5040 1504 5046 1516
rect 5077 1513 5089 1516
rect 5123 1513 5135 1547
rect 5077 1507 5135 1513
rect 5718 1504 5724 1556
rect 5776 1544 5782 1556
rect 5813 1547 5871 1553
rect 5813 1544 5825 1547
rect 5776 1516 5825 1544
rect 5776 1504 5782 1516
rect 5813 1513 5825 1516
rect 5859 1513 5871 1547
rect 5813 1507 5871 1513
rect 6454 1504 6460 1556
rect 6512 1544 6518 1556
rect 6549 1547 6607 1553
rect 6549 1544 6561 1547
rect 6512 1516 6561 1544
rect 6512 1504 6518 1516
rect 6549 1513 6561 1516
rect 6595 1513 6607 1547
rect 6549 1507 6607 1513
rect 7098 1504 7104 1556
rect 7156 1544 7162 1556
rect 7285 1547 7343 1553
rect 7285 1544 7297 1547
rect 7156 1516 7297 1544
rect 7156 1504 7162 1516
rect 7285 1513 7297 1516
rect 7331 1513 7343 1547
rect 7285 1507 7343 1513
rect 7834 1504 7840 1556
rect 7892 1544 7898 1556
rect 8021 1547 8079 1553
rect 8021 1544 8033 1547
rect 7892 1516 8033 1544
rect 7892 1504 7898 1516
rect 8021 1513 8033 1516
rect 8067 1513 8079 1547
rect 8021 1507 8079 1513
rect 8570 1504 8576 1556
rect 8628 1544 8634 1556
rect 8941 1547 8999 1553
rect 8941 1544 8953 1547
rect 8628 1516 8953 1544
rect 8628 1504 8634 1516
rect 8941 1513 8953 1516
rect 8987 1513 8999 1547
rect 8941 1507 8999 1513
rect 9306 1504 9312 1556
rect 9364 1544 9370 1556
rect 9493 1547 9551 1553
rect 9493 1544 9505 1547
rect 9364 1516 9505 1544
rect 9364 1504 9370 1516
rect 9493 1513 9505 1516
rect 9539 1513 9551 1547
rect 9493 1507 9551 1513
rect 10042 1504 10048 1556
rect 10100 1544 10106 1556
rect 10229 1547 10287 1553
rect 10229 1544 10241 1547
rect 10100 1516 10241 1544
rect 10100 1504 10106 1516
rect 10229 1513 10241 1516
rect 10275 1513 10287 1547
rect 10229 1507 10287 1513
rect 10778 1504 10784 1556
rect 10836 1544 10842 1556
rect 10965 1547 11023 1553
rect 10965 1544 10977 1547
rect 10836 1516 10977 1544
rect 10836 1504 10842 1516
rect 10965 1513 10977 1516
rect 11011 1513 11023 1547
rect 10965 1507 11023 1513
rect 11606 1504 11612 1556
rect 11664 1544 11670 1556
rect 11701 1547 11759 1553
rect 11701 1544 11713 1547
rect 11664 1516 11713 1544
rect 11664 1504 11670 1516
rect 11701 1513 11713 1516
rect 11747 1513 11759 1547
rect 11701 1507 11759 1513
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 12437 1547 12495 1553
rect 12437 1544 12449 1547
rect 12308 1516 12449 1544
rect 12308 1504 12314 1516
rect 12437 1513 12449 1516
rect 12483 1513 12495 1547
rect 12437 1507 12495 1513
rect 13173 1547 13231 1553
rect 13173 1513 13185 1547
rect 13219 1544 13231 1547
rect 13262 1544 13268 1556
rect 13219 1516 13268 1544
rect 13219 1513 13231 1516
rect 13173 1507 13231 1513
rect 13262 1504 13268 1516
rect 13320 1504 13326 1556
rect 13446 1504 13452 1556
rect 13504 1504 13510 1556
rect 13722 1504 13728 1556
rect 13780 1504 13786 1556
rect 13832 1380 14044 1408
rect 1302 1300 1308 1352
rect 1360 1340 1366 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1360 1312 1409 1340
rect 1360 1300 1366 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 1578 1300 1584 1352
rect 1636 1340 1642 1352
rect 2685 1343 2743 1349
rect 1636 1312 2360 1340
rect 1636 1300 1642 1312
rect 2222 1232 2228 1284
rect 2280 1232 2286 1284
rect 2332 1272 2360 1312
rect 2685 1309 2697 1343
rect 2731 1340 2743 1343
rect 2774 1340 2780 1352
rect 2731 1312 2780 1340
rect 2731 1309 2743 1312
rect 2685 1303 2743 1309
rect 2774 1300 2780 1312
rect 2832 1300 2838 1352
rect 2884 1312 3556 1340
rect 2884 1272 2912 1312
rect 2332 1244 2912 1272
rect 3421 1275 3479 1281
rect 3421 1241 3433 1275
rect 3467 1241 3479 1275
rect 3528 1272 3556 1312
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4246 1300 4252 1352
rect 4304 1340 4310 1352
rect 4525 1343 4583 1349
rect 4525 1340 4537 1343
rect 4304 1312 4537 1340
rect 4304 1300 4310 1312
rect 4525 1309 4537 1312
rect 4571 1309 4583 1343
rect 4525 1303 4583 1309
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 5261 1343 5319 1349
rect 5261 1340 5273 1343
rect 5040 1312 5273 1340
rect 5040 1300 5046 1312
rect 5261 1309 5273 1312
rect 5307 1309 5319 1343
rect 5261 1303 5319 1309
rect 5718 1300 5724 1352
rect 5776 1340 5782 1352
rect 5997 1343 6055 1349
rect 5997 1340 6009 1343
rect 5776 1312 6009 1340
rect 5776 1300 5782 1312
rect 5997 1309 6009 1312
rect 6043 1309 6055 1343
rect 5997 1303 6055 1309
rect 6454 1300 6460 1352
rect 6512 1340 6518 1352
rect 6733 1343 6791 1349
rect 6733 1340 6745 1343
rect 6512 1312 6745 1340
rect 6512 1300 6518 1312
rect 6733 1309 6745 1312
rect 6779 1309 6791 1343
rect 6733 1303 6791 1309
rect 7466 1300 7472 1352
rect 7524 1300 7530 1352
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 8720 1312 9137 1340
rect 8720 1300 8726 1312
rect 9125 1309 9137 1312
rect 9171 1309 9183 1343
rect 9125 1303 9183 1309
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 10410 1300 10416 1352
rect 10468 1300 10474 1352
rect 10870 1300 10876 1352
rect 10928 1340 10934 1352
rect 11149 1343 11207 1349
rect 11149 1340 11161 1343
rect 10928 1312 11161 1340
rect 10928 1300 10934 1312
rect 11149 1309 11161 1312
rect 11195 1309 11207 1343
rect 11149 1303 11207 1309
rect 11606 1300 11612 1352
rect 11664 1340 11670 1352
rect 11885 1343 11943 1349
rect 11885 1340 11897 1343
rect 11664 1312 11897 1340
rect 11664 1300 11670 1312
rect 11885 1309 11897 1312
rect 11931 1309 11943 1343
rect 11885 1303 11943 1309
rect 12342 1300 12348 1352
rect 12400 1340 12406 1352
rect 12621 1343 12679 1349
rect 12621 1340 12633 1343
rect 12400 1312 12633 1340
rect 12400 1300 12406 1312
rect 12621 1309 12633 1312
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 13078 1300 13084 1352
rect 13136 1300 13142 1352
rect 13354 1300 13360 1352
rect 13412 1300 13418 1352
rect 13633 1343 13691 1349
rect 13633 1309 13645 1343
rect 13679 1340 13691 1343
rect 13832 1340 13860 1380
rect 13679 1312 13860 1340
rect 13679 1309 13691 1312
rect 13633 1303 13691 1309
rect 13906 1300 13912 1352
rect 13964 1300 13970 1352
rect 14016 1340 14044 1380
rect 14550 1340 14556 1352
rect 14016 1312 14556 1340
rect 14550 1300 14556 1312
rect 14608 1300 14614 1352
rect 15470 1300 15476 1352
rect 15528 1300 15534 1352
rect 4065 1275 4123 1281
rect 4065 1272 4077 1275
rect 3528 1244 4077 1272
rect 3421 1235 3479 1241
rect 4065 1241 4077 1244
rect 4111 1241 4123 1275
rect 12526 1272 12532 1284
rect 4065 1235 4123 1241
rect 5000 1244 12532 1272
rect 3436 1204 3464 1235
rect 5000 1204 5028 1244
rect 12526 1232 12532 1244
rect 12584 1232 12590 1284
rect 14185 1275 14243 1281
rect 14185 1272 14197 1275
rect 12912 1244 14197 1272
rect 12912 1213 12940 1244
rect 14185 1241 14197 1244
rect 14231 1241 14243 1275
rect 14185 1235 14243 1241
rect 14369 1275 14427 1281
rect 14369 1241 14381 1275
rect 14415 1272 14427 1275
rect 15488 1272 15516 1300
rect 14415 1244 15516 1272
rect 14415 1241 14427 1244
rect 14369 1235 14427 1241
rect 3436 1176 5028 1204
rect 12897 1207 12955 1213
rect 12897 1173 12909 1207
rect 12943 1173 12955 1207
rect 12897 1167 12955 1173
rect 1104 1114 14971 1136
rect 1104 1062 4376 1114
rect 4428 1062 4440 1114
rect 4492 1062 4504 1114
rect 4556 1062 4568 1114
rect 4620 1062 4632 1114
rect 4684 1062 7803 1114
rect 7855 1062 7867 1114
rect 7919 1062 7931 1114
rect 7983 1062 7995 1114
rect 8047 1062 8059 1114
rect 8111 1062 11230 1114
rect 11282 1062 11294 1114
rect 11346 1062 11358 1114
rect 11410 1062 11422 1114
rect 11474 1062 11486 1114
rect 11538 1062 14657 1114
rect 14709 1062 14721 1114
rect 14773 1062 14785 1114
rect 14837 1062 14849 1114
rect 14901 1062 14913 1114
rect 14965 1062 14971 1114
rect 1104 1040 14971 1062
rect 2222 960 2228 1012
rect 2280 1000 2286 1012
rect 8386 1000 8392 1012
rect 2280 972 8392 1000
rect 2280 960 2286 972
rect 8386 960 8392 972
rect 8444 960 8450 1012
rect 13078 960 13084 1012
rect 13136 1000 13142 1012
rect 15286 1000 15292 1012
rect 13136 972 15292 1000
rect 13136 960 13142 972
rect 15286 960 15292 972
rect 15344 960 15350 1012
<< via1 >>
rect 4376 43494 4428 43546
rect 4440 43494 4492 43546
rect 4504 43494 4556 43546
rect 4568 43494 4620 43546
rect 4632 43494 4684 43546
rect 7803 43494 7855 43546
rect 7867 43494 7919 43546
rect 7931 43494 7983 43546
rect 7995 43494 8047 43546
rect 8059 43494 8111 43546
rect 11230 43494 11282 43546
rect 11294 43494 11346 43546
rect 11358 43494 11410 43546
rect 11422 43494 11474 43546
rect 11486 43494 11538 43546
rect 14657 43494 14709 43546
rect 14721 43494 14773 43546
rect 14785 43494 14837 43546
rect 14849 43494 14901 43546
rect 14913 43494 14965 43546
rect 572 43392 624 43444
rect 2780 43392 2832 43444
rect 3516 43392 3568 43444
rect 4252 43392 4304 43444
rect 4988 43392 5040 43444
rect 5724 43392 5776 43444
rect 6460 43392 6512 43444
rect 7196 43392 7248 43444
rect 8208 43435 8260 43444
rect 8208 43401 8217 43435
rect 8217 43401 8251 43435
rect 8251 43401 8260 43435
rect 8208 43392 8260 43401
rect 8668 43392 8720 43444
rect 9404 43392 9456 43444
rect 10140 43392 10192 43444
rect 10876 43392 10928 43444
rect 12348 43392 12400 43444
rect 13084 43392 13136 43444
rect 13820 43392 13872 43444
rect 1768 43256 1820 43308
rect 2136 43299 2188 43308
rect 2136 43265 2145 43299
rect 2145 43265 2179 43299
rect 2179 43265 2188 43299
rect 2136 43256 2188 43265
rect 2504 43299 2556 43308
rect 2504 43265 2513 43299
rect 2513 43265 2547 43299
rect 2547 43265 2556 43299
rect 2504 43256 2556 43265
rect 3056 43256 3108 43308
rect 3792 43299 3844 43308
rect 3792 43265 3801 43299
rect 3801 43265 3835 43299
rect 3835 43265 3844 43299
rect 3792 43256 3844 43265
rect 4344 43299 4396 43308
rect 4344 43265 4353 43299
rect 4353 43265 4387 43299
rect 4387 43265 4396 43299
rect 4344 43256 4396 43265
rect 5080 43299 5132 43308
rect 5080 43265 5089 43299
rect 5089 43265 5123 43299
rect 5123 43265 5132 43299
rect 5080 43256 5132 43265
rect 5816 43299 5868 43308
rect 5816 43265 5825 43299
rect 5825 43265 5859 43299
rect 5859 43265 5868 43299
rect 5816 43256 5868 43265
rect 6552 43299 6604 43308
rect 6552 43265 6561 43299
rect 6561 43265 6595 43299
rect 6595 43265 6604 43299
rect 6552 43256 6604 43265
rect 7288 43299 7340 43308
rect 7288 43265 7297 43299
rect 7297 43265 7331 43299
rect 7331 43265 7340 43299
rect 7288 43256 7340 43265
rect 8024 43299 8076 43308
rect 8024 43265 8033 43299
rect 8033 43265 8067 43299
rect 8067 43265 8076 43299
rect 8024 43256 8076 43265
rect 8944 43299 8996 43308
rect 8944 43265 8953 43299
rect 8953 43265 8987 43299
rect 8987 43265 8996 43299
rect 8944 43256 8996 43265
rect 9312 43256 9364 43308
rect 10232 43299 10284 43308
rect 10232 43265 10241 43299
rect 10241 43265 10275 43299
rect 10275 43265 10284 43299
rect 10232 43256 10284 43265
rect 11612 43299 11664 43308
rect 11612 43265 11621 43299
rect 11621 43265 11655 43299
rect 11655 43265 11664 43299
rect 11612 43256 11664 43265
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 12532 43299 12584 43308
rect 12532 43265 12541 43299
rect 12541 43265 12575 43299
rect 12575 43265 12584 43299
rect 12532 43256 12584 43265
rect 13268 43256 13320 43308
rect 13636 43299 13688 43308
rect 13636 43265 13645 43299
rect 13645 43265 13679 43299
rect 13679 43265 13688 43299
rect 13636 43256 13688 43265
rect 14096 43299 14148 43308
rect 14096 43265 14105 43299
rect 14105 43265 14139 43299
rect 14139 43265 14148 43299
rect 14096 43256 14148 43265
rect 14556 43188 14608 43240
rect 2044 43120 2096 43172
rect 1400 43052 1452 43104
rect 11704 43052 11756 43104
rect 2663 42950 2715 43002
rect 2727 42950 2779 43002
rect 2791 42950 2843 43002
rect 2855 42950 2907 43002
rect 2919 42950 2971 43002
rect 6090 42950 6142 43002
rect 6154 42950 6206 43002
rect 6218 42950 6270 43002
rect 6282 42950 6334 43002
rect 6346 42950 6398 43002
rect 9517 42950 9569 43002
rect 9581 42950 9633 43002
rect 9645 42950 9697 43002
rect 9709 42950 9761 43002
rect 9773 42950 9825 43002
rect 12944 42950 12996 43002
rect 13008 42950 13060 43002
rect 13072 42950 13124 43002
rect 13136 42950 13188 43002
rect 13200 42950 13252 43002
rect 2136 42848 2188 42900
rect 3056 42848 3108 42900
rect 3792 42848 3844 42900
rect 4344 42848 4396 42900
rect 5816 42848 5868 42900
rect 6552 42848 6604 42900
rect 7288 42848 7340 42900
rect 8024 42848 8076 42900
rect 8944 42848 8996 42900
rect 9312 42891 9364 42900
rect 9312 42857 9321 42891
rect 9321 42857 9355 42891
rect 9355 42857 9364 42891
rect 9312 42848 9364 42857
rect 10232 42848 10284 42900
rect 11612 42848 11664 42900
rect 12072 42848 12124 42900
rect 12532 42848 12584 42900
rect 13268 42848 13320 42900
rect 13636 42848 13688 42900
rect 14096 42848 14148 42900
rect 15292 42712 15344 42764
rect 2228 42687 2280 42696
rect 2228 42653 2237 42687
rect 2237 42653 2271 42687
rect 2271 42653 2280 42687
rect 2228 42644 2280 42653
rect 2964 42687 3016 42696
rect 2964 42653 2973 42687
rect 2973 42653 3007 42687
rect 3007 42653 3016 42687
rect 2964 42644 3016 42653
rect 3516 42687 3568 42696
rect 3516 42653 3525 42687
rect 3525 42653 3559 42687
rect 3559 42653 3568 42687
rect 3516 42644 3568 42653
rect 1216 42576 1268 42628
rect 5908 42687 5960 42696
rect 5908 42653 5917 42687
rect 5917 42653 5951 42687
rect 5951 42653 5960 42687
rect 5908 42644 5960 42653
rect 6644 42687 6696 42696
rect 6644 42653 6653 42687
rect 6653 42653 6687 42687
rect 6687 42653 6696 42687
rect 6644 42644 6696 42653
rect 7288 42687 7340 42696
rect 7288 42653 7297 42687
rect 7297 42653 7331 42687
rect 7331 42653 7340 42687
rect 7288 42644 7340 42653
rect 8208 42644 8260 42696
rect 8760 42687 8812 42696
rect 8760 42653 8769 42687
rect 8769 42653 8803 42687
rect 8803 42653 8812 42687
rect 8760 42644 8812 42653
rect 9496 42687 9548 42696
rect 9496 42653 9505 42687
rect 9505 42653 9539 42687
rect 9539 42653 9548 42687
rect 9496 42644 9548 42653
rect 10232 42687 10284 42696
rect 10232 42653 10241 42687
rect 10241 42653 10275 42687
rect 10275 42653 10284 42687
rect 10232 42644 10284 42653
rect 10968 42687 11020 42696
rect 10968 42653 10977 42687
rect 10977 42653 11011 42687
rect 11011 42653 11020 42687
rect 10968 42644 11020 42653
rect 11704 42687 11756 42696
rect 11704 42653 11713 42687
rect 11713 42653 11747 42687
rect 11747 42653 11756 42687
rect 11704 42644 11756 42653
rect 12440 42687 12492 42696
rect 12440 42653 12449 42687
rect 12449 42653 12483 42687
rect 12483 42653 12492 42687
rect 12440 42644 12492 42653
rect 13176 42687 13228 42696
rect 13176 42653 13185 42687
rect 13185 42653 13219 42687
rect 13219 42653 13228 42687
rect 13176 42644 13228 42653
rect 14096 42644 14148 42696
rect 13544 42619 13596 42628
rect 13544 42585 13553 42619
rect 13553 42585 13587 42619
rect 13587 42585 13596 42619
rect 13544 42576 13596 42585
rect 14280 42508 14332 42560
rect 4376 42406 4428 42458
rect 4440 42406 4492 42458
rect 4504 42406 4556 42458
rect 4568 42406 4620 42458
rect 4632 42406 4684 42458
rect 7803 42406 7855 42458
rect 7867 42406 7919 42458
rect 7931 42406 7983 42458
rect 7995 42406 8047 42458
rect 8059 42406 8111 42458
rect 11230 42406 11282 42458
rect 11294 42406 11346 42458
rect 11358 42406 11410 42458
rect 11422 42406 11474 42458
rect 11486 42406 11538 42458
rect 14657 42406 14709 42458
rect 14721 42406 14773 42458
rect 14785 42406 14837 42458
rect 14849 42406 14901 42458
rect 14913 42406 14965 42458
rect 2228 42304 2280 42356
rect 2964 42304 3016 42356
rect 5908 42304 5960 42356
rect 6644 42304 6696 42356
rect 7288 42304 7340 42356
rect 8208 42304 8260 42356
rect 8760 42304 8812 42356
rect 9496 42304 9548 42356
rect 10232 42304 10284 42356
rect 10968 42304 11020 42356
rect 11704 42304 11756 42356
rect 12440 42304 12492 42356
rect 13176 42304 13228 42356
rect 13544 42304 13596 42356
rect 14280 42347 14332 42356
rect 14280 42313 14289 42347
rect 14289 42313 14323 42347
rect 14323 42313 14332 42347
rect 14280 42304 14332 42313
rect 2412 42236 2464 42288
rect 2228 42211 2280 42220
rect 2228 42177 2237 42211
rect 2237 42177 2271 42211
rect 2271 42177 2280 42211
rect 2228 42168 2280 42177
rect 3056 42211 3108 42220
rect 3056 42177 3065 42211
rect 3065 42177 3099 42211
rect 3099 42177 3108 42211
rect 3056 42168 3108 42177
rect 5724 42211 5776 42220
rect 5724 42177 5733 42211
rect 5733 42177 5767 42211
rect 5767 42177 5776 42211
rect 5724 42168 5776 42177
rect 6552 42211 6604 42220
rect 6552 42177 6561 42211
rect 6561 42177 6595 42211
rect 6595 42177 6604 42211
rect 6552 42168 6604 42177
rect 7288 42211 7340 42220
rect 7288 42177 7297 42211
rect 7297 42177 7331 42211
rect 7331 42177 7340 42211
rect 7288 42168 7340 42177
rect 8116 42211 8168 42220
rect 8116 42177 8125 42211
rect 8125 42177 8159 42211
rect 8159 42177 8168 42211
rect 8116 42168 8168 42177
rect 14096 42236 14148 42288
rect 3608 42100 3660 42152
rect 3240 42032 3292 42084
rect 10968 42211 11020 42220
rect 10968 42177 10977 42211
rect 10977 42177 11011 42211
rect 11011 42177 11020 42211
rect 10968 42168 11020 42177
rect 11704 42211 11756 42220
rect 11704 42177 11713 42211
rect 11713 42177 11747 42211
rect 11747 42177 11756 42211
rect 11704 42168 11756 42177
rect 12440 42211 12492 42220
rect 12440 42177 12449 42211
rect 12449 42177 12483 42211
rect 12483 42177 12492 42211
rect 12440 42168 12492 42177
rect 14004 42168 14056 42220
rect 14188 42211 14240 42220
rect 14188 42177 14197 42211
rect 14197 42177 14231 42211
rect 14231 42177 14240 42211
rect 14188 42168 14240 42177
rect 15752 42168 15804 42220
rect 15108 41964 15160 42016
rect 2663 41862 2715 41914
rect 2727 41862 2779 41914
rect 2791 41862 2843 41914
rect 2855 41862 2907 41914
rect 2919 41862 2971 41914
rect 6090 41862 6142 41914
rect 6154 41862 6206 41914
rect 6218 41862 6270 41914
rect 6282 41862 6334 41914
rect 6346 41862 6398 41914
rect 9517 41862 9569 41914
rect 9581 41862 9633 41914
rect 9645 41862 9697 41914
rect 9709 41862 9761 41914
rect 9773 41862 9825 41914
rect 12944 41862 12996 41914
rect 13008 41862 13060 41914
rect 13072 41862 13124 41914
rect 13136 41862 13188 41914
rect 13200 41862 13252 41914
rect 3056 41760 3108 41812
rect 14188 41760 14240 41812
rect 14004 41624 14056 41676
rect 15016 41624 15068 41676
rect 6920 41556 6972 41608
rect 15476 41556 15528 41608
rect 4376 41318 4428 41370
rect 4440 41318 4492 41370
rect 4504 41318 4556 41370
rect 4568 41318 4620 41370
rect 4632 41318 4684 41370
rect 7803 41318 7855 41370
rect 7867 41318 7919 41370
rect 7931 41318 7983 41370
rect 7995 41318 8047 41370
rect 8059 41318 8111 41370
rect 11230 41318 11282 41370
rect 11294 41318 11346 41370
rect 11358 41318 11410 41370
rect 11422 41318 11474 41370
rect 11486 41318 11538 41370
rect 14657 41318 14709 41370
rect 14721 41318 14773 41370
rect 14785 41318 14837 41370
rect 14849 41318 14901 41370
rect 14913 41318 14965 41370
rect 756 41080 808 41132
rect 8208 40876 8260 40928
rect 2663 40774 2715 40826
rect 2727 40774 2779 40826
rect 2791 40774 2843 40826
rect 2855 40774 2907 40826
rect 2919 40774 2971 40826
rect 6090 40774 6142 40826
rect 6154 40774 6206 40826
rect 6218 40774 6270 40826
rect 6282 40774 6334 40826
rect 6346 40774 6398 40826
rect 9517 40774 9569 40826
rect 9581 40774 9633 40826
rect 9645 40774 9697 40826
rect 9709 40774 9761 40826
rect 9773 40774 9825 40826
rect 12944 40774 12996 40826
rect 13008 40774 13060 40826
rect 13072 40774 13124 40826
rect 13136 40774 13188 40826
rect 13200 40774 13252 40826
rect 4376 40230 4428 40282
rect 4440 40230 4492 40282
rect 4504 40230 4556 40282
rect 4568 40230 4620 40282
rect 4632 40230 4684 40282
rect 7803 40230 7855 40282
rect 7867 40230 7919 40282
rect 7931 40230 7983 40282
rect 7995 40230 8047 40282
rect 8059 40230 8111 40282
rect 11230 40230 11282 40282
rect 11294 40230 11346 40282
rect 11358 40230 11410 40282
rect 11422 40230 11474 40282
rect 11486 40230 11538 40282
rect 14657 40230 14709 40282
rect 14721 40230 14773 40282
rect 14785 40230 14837 40282
rect 14849 40230 14901 40282
rect 14913 40230 14965 40282
rect 1400 40035 1452 40044
rect 1400 40001 1409 40035
rect 1409 40001 1443 40035
rect 1443 40001 1452 40035
rect 1400 39992 1452 40001
rect 13360 40035 13412 40044
rect 13360 40001 13369 40035
rect 13369 40001 13403 40035
rect 13403 40001 13412 40035
rect 13360 39992 13412 40001
rect 10968 39924 11020 39976
rect 7380 39788 7432 39840
rect 14004 39788 14056 39840
rect 14188 39831 14240 39840
rect 14188 39797 14197 39831
rect 14197 39797 14231 39831
rect 14231 39797 14240 39831
rect 14188 39788 14240 39797
rect 2663 39686 2715 39738
rect 2727 39686 2779 39738
rect 2791 39686 2843 39738
rect 2855 39686 2907 39738
rect 2919 39686 2971 39738
rect 6090 39686 6142 39738
rect 6154 39686 6206 39738
rect 6218 39686 6270 39738
rect 6282 39686 6334 39738
rect 6346 39686 6398 39738
rect 9517 39686 9569 39738
rect 9581 39686 9633 39738
rect 9645 39686 9697 39738
rect 9709 39686 9761 39738
rect 9773 39686 9825 39738
rect 12944 39686 12996 39738
rect 13008 39686 13060 39738
rect 13072 39686 13124 39738
rect 13136 39686 13188 39738
rect 13200 39686 13252 39738
rect 756 39380 808 39432
rect 8392 39380 8444 39432
rect 10968 39584 11020 39636
rect 13360 39584 13412 39636
rect 7380 39312 7432 39364
rect 12716 39423 12768 39432
rect 12716 39389 12725 39423
rect 12725 39389 12759 39423
rect 12759 39389 12768 39423
rect 12716 39380 12768 39389
rect 13360 39380 13412 39432
rect 7564 39244 7616 39296
rect 13912 39355 13964 39364
rect 13912 39321 13921 39355
rect 13921 39321 13955 39355
rect 13955 39321 13964 39355
rect 13912 39312 13964 39321
rect 14372 39287 14424 39296
rect 14372 39253 14381 39287
rect 14381 39253 14415 39287
rect 14415 39253 14424 39287
rect 14372 39244 14424 39253
rect 4376 39142 4428 39194
rect 4440 39142 4492 39194
rect 4504 39142 4556 39194
rect 4568 39142 4620 39194
rect 4632 39142 4684 39194
rect 7803 39142 7855 39194
rect 7867 39142 7919 39194
rect 7931 39142 7983 39194
rect 7995 39142 8047 39194
rect 8059 39142 8111 39194
rect 11230 39142 11282 39194
rect 11294 39142 11346 39194
rect 11358 39142 11410 39194
rect 11422 39142 11474 39194
rect 11486 39142 11538 39194
rect 14657 39142 14709 39194
rect 14721 39142 14773 39194
rect 14785 39142 14837 39194
rect 14849 39142 14901 39194
rect 14913 39142 14965 39194
rect 5080 39040 5132 39092
rect 12716 39040 12768 39092
rect 7564 38972 7616 39024
rect 5172 38947 5224 38956
rect 5172 38913 5181 38947
rect 5181 38913 5215 38947
rect 5215 38913 5224 38947
rect 5172 38904 5224 38913
rect 12624 38904 12676 38956
rect 12808 38904 12860 38956
rect 13452 38904 13504 38956
rect 13268 38700 13320 38752
rect 13636 38743 13688 38752
rect 13636 38709 13645 38743
rect 13645 38709 13679 38743
rect 13679 38709 13688 38743
rect 13636 38700 13688 38709
rect 14188 38743 14240 38752
rect 14188 38709 14197 38743
rect 14197 38709 14231 38743
rect 14231 38709 14240 38743
rect 14188 38700 14240 38709
rect 14464 38700 14516 38752
rect 2663 38598 2715 38650
rect 2727 38598 2779 38650
rect 2791 38598 2843 38650
rect 2855 38598 2907 38650
rect 2919 38598 2971 38650
rect 6090 38598 6142 38650
rect 6154 38598 6206 38650
rect 6218 38598 6270 38650
rect 6282 38598 6334 38650
rect 6346 38598 6398 38650
rect 9517 38598 9569 38650
rect 9581 38598 9633 38650
rect 9645 38598 9697 38650
rect 9709 38598 9761 38650
rect 9773 38598 9825 38650
rect 12944 38598 12996 38650
rect 13008 38598 13060 38650
rect 13072 38598 13124 38650
rect 13136 38598 13188 38650
rect 13200 38598 13252 38650
rect 5172 38496 5224 38548
rect 13360 38496 13412 38548
rect 12440 38428 12492 38480
rect 12716 38428 12768 38480
rect 756 38292 808 38344
rect 2136 38292 2188 38344
rect 11612 38292 11664 38344
rect 9404 38224 9456 38276
rect 13176 38335 13228 38344
rect 13176 38301 13185 38335
rect 13185 38301 13219 38335
rect 13219 38301 13228 38335
rect 13176 38292 13228 38301
rect 13268 38292 13320 38344
rect 13360 38292 13412 38344
rect 12624 38156 12676 38208
rect 13268 38156 13320 38208
rect 13820 38199 13872 38208
rect 13820 38165 13829 38199
rect 13829 38165 13863 38199
rect 13863 38165 13872 38199
rect 13820 38156 13872 38165
rect 14372 38199 14424 38208
rect 14372 38165 14381 38199
rect 14381 38165 14415 38199
rect 14415 38165 14424 38199
rect 14372 38156 14424 38165
rect 4376 38054 4428 38106
rect 4440 38054 4492 38106
rect 4504 38054 4556 38106
rect 4568 38054 4620 38106
rect 4632 38054 4684 38106
rect 7803 38054 7855 38106
rect 7867 38054 7919 38106
rect 7931 38054 7983 38106
rect 7995 38054 8047 38106
rect 8059 38054 8111 38106
rect 11230 38054 11282 38106
rect 11294 38054 11346 38106
rect 11358 38054 11410 38106
rect 11422 38054 11474 38106
rect 11486 38054 11538 38106
rect 14657 38054 14709 38106
rect 14721 38054 14773 38106
rect 14785 38054 14837 38106
rect 14849 38054 14901 38106
rect 14913 38054 14965 38106
rect 11796 37952 11848 38004
rect 12532 37952 12584 38004
rect 12440 37884 12492 37936
rect 13176 37952 13228 38004
rect 756 37816 808 37868
rect 10784 37816 10836 37868
rect 12072 37859 12124 37868
rect 12072 37825 12081 37859
rect 12081 37825 12115 37859
rect 12115 37825 12124 37859
rect 12072 37816 12124 37825
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 13084 37859 13136 37868
rect 13084 37825 13093 37859
rect 13093 37825 13127 37859
rect 13127 37825 13136 37859
rect 13084 37816 13136 37825
rect 13268 37816 13320 37868
rect 12348 37680 12400 37732
rect 5724 37612 5776 37664
rect 6552 37612 6604 37664
rect 12624 37612 12676 37664
rect 13544 37612 13596 37664
rect 13636 37655 13688 37664
rect 13636 37621 13645 37655
rect 13645 37621 13679 37655
rect 13679 37621 13688 37655
rect 13636 37612 13688 37621
rect 14188 37655 14240 37664
rect 14188 37621 14197 37655
rect 14197 37621 14231 37655
rect 14231 37621 14240 37655
rect 14188 37612 14240 37621
rect 2663 37510 2715 37562
rect 2727 37510 2779 37562
rect 2791 37510 2843 37562
rect 2855 37510 2907 37562
rect 2919 37510 2971 37562
rect 6090 37510 6142 37562
rect 6154 37510 6206 37562
rect 6218 37510 6270 37562
rect 6282 37510 6334 37562
rect 6346 37510 6398 37562
rect 9517 37510 9569 37562
rect 9581 37510 9633 37562
rect 9645 37510 9697 37562
rect 9709 37510 9761 37562
rect 9773 37510 9825 37562
rect 12944 37510 12996 37562
rect 13008 37510 13060 37562
rect 13072 37510 13124 37562
rect 13136 37510 13188 37562
rect 13200 37510 13252 37562
rect 10784 37451 10836 37460
rect 10784 37417 10793 37451
rect 10793 37417 10827 37451
rect 10827 37417 10836 37451
rect 10784 37408 10836 37417
rect 12072 37408 12124 37460
rect 12348 37451 12400 37460
rect 12348 37417 12357 37451
rect 12357 37417 12391 37451
rect 12391 37417 12400 37451
rect 12348 37408 12400 37417
rect 12624 37272 12676 37324
rect 10968 37247 11020 37256
rect 10968 37213 10977 37247
rect 10977 37213 11011 37247
rect 11011 37213 11020 37247
rect 10968 37204 11020 37213
rect 6552 37136 6604 37188
rect 11888 37204 11940 37256
rect 12808 37247 12860 37256
rect 12808 37213 12817 37247
rect 12817 37213 12851 37247
rect 12851 37213 12860 37247
rect 12808 37204 12860 37213
rect 12900 37204 12952 37256
rect 13268 37204 13320 37256
rect 12164 37136 12216 37188
rect 13544 37179 13596 37188
rect 13544 37145 13553 37179
rect 13553 37145 13587 37179
rect 13587 37145 13596 37179
rect 13544 37136 13596 37145
rect 12716 37068 12768 37120
rect 13176 37111 13228 37120
rect 13176 37077 13185 37111
rect 13185 37077 13219 37111
rect 13219 37077 13228 37111
rect 13176 37068 13228 37077
rect 13636 37111 13688 37120
rect 13636 37077 13645 37111
rect 13645 37077 13679 37111
rect 13679 37077 13688 37111
rect 13636 37068 13688 37077
rect 14372 37111 14424 37120
rect 14372 37077 14381 37111
rect 14381 37077 14415 37111
rect 14415 37077 14424 37111
rect 14372 37068 14424 37077
rect 4376 36966 4428 37018
rect 4440 36966 4492 37018
rect 4504 36966 4556 37018
rect 4568 36966 4620 37018
rect 4632 36966 4684 37018
rect 7803 36966 7855 37018
rect 7867 36966 7919 37018
rect 7931 36966 7983 37018
rect 7995 36966 8047 37018
rect 8059 36966 8111 37018
rect 11230 36966 11282 37018
rect 11294 36966 11346 37018
rect 11358 36966 11410 37018
rect 11422 36966 11474 37018
rect 11486 36966 11538 37018
rect 14657 36966 14709 37018
rect 14721 36966 14773 37018
rect 14785 36966 14837 37018
rect 14849 36966 14901 37018
rect 14913 36966 14965 37018
rect 2228 36864 2280 36916
rect 10968 36864 11020 36916
rect 11612 36907 11664 36916
rect 11612 36873 11621 36907
rect 11621 36873 11655 36907
rect 11655 36873 11664 36907
rect 11612 36864 11664 36873
rect 11888 36907 11940 36916
rect 11888 36873 11897 36907
rect 11897 36873 11931 36907
rect 11931 36873 11940 36907
rect 11888 36864 11940 36873
rect 12348 36864 12400 36916
rect 13176 36864 13228 36916
rect 756 36728 808 36780
rect 4252 36728 4304 36780
rect 5172 36660 5224 36712
rect 8300 36592 8352 36644
rect 11336 36592 11388 36644
rect 11888 36660 11940 36712
rect 12716 36771 12768 36780
rect 12716 36737 12725 36771
rect 12725 36737 12759 36771
rect 12759 36737 12768 36771
rect 12716 36728 12768 36737
rect 12992 36771 13044 36780
rect 12992 36737 13001 36771
rect 13001 36737 13035 36771
rect 13035 36737 13044 36771
rect 12992 36728 13044 36737
rect 13452 36728 13504 36780
rect 13360 36592 13412 36644
rect 13452 36592 13504 36644
rect 13636 36660 13688 36712
rect 12532 36567 12584 36576
rect 12532 36533 12541 36567
rect 12541 36533 12575 36567
rect 12575 36533 12584 36567
rect 12532 36524 12584 36533
rect 13820 36567 13872 36576
rect 13820 36533 13829 36567
rect 13829 36533 13863 36567
rect 13863 36533 13872 36567
rect 13820 36524 13872 36533
rect 15292 36524 15344 36576
rect 2663 36422 2715 36474
rect 2727 36422 2779 36474
rect 2791 36422 2843 36474
rect 2855 36422 2907 36474
rect 2919 36422 2971 36474
rect 6090 36422 6142 36474
rect 6154 36422 6206 36474
rect 6218 36422 6270 36474
rect 6282 36422 6334 36474
rect 6346 36422 6398 36474
rect 9517 36422 9569 36474
rect 9581 36422 9633 36474
rect 9645 36422 9697 36474
rect 9709 36422 9761 36474
rect 9773 36422 9825 36474
rect 12944 36422 12996 36474
rect 13008 36422 13060 36474
rect 13072 36422 13124 36474
rect 13136 36422 13188 36474
rect 13200 36422 13252 36474
rect 7288 36320 7340 36372
rect 12164 36363 12216 36372
rect 12164 36329 12173 36363
rect 12173 36329 12207 36363
rect 12207 36329 12216 36363
rect 12164 36320 12216 36329
rect 12532 36320 12584 36372
rect 12716 36320 12768 36372
rect 13452 36320 13504 36372
rect 12624 36252 12676 36304
rect 12900 36252 12952 36304
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 12440 36116 12492 36168
rect 12624 36159 12676 36168
rect 12624 36125 12633 36159
rect 12633 36125 12667 36159
rect 12667 36125 12676 36159
rect 12624 36116 12676 36125
rect 12716 36116 12768 36168
rect 12808 36116 12860 36168
rect 13176 36116 13228 36168
rect 13452 36116 13504 36168
rect 10968 36048 11020 36100
rect 13360 35980 13412 36032
rect 13728 35980 13780 36032
rect 15108 35980 15160 36032
rect 4376 35878 4428 35930
rect 4440 35878 4492 35930
rect 4504 35878 4556 35930
rect 4568 35878 4620 35930
rect 4632 35878 4684 35930
rect 7803 35878 7855 35930
rect 7867 35878 7919 35930
rect 7931 35878 7983 35930
rect 7995 35878 8047 35930
rect 8059 35878 8111 35930
rect 11230 35878 11282 35930
rect 11294 35878 11346 35930
rect 11358 35878 11410 35930
rect 11422 35878 11474 35930
rect 11486 35878 11538 35930
rect 14657 35878 14709 35930
rect 14721 35878 14773 35930
rect 14785 35878 14837 35930
rect 14849 35878 14901 35930
rect 14913 35878 14965 35930
rect 10416 35683 10468 35692
rect 10416 35649 10425 35683
rect 10425 35649 10459 35683
rect 10459 35649 10468 35683
rect 10416 35640 10468 35649
rect 10692 35683 10744 35692
rect 10692 35649 10701 35683
rect 10701 35649 10735 35683
rect 10735 35649 10744 35683
rect 10692 35640 10744 35649
rect 11980 35708 12032 35760
rect 13452 35708 13504 35760
rect 11888 35640 11940 35692
rect 11520 35615 11572 35624
rect 11520 35581 11529 35615
rect 11529 35581 11563 35615
rect 11563 35581 11572 35615
rect 11520 35572 11572 35581
rect 12440 35572 12492 35624
rect 13176 35572 13228 35624
rect 10968 35504 11020 35556
rect 14004 35640 14056 35692
rect 11152 35436 11204 35488
rect 12532 35479 12584 35488
rect 12532 35445 12541 35479
rect 12541 35445 12575 35479
rect 12575 35445 12584 35479
rect 12532 35436 12584 35445
rect 15108 35504 15160 35556
rect 13820 35479 13872 35488
rect 13820 35445 13829 35479
rect 13829 35445 13863 35479
rect 13863 35445 13872 35479
rect 13820 35436 13872 35445
rect 14372 35479 14424 35488
rect 14372 35445 14381 35479
rect 14381 35445 14415 35479
rect 14415 35445 14424 35479
rect 14372 35436 14424 35445
rect 2663 35334 2715 35386
rect 2727 35334 2779 35386
rect 2791 35334 2843 35386
rect 2855 35334 2907 35386
rect 2919 35334 2971 35386
rect 6090 35334 6142 35386
rect 6154 35334 6206 35386
rect 6218 35334 6270 35386
rect 6282 35334 6334 35386
rect 6346 35334 6398 35386
rect 9517 35334 9569 35386
rect 9581 35334 9633 35386
rect 9645 35334 9697 35386
rect 9709 35334 9761 35386
rect 9773 35334 9825 35386
rect 12944 35334 12996 35386
rect 13008 35334 13060 35386
rect 13072 35334 13124 35386
rect 13136 35334 13188 35386
rect 13200 35334 13252 35386
rect 1768 35275 1820 35284
rect 1768 35241 1777 35275
rect 1777 35241 1811 35275
rect 1811 35241 1820 35275
rect 1768 35232 1820 35241
rect 10416 35232 10468 35284
rect 10692 35232 10744 35284
rect 13636 35232 13688 35284
rect 5908 35096 5960 35148
rect 11796 35096 11848 35148
rect 756 35028 808 35080
rect 1952 35071 2004 35080
rect 1952 35037 1961 35071
rect 1961 35037 1995 35071
rect 1995 35037 2004 35071
rect 1952 35028 2004 35037
rect 9680 35071 9732 35080
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 9680 35028 9732 35037
rect 9036 34960 9088 35012
rect 11060 35028 11112 35080
rect 12348 35096 12400 35148
rect 12072 34960 12124 35012
rect 12624 35028 12676 35080
rect 13728 35028 13780 35080
rect 13544 35003 13596 35012
rect 13544 34969 13553 35003
rect 13553 34969 13587 35003
rect 13587 34969 13596 35003
rect 13544 34960 13596 34969
rect 13912 35003 13964 35012
rect 13912 34969 13921 35003
rect 13921 34969 13955 35003
rect 13955 34969 13964 35003
rect 13912 34960 13964 34969
rect 11704 34935 11756 34944
rect 11704 34901 11713 34935
rect 11713 34901 11747 34935
rect 11747 34901 11756 34935
rect 11704 34892 11756 34901
rect 12900 34935 12952 34944
rect 12900 34901 12909 34935
rect 12909 34901 12943 34935
rect 12943 34901 12952 34935
rect 12900 34892 12952 34901
rect 13176 34935 13228 34944
rect 13176 34901 13185 34935
rect 13185 34901 13219 34935
rect 13219 34901 13228 34935
rect 13176 34892 13228 34901
rect 14096 34935 14148 34944
rect 14096 34901 14105 34935
rect 14105 34901 14139 34935
rect 14139 34901 14148 34935
rect 14096 34892 14148 34901
rect 4376 34790 4428 34842
rect 4440 34790 4492 34842
rect 4504 34790 4556 34842
rect 4568 34790 4620 34842
rect 4632 34790 4684 34842
rect 7803 34790 7855 34842
rect 7867 34790 7919 34842
rect 7931 34790 7983 34842
rect 7995 34790 8047 34842
rect 8059 34790 8111 34842
rect 11230 34790 11282 34842
rect 11294 34790 11346 34842
rect 11358 34790 11410 34842
rect 11422 34790 11474 34842
rect 11486 34790 11538 34842
rect 14657 34790 14709 34842
rect 14721 34790 14773 34842
rect 14785 34790 14837 34842
rect 14849 34790 14901 34842
rect 14913 34790 14965 34842
rect 1952 34688 2004 34740
rect 9680 34688 9732 34740
rect 4804 34620 4856 34672
rect 5448 34620 5500 34672
rect 9036 34620 9088 34672
rect 10968 34731 11020 34740
rect 10968 34697 10977 34731
rect 10977 34697 11011 34731
rect 11011 34697 11020 34731
rect 10968 34688 11020 34697
rect 11152 34688 11204 34740
rect 12072 34688 12124 34740
rect 12900 34688 12952 34740
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 1952 34595 2004 34604
rect 1952 34561 1961 34595
rect 1961 34561 1995 34595
rect 1995 34561 2004 34595
rect 1952 34552 2004 34561
rect 5816 34552 5868 34604
rect 6460 34484 6512 34536
rect 8300 34484 8352 34536
rect 9220 34595 9272 34604
rect 9220 34561 9229 34595
rect 9229 34561 9263 34595
rect 9263 34561 9272 34595
rect 9220 34552 9272 34561
rect 9312 34552 9364 34604
rect 9956 34595 10008 34604
rect 9956 34561 9965 34595
rect 9965 34561 9999 34595
rect 9999 34561 10008 34595
rect 9956 34552 10008 34561
rect 11888 34620 11940 34672
rect 10784 34552 10836 34604
rect 11796 34595 11848 34604
rect 11796 34561 11805 34595
rect 11805 34561 11839 34595
rect 11839 34561 11848 34595
rect 11796 34552 11848 34561
rect 12256 34595 12308 34604
rect 12256 34561 12265 34595
rect 12265 34561 12299 34595
rect 12299 34561 12308 34595
rect 12256 34552 12308 34561
rect 13176 34688 13228 34740
rect 10140 34416 10192 34468
rect 11980 34416 12032 34468
rect 12440 34416 12492 34468
rect 12716 34484 12768 34536
rect 13452 34552 13504 34604
rect 12808 34416 12860 34468
rect 13268 34348 13320 34400
rect 13636 34391 13688 34400
rect 13636 34357 13645 34391
rect 13645 34357 13679 34391
rect 13679 34357 13688 34391
rect 13636 34348 13688 34357
rect 14188 34391 14240 34400
rect 14188 34357 14197 34391
rect 14197 34357 14231 34391
rect 14231 34357 14240 34391
rect 14188 34348 14240 34357
rect 2663 34246 2715 34298
rect 2727 34246 2779 34298
rect 2791 34246 2843 34298
rect 2855 34246 2907 34298
rect 2919 34246 2971 34298
rect 6090 34246 6142 34298
rect 6154 34246 6206 34298
rect 6218 34246 6270 34298
rect 6282 34246 6334 34298
rect 6346 34246 6398 34298
rect 9517 34246 9569 34298
rect 9581 34246 9633 34298
rect 9645 34246 9697 34298
rect 9709 34246 9761 34298
rect 9773 34246 9825 34298
rect 12944 34246 12996 34298
rect 13008 34246 13060 34298
rect 13072 34246 13124 34298
rect 13136 34246 13188 34298
rect 13200 34246 13252 34298
rect 1952 34144 2004 34196
rect 9312 34144 9364 34196
rect 9956 34144 10008 34196
rect 10784 34144 10836 34196
rect 11704 34144 11756 34196
rect 13728 34076 13780 34128
rect 7104 33940 7156 33992
rect 9128 33983 9180 33992
rect 9128 33949 9137 33983
rect 9137 33949 9171 33983
rect 9171 33949 9180 33983
rect 9128 33940 9180 33949
rect 9404 33983 9456 33992
rect 9404 33949 9413 33983
rect 9413 33949 9447 33983
rect 9447 33949 9456 33983
rect 9404 33940 9456 33949
rect 9588 33940 9640 33992
rect 13820 34008 13872 34060
rect 9864 33872 9916 33924
rect 11612 33983 11664 33992
rect 11612 33949 11621 33983
rect 11621 33949 11655 33983
rect 11655 33949 11664 33983
rect 11612 33940 11664 33949
rect 12256 33940 12308 33992
rect 13176 33983 13228 33992
rect 13176 33949 13185 33983
rect 13185 33949 13219 33983
rect 13219 33949 13228 33983
rect 13176 33940 13228 33949
rect 13360 33940 13412 33992
rect 11704 33804 11756 33856
rect 12716 33804 12768 33856
rect 13912 33915 13964 33924
rect 13912 33881 13921 33915
rect 13921 33881 13955 33915
rect 13955 33881 13964 33915
rect 13912 33872 13964 33881
rect 14004 33872 14056 33924
rect 14372 33847 14424 33856
rect 14372 33813 14381 33847
rect 14381 33813 14415 33847
rect 14415 33813 14424 33847
rect 14372 33804 14424 33813
rect 4376 33702 4428 33754
rect 4440 33702 4492 33754
rect 4504 33702 4556 33754
rect 4568 33702 4620 33754
rect 4632 33702 4684 33754
rect 7803 33702 7855 33754
rect 7867 33702 7919 33754
rect 7931 33702 7983 33754
rect 7995 33702 8047 33754
rect 8059 33702 8111 33754
rect 11230 33702 11282 33754
rect 11294 33702 11346 33754
rect 11358 33702 11410 33754
rect 11422 33702 11474 33754
rect 11486 33702 11538 33754
rect 14657 33702 14709 33754
rect 14721 33702 14773 33754
rect 14785 33702 14837 33754
rect 14849 33702 14901 33754
rect 14913 33702 14965 33754
rect 3700 33600 3752 33652
rect 6460 33600 6512 33652
rect 9404 33600 9456 33652
rect 9588 33643 9640 33652
rect 9588 33609 9597 33643
rect 9597 33609 9631 33643
rect 9631 33609 9640 33643
rect 9588 33600 9640 33609
rect 9864 33643 9916 33652
rect 9864 33609 9873 33643
rect 9873 33609 9907 33643
rect 9907 33609 9916 33643
rect 9864 33600 9916 33609
rect 13268 33600 13320 33652
rect 756 33464 808 33516
rect 8300 33507 8352 33516
rect 8300 33473 8309 33507
rect 8309 33473 8343 33507
rect 8343 33473 8352 33507
rect 8300 33464 8352 33473
rect 6460 33396 6512 33448
rect 7012 33328 7064 33380
rect 10600 33507 10652 33516
rect 10600 33473 10609 33507
rect 10609 33473 10643 33507
rect 10643 33473 10652 33507
rect 10600 33464 10652 33473
rect 11888 33464 11940 33516
rect 12348 33464 12400 33516
rect 12716 33464 12768 33516
rect 13728 33532 13780 33584
rect 11520 33439 11572 33448
rect 11520 33405 11529 33439
rect 11529 33405 11563 33439
rect 11563 33405 11572 33439
rect 11520 33396 11572 33405
rect 13452 33396 13504 33448
rect 12808 33260 12860 33312
rect 14280 33328 14332 33380
rect 13636 33303 13688 33312
rect 13636 33269 13645 33303
rect 13645 33269 13679 33303
rect 13679 33269 13688 33303
rect 13636 33260 13688 33269
rect 14188 33303 14240 33312
rect 14188 33269 14197 33303
rect 14197 33269 14231 33303
rect 14231 33269 14240 33303
rect 14188 33260 14240 33269
rect 2663 33158 2715 33210
rect 2727 33158 2779 33210
rect 2791 33158 2843 33210
rect 2855 33158 2907 33210
rect 2919 33158 2971 33210
rect 6090 33158 6142 33210
rect 6154 33158 6206 33210
rect 6218 33158 6270 33210
rect 6282 33158 6334 33210
rect 6346 33158 6398 33210
rect 9517 33158 9569 33210
rect 9581 33158 9633 33210
rect 9645 33158 9697 33210
rect 9709 33158 9761 33210
rect 9773 33158 9825 33210
rect 12944 33158 12996 33210
rect 13008 33158 13060 33210
rect 13072 33158 13124 33210
rect 13136 33158 13188 33210
rect 13200 33158 13252 33210
rect 10600 33056 10652 33108
rect 11060 33056 11112 33108
rect 11428 33031 11480 33040
rect 11428 32997 11437 33031
rect 11437 32997 11471 33031
rect 11471 32997 11480 33031
rect 11428 32988 11480 32997
rect 13728 33056 13780 33108
rect 15568 32988 15620 33040
rect 756 32852 808 32904
rect 9956 32852 10008 32904
rect 1676 32716 1728 32768
rect 10968 32716 11020 32768
rect 11428 32852 11480 32904
rect 12072 32784 12124 32836
rect 12900 32852 12952 32904
rect 13360 32895 13412 32904
rect 13360 32861 13369 32895
rect 13369 32861 13403 32895
rect 13403 32861 13412 32895
rect 13360 32852 13412 32861
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 11796 32716 11848 32768
rect 12624 32716 12676 32768
rect 15108 32784 15160 32836
rect 14280 32759 14332 32768
rect 14280 32725 14289 32759
rect 14289 32725 14323 32759
rect 14323 32725 14332 32759
rect 14280 32716 14332 32725
rect 4376 32614 4428 32666
rect 4440 32614 4492 32666
rect 4504 32614 4556 32666
rect 4568 32614 4620 32666
rect 4632 32614 4684 32666
rect 7803 32614 7855 32666
rect 7867 32614 7919 32666
rect 7931 32614 7983 32666
rect 7995 32614 8047 32666
rect 8059 32614 8111 32666
rect 11230 32614 11282 32666
rect 11294 32614 11346 32666
rect 11358 32614 11410 32666
rect 11422 32614 11474 32666
rect 11486 32614 11538 32666
rect 14657 32614 14709 32666
rect 14721 32614 14773 32666
rect 14785 32614 14837 32666
rect 14849 32614 14901 32666
rect 14913 32614 14965 32666
rect 1676 32512 1728 32564
rect 11060 32512 11112 32564
rect 11336 32512 11388 32564
rect 13268 32512 13320 32564
rect 7104 32376 7156 32428
rect 7656 32376 7708 32428
rect 8392 32444 8444 32496
rect 9128 32444 9180 32496
rect 10048 32444 10100 32496
rect 10968 32444 11020 32496
rect 12440 32444 12492 32496
rect 11796 32419 11848 32428
rect 11796 32385 11803 32419
rect 11803 32385 11837 32419
rect 11837 32385 11848 32419
rect 11796 32376 11848 32385
rect 12164 32376 12216 32428
rect 13728 32419 13780 32428
rect 13728 32385 13737 32419
rect 13737 32385 13771 32419
rect 13771 32385 13780 32419
rect 13728 32376 13780 32385
rect 14188 32419 14240 32428
rect 14188 32385 14197 32419
rect 14197 32385 14231 32419
rect 14231 32385 14240 32419
rect 14188 32376 14240 32385
rect 12716 32308 12768 32360
rect 13636 32308 13688 32360
rect 9036 32215 9088 32224
rect 9036 32181 9045 32215
rect 9045 32181 9079 32215
rect 9079 32181 9088 32215
rect 9036 32172 9088 32181
rect 10416 32215 10468 32224
rect 10416 32181 10425 32215
rect 10425 32181 10459 32215
rect 10459 32181 10468 32215
rect 10416 32172 10468 32181
rect 11152 32215 11204 32224
rect 11152 32181 11161 32215
rect 11161 32181 11195 32215
rect 11195 32181 11204 32215
rect 11152 32172 11204 32181
rect 11612 32172 11664 32224
rect 12716 32172 12768 32224
rect 13912 32172 13964 32224
rect 14004 32215 14056 32224
rect 14004 32181 14013 32215
rect 14013 32181 14047 32215
rect 14047 32181 14056 32215
rect 14004 32172 14056 32181
rect 14372 32215 14424 32224
rect 14372 32181 14381 32215
rect 14381 32181 14415 32215
rect 14415 32181 14424 32215
rect 14372 32172 14424 32181
rect 2663 32070 2715 32122
rect 2727 32070 2779 32122
rect 2791 32070 2843 32122
rect 2855 32070 2907 32122
rect 2919 32070 2971 32122
rect 6090 32070 6142 32122
rect 6154 32070 6206 32122
rect 6218 32070 6270 32122
rect 6282 32070 6334 32122
rect 6346 32070 6398 32122
rect 9517 32070 9569 32122
rect 9581 32070 9633 32122
rect 9645 32070 9697 32122
rect 9709 32070 9761 32122
rect 9773 32070 9825 32122
rect 12944 32070 12996 32122
rect 13008 32070 13060 32122
rect 13072 32070 13124 32122
rect 13136 32070 13188 32122
rect 13200 32070 13252 32122
rect 1768 31968 1820 32020
rect 10140 31968 10192 32020
rect 11152 31968 11204 32020
rect 8208 31900 8260 31952
rect 11336 31943 11388 31952
rect 11336 31909 11345 31943
rect 11345 31909 11379 31943
rect 11379 31909 11388 31943
rect 11336 31900 11388 31909
rect 11704 31900 11756 31952
rect 6920 31875 6972 31884
rect 6920 31841 6929 31875
rect 6929 31841 6963 31875
rect 6963 31841 6972 31875
rect 6920 31832 6972 31841
rect 12164 32011 12216 32020
rect 12164 31977 12173 32011
rect 12173 31977 12207 32011
rect 12207 31977 12216 32011
rect 12164 31968 12216 31977
rect 12440 31968 12492 32020
rect 14188 31968 14240 32020
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 8116 31764 8168 31816
rect 9220 31764 9272 31816
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 12532 31832 12584 31884
rect 12624 31764 12676 31816
rect 12992 31807 13044 31816
rect 12992 31773 13001 31807
rect 13001 31773 13035 31807
rect 13035 31773 13044 31807
rect 12992 31764 13044 31773
rect 15660 31764 15712 31816
rect 7472 31696 7524 31748
rect 11520 31628 11572 31680
rect 11704 31628 11756 31680
rect 11796 31628 11848 31680
rect 12256 31628 12308 31680
rect 12440 31628 12492 31680
rect 13360 31628 13412 31680
rect 13912 31628 13964 31680
rect 14188 31671 14240 31680
rect 14188 31637 14197 31671
rect 14197 31637 14231 31671
rect 14231 31637 14240 31671
rect 14188 31628 14240 31637
rect 4376 31526 4428 31578
rect 4440 31526 4492 31578
rect 4504 31526 4556 31578
rect 4568 31526 4620 31578
rect 4632 31526 4684 31578
rect 7803 31526 7855 31578
rect 7867 31526 7919 31578
rect 7931 31526 7983 31578
rect 7995 31526 8047 31578
rect 8059 31526 8111 31578
rect 11230 31526 11282 31578
rect 11294 31526 11346 31578
rect 11358 31526 11410 31578
rect 11422 31526 11474 31578
rect 11486 31526 11538 31578
rect 14657 31526 14709 31578
rect 14721 31526 14773 31578
rect 14785 31526 14837 31578
rect 14849 31526 14901 31578
rect 14913 31526 14965 31578
rect 10968 31467 11020 31476
rect 10968 31433 10977 31467
rect 10977 31433 11011 31467
rect 11011 31433 11020 31467
rect 10968 31424 11020 31433
rect 11980 31424 12032 31476
rect 756 31288 808 31340
rect 5448 31288 5500 31340
rect 8300 31288 8352 31340
rect 9220 31356 9272 31408
rect 10508 31288 10560 31340
rect 11152 31331 11204 31340
rect 11152 31297 11161 31331
rect 11161 31297 11195 31331
rect 11195 31297 11204 31331
rect 11152 31288 11204 31297
rect 12164 31356 12216 31408
rect 14280 31356 14332 31408
rect 15384 31288 15436 31340
rect 1584 31127 1636 31136
rect 1584 31093 1593 31127
rect 1593 31093 1627 31127
rect 1627 31093 1636 31127
rect 1584 31084 1636 31093
rect 7564 31084 7616 31136
rect 11520 31263 11572 31272
rect 8300 31127 8352 31136
rect 8300 31093 8309 31127
rect 8309 31093 8343 31127
rect 8343 31093 8352 31127
rect 8300 31084 8352 31093
rect 11520 31229 11529 31263
rect 11529 31229 11563 31263
rect 11563 31229 11572 31263
rect 11520 31220 11572 31229
rect 12256 31220 12308 31272
rect 9864 31084 9916 31136
rect 11796 31084 11848 31136
rect 13268 31152 13320 31204
rect 12256 31084 12308 31136
rect 12624 31084 12676 31136
rect 13544 31084 13596 31136
rect 13636 31127 13688 31136
rect 13636 31093 13645 31127
rect 13645 31093 13679 31127
rect 13679 31093 13688 31127
rect 13636 31084 13688 31093
rect 15292 31084 15344 31136
rect 2663 30982 2715 31034
rect 2727 30982 2779 31034
rect 2791 30982 2843 31034
rect 2855 30982 2907 31034
rect 2919 30982 2971 31034
rect 6090 30982 6142 31034
rect 6154 30982 6206 31034
rect 6218 30982 6270 31034
rect 6282 30982 6334 31034
rect 6346 30982 6398 31034
rect 9517 30982 9569 31034
rect 9581 30982 9633 31034
rect 9645 30982 9697 31034
rect 9709 30982 9761 31034
rect 9773 30982 9825 31034
rect 12944 30982 12996 31034
rect 13008 30982 13060 31034
rect 13072 30982 13124 31034
rect 13136 30982 13188 31034
rect 13200 30982 13252 31034
rect 1584 30880 1636 30932
rect 5356 30880 5408 30932
rect 10324 30923 10376 30932
rect 10324 30889 10333 30923
rect 10333 30889 10367 30923
rect 10367 30889 10376 30923
rect 10324 30880 10376 30889
rect 11152 30880 11204 30932
rect 11520 30923 11572 30932
rect 11520 30889 11529 30923
rect 11529 30889 11563 30923
rect 11563 30889 11572 30923
rect 11520 30880 11572 30889
rect 11796 30923 11848 30932
rect 11796 30889 11805 30923
rect 11805 30889 11839 30923
rect 11839 30889 11848 30923
rect 11796 30880 11848 30889
rect 12072 30923 12124 30932
rect 12072 30889 12081 30923
rect 12081 30889 12115 30923
rect 12115 30889 12124 30923
rect 12072 30880 12124 30889
rect 9680 30719 9732 30728
rect 9680 30685 9689 30719
rect 9689 30685 9723 30719
rect 9723 30685 9732 30719
rect 9680 30676 9732 30685
rect 10876 30719 10928 30728
rect 10876 30685 10885 30719
rect 10885 30685 10919 30719
rect 10919 30685 10928 30719
rect 10876 30676 10928 30685
rect 12624 30880 12676 30932
rect 13452 30744 13504 30796
rect 12440 30719 12492 30728
rect 12440 30685 12449 30719
rect 12449 30685 12483 30719
rect 12483 30685 12492 30719
rect 12440 30676 12492 30685
rect 3792 30540 3844 30592
rect 9956 30540 10008 30592
rect 12900 30608 12952 30660
rect 12992 30651 13044 30660
rect 12992 30617 13001 30651
rect 13001 30617 13035 30651
rect 13035 30617 13044 30651
rect 12992 30608 13044 30617
rect 13360 30651 13412 30660
rect 13360 30617 13369 30651
rect 13369 30617 13403 30651
rect 13403 30617 13412 30651
rect 13360 30608 13412 30617
rect 12716 30540 12768 30592
rect 14556 30608 14608 30660
rect 15108 30540 15160 30592
rect 4376 30438 4428 30490
rect 4440 30438 4492 30490
rect 4504 30438 4556 30490
rect 4568 30438 4620 30490
rect 4632 30438 4684 30490
rect 7803 30438 7855 30490
rect 7867 30438 7919 30490
rect 7931 30438 7983 30490
rect 7995 30438 8047 30490
rect 8059 30438 8111 30490
rect 11230 30438 11282 30490
rect 11294 30438 11346 30490
rect 11358 30438 11410 30490
rect 11422 30438 11474 30490
rect 11486 30438 11538 30490
rect 14657 30438 14709 30490
rect 14721 30438 14773 30490
rect 14785 30438 14837 30490
rect 14849 30438 14901 30490
rect 14913 30438 14965 30490
rect 7104 30336 7156 30388
rect 9128 30336 9180 30388
rect 13728 30336 13780 30388
rect 756 30200 808 30252
rect 6828 30268 6880 30320
rect 7196 30268 7248 30320
rect 8484 30268 8536 30320
rect 7012 30200 7064 30252
rect 7380 30200 7432 30252
rect 9036 30132 9088 30184
rect 10416 30243 10468 30252
rect 10416 30209 10425 30243
rect 10425 30209 10459 30243
rect 10459 30209 10468 30243
rect 10416 30200 10468 30209
rect 12808 30243 12860 30252
rect 12808 30209 12817 30243
rect 12817 30209 12851 30243
rect 12851 30209 12860 30243
rect 12808 30200 12860 30209
rect 14004 30243 14056 30252
rect 14004 30209 14013 30243
rect 14013 30209 14047 30243
rect 14047 30209 14056 30243
rect 14004 30200 14056 30209
rect 9312 30132 9364 30184
rect 9772 30132 9824 30184
rect 9864 30175 9916 30184
rect 9864 30141 9873 30175
rect 9873 30141 9907 30175
rect 9907 30141 9916 30175
rect 9864 30132 9916 30141
rect 3884 30064 3936 30116
rect 2412 29996 2464 30048
rect 7380 30039 7432 30048
rect 7380 30005 7389 30039
rect 7389 30005 7423 30039
rect 7423 30005 7432 30039
rect 7380 29996 7432 30005
rect 9680 30064 9732 30116
rect 10324 30132 10376 30184
rect 11612 30175 11664 30184
rect 11612 30141 11621 30175
rect 11621 30141 11655 30175
rect 11655 30141 11664 30175
rect 11612 30132 11664 30141
rect 11796 30175 11848 30184
rect 11796 30141 11805 30175
rect 11805 30141 11839 30175
rect 11839 30141 11848 30175
rect 11796 30132 11848 30141
rect 11888 30064 11940 30116
rect 13360 30132 13412 30184
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 12072 29996 12124 30048
rect 13912 30064 13964 30116
rect 12624 29996 12676 30048
rect 14280 30039 14332 30048
rect 14280 30005 14289 30039
rect 14289 30005 14323 30039
rect 14323 30005 14332 30039
rect 14280 29996 14332 30005
rect 15752 29996 15804 30048
rect 2663 29894 2715 29946
rect 2727 29894 2779 29946
rect 2791 29894 2843 29946
rect 2855 29894 2907 29946
rect 2919 29894 2971 29946
rect 6090 29894 6142 29946
rect 6154 29894 6206 29946
rect 6218 29894 6270 29946
rect 6282 29894 6334 29946
rect 6346 29894 6398 29946
rect 9517 29894 9569 29946
rect 9581 29894 9633 29946
rect 9645 29894 9697 29946
rect 9709 29894 9761 29946
rect 9773 29894 9825 29946
rect 12944 29894 12996 29946
rect 13008 29894 13060 29946
rect 13072 29894 13124 29946
rect 13136 29894 13188 29946
rect 13200 29894 13252 29946
rect 2044 29792 2096 29844
rect 2412 29792 2464 29844
rect 7380 29792 7432 29844
rect 8300 29792 8352 29844
rect 8760 29767 8812 29776
rect 8760 29733 8769 29767
rect 8769 29733 8803 29767
rect 8803 29733 8812 29767
rect 8760 29724 8812 29733
rect 8944 29724 8996 29776
rect 4252 29656 4304 29708
rect 5540 29699 5592 29708
rect 5540 29665 5549 29699
rect 5549 29665 5583 29699
rect 5583 29665 5592 29699
rect 5540 29656 5592 29665
rect 7656 29656 7708 29708
rect 9220 29656 9272 29708
rect 10876 29792 10928 29844
rect 11060 29792 11112 29844
rect 12164 29792 12216 29844
rect 13452 29835 13504 29844
rect 13452 29801 13461 29835
rect 13461 29801 13495 29835
rect 13495 29801 13504 29835
rect 13452 29792 13504 29801
rect 12256 29767 12308 29776
rect 12256 29733 12265 29767
rect 12265 29733 12299 29767
rect 12299 29733 12308 29767
rect 12256 29724 12308 29733
rect 13820 29724 13872 29776
rect 756 29588 808 29640
rect 5816 29631 5868 29640
rect 3884 29520 3936 29572
rect 5816 29597 5823 29631
rect 5823 29597 5857 29631
rect 5857 29597 5868 29631
rect 5816 29588 5868 29597
rect 6828 29588 6880 29640
rect 6552 29495 6604 29504
rect 6552 29461 6561 29495
rect 6561 29461 6595 29495
rect 6595 29461 6604 29495
rect 6552 29452 6604 29461
rect 6736 29452 6788 29504
rect 7840 29631 7892 29640
rect 7840 29597 7849 29631
rect 7849 29597 7883 29631
rect 7883 29597 7892 29631
rect 7840 29588 7892 29597
rect 8116 29631 8168 29640
rect 8116 29597 8125 29631
rect 8125 29597 8159 29631
rect 8159 29597 8168 29631
rect 8116 29588 8168 29597
rect 8944 29631 8996 29640
rect 8944 29597 8953 29631
rect 8953 29597 8987 29631
rect 8987 29597 8996 29631
rect 8944 29588 8996 29597
rect 9864 29631 9916 29640
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10048 29588 10100 29640
rect 11060 29631 11112 29640
rect 11060 29597 11069 29631
rect 11069 29597 11103 29631
rect 11103 29597 11112 29631
rect 11060 29588 11112 29597
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 12164 29656 12216 29708
rect 12624 29631 12676 29640
rect 12624 29597 12658 29631
rect 12658 29597 12676 29631
rect 12624 29588 12676 29597
rect 11796 29520 11848 29572
rect 13820 29588 13872 29640
rect 14372 29520 14424 29572
rect 10048 29452 10100 29504
rect 10416 29452 10468 29504
rect 12440 29452 12492 29504
rect 13912 29452 13964 29504
rect 14096 29495 14148 29504
rect 14096 29461 14105 29495
rect 14105 29461 14139 29495
rect 14139 29461 14148 29495
rect 14096 29452 14148 29461
rect 4376 29350 4428 29402
rect 4440 29350 4492 29402
rect 4504 29350 4556 29402
rect 4568 29350 4620 29402
rect 4632 29350 4684 29402
rect 7803 29350 7855 29402
rect 7867 29350 7919 29402
rect 7931 29350 7983 29402
rect 7995 29350 8047 29402
rect 8059 29350 8111 29402
rect 11230 29350 11282 29402
rect 11294 29350 11346 29402
rect 11358 29350 11410 29402
rect 11422 29350 11474 29402
rect 11486 29350 11538 29402
rect 14657 29350 14709 29402
rect 14721 29350 14773 29402
rect 14785 29350 14837 29402
rect 14849 29350 14901 29402
rect 14913 29350 14965 29402
rect 6552 29248 6604 29300
rect 8300 29248 8352 29300
rect 6736 29044 6788 29096
rect 6828 29087 6880 29096
rect 6828 29053 6837 29087
rect 6837 29053 6871 29087
rect 6871 29053 6880 29087
rect 6828 29044 6880 29053
rect 7840 29155 7892 29164
rect 7840 29121 7874 29155
rect 7874 29121 7892 29155
rect 7840 29112 7892 29121
rect 8024 29155 8076 29164
rect 8024 29121 8033 29155
rect 8033 29121 8067 29155
rect 8067 29121 8076 29155
rect 8024 29112 8076 29121
rect 9864 29248 9916 29300
rect 12716 29291 12768 29300
rect 12716 29257 12725 29291
rect 12725 29257 12759 29291
rect 12759 29257 12768 29291
rect 12716 29248 12768 29257
rect 12808 29248 12860 29300
rect 9036 29155 9088 29164
rect 5264 28976 5316 29028
rect 9036 29121 9045 29155
rect 9045 29121 9088 29155
rect 9036 29112 9088 29121
rect 8760 29087 8812 29096
rect 8760 29053 8769 29087
rect 8769 29053 8803 29087
rect 8803 29053 8812 29087
rect 8760 29044 8812 29053
rect 8668 28976 8720 29028
rect 11796 29112 11848 29164
rect 14188 29180 14240 29232
rect 11888 29044 11940 29096
rect 12900 29155 12952 29164
rect 12900 29121 12909 29155
rect 12909 29121 12943 29155
rect 12943 29121 12952 29155
rect 12900 29112 12952 29121
rect 12992 29112 13044 29164
rect 14004 29112 14056 29164
rect 13268 29044 13320 29096
rect 11796 29019 11848 29028
rect 11796 28985 11805 29019
rect 11805 28985 11839 29019
rect 11839 28985 11848 29019
rect 11796 28976 11848 28985
rect 10140 28908 10192 28960
rect 10692 28908 10744 28960
rect 12256 28908 12308 28960
rect 13636 28951 13688 28960
rect 13636 28917 13645 28951
rect 13645 28917 13679 28951
rect 13679 28917 13688 28951
rect 13636 28908 13688 28917
rect 14188 28951 14240 28960
rect 14188 28917 14197 28951
rect 14197 28917 14231 28951
rect 14231 28917 14240 28951
rect 14188 28908 14240 28917
rect 2663 28806 2715 28858
rect 2727 28806 2779 28858
rect 2791 28806 2843 28858
rect 2855 28806 2907 28858
rect 2919 28806 2971 28858
rect 6090 28806 6142 28858
rect 6154 28806 6206 28858
rect 6218 28806 6270 28858
rect 6282 28806 6334 28858
rect 6346 28806 6398 28858
rect 9517 28806 9569 28858
rect 9581 28806 9633 28858
rect 9645 28806 9697 28858
rect 9709 28806 9761 28858
rect 9773 28806 9825 28858
rect 12944 28806 12996 28858
rect 13008 28806 13060 28858
rect 13072 28806 13124 28858
rect 13136 28806 13188 28858
rect 13200 28806 13252 28858
rect 5540 28704 5592 28756
rect 6000 28704 6052 28756
rect 8024 28704 8076 28756
rect 10784 28704 10836 28756
rect 8760 28636 8812 28688
rect 10140 28636 10192 28688
rect 9680 28568 9732 28620
rect 10324 28568 10376 28620
rect 12256 28704 12308 28756
rect 12624 28704 12676 28756
rect 13820 28704 13872 28756
rect 12348 28679 12400 28688
rect 12348 28645 12357 28679
rect 12357 28645 12391 28679
rect 12391 28645 12400 28679
rect 12348 28636 12400 28645
rect 756 28500 808 28552
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 3792 28364 3844 28416
rect 8852 28500 8904 28552
rect 7104 28364 7156 28416
rect 10692 28543 10744 28552
rect 10692 28509 10701 28543
rect 10701 28509 10735 28543
rect 10735 28509 10744 28543
rect 10692 28500 10744 28509
rect 10784 28543 10836 28552
rect 10784 28509 10818 28543
rect 10818 28509 10836 28543
rect 10784 28500 10836 28509
rect 10968 28543 11020 28552
rect 10968 28509 10977 28543
rect 10977 28509 11011 28543
rect 11011 28509 11020 28543
rect 10968 28500 11020 28509
rect 12072 28500 12124 28552
rect 12624 28543 12676 28552
rect 12624 28509 12633 28543
rect 12633 28509 12667 28543
rect 12667 28509 12676 28543
rect 12624 28500 12676 28509
rect 12900 28543 12952 28552
rect 12900 28509 12909 28543
rect 12909 28509 12943 28543
rect 12943 28509 12952 28543
rect 12900 28500 12952 28509
rect 13544 28500 13596 28552
rect 14004 28500 14056 28552
rect 14372 28500 14424 28552
rect 14556 28500 14608 28552
rect 12348 28364 12400 28416
rect 13820 28407 13872 28416
rect 13820 28373 13829 28407
rect 13829 28373 13863 28407
rect 13863 28373 13872 28407
rect 13820 28364 13872 28373
rect 14372 28407 14424 28416
rect 14372 28373 14381 28407
rect 14381 28373 14415 28407
rect 14415 28373 14424 28407
rect 14372 28364 14424 28373
rect 4376 28262 4428 28314
rect 4440 28262 4492 28314
rect 4504 28262 4556 28314
rect 4568 28262 4620 28314
rect 4632 28262 4684 28314
rect 7803 28262 7855 28314
rect 7867 28262 7919 28314
rect 7931 28262 7983 28314
rect 7995 28262 8047 28314
rect 8059 28262 8111 28314
rect 11230 28262 11282 28314
rect 11294 28262 11346 28314
rect 11358 28262 11410 28314
rect 11422 28262 11474 28314
rect 11486 28262 11538 28314
rect 14657 28262 14709 28314
rect 14721 28262 14773 28314
rect 14785 28262 14837 28314
rect 14849 28262 14901 28314
rect 14913 28262 14965 28314
rect 1584 28160 1636 28212
rect 1952 28160 2004 28212
rect 10140 28160 10192 28212
rect 10508 28160 10560 28212
rect 10968 28160 11020 28212
rect 11704 28160 11756 28212
rect 9772 28092 9824 28144
rect 10876 28092 10928 28144
rect 1492 28067 1544 28076
rect 1492 28033 1501 28067
rect 1501 28033 1535 28067
rect 1535 28033 1544 28067
rect 1492 28024 1544 28033
rect 7564 28024 7616 28076
rect 8208 28024 8260 28076
rect 1676 27820 1728 27872
rect 6644 27820 6696 27872
rect 8392 27820 8444 27872
rect 9128 27820 9180 27872
rect 9864 28024 9916 28076
rect 11980 28097 12032 28144
rect 11980 28092 12005 28097
rect 12005 28092 12032 28097
rect 12900 28160 12952 28212
rect 14280 28160 14332 28212
rect 13912 28135 13964 28144
rect 13912 28101 13921 28135
rect 13921 28101 13955 28135
rect 13955 28101 13964 28135
rect 13912 28092 13964 28101
rect 12072 28024 12124 28076
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 12624 28024 12676 28076
rect 15108 27888 15160 27940
rect 10048 27820 10100 27872
rect 10508 27820 10560 27872
rect 12808 27820 12860 27872
rect 13636 27863 13688 27872
rect 13636 27829 13645 27863
rect 13645 27829 13679 27863
rect 13679 27829 13688 27863
rect 13636 27820 13688 27829
rect 14188 27863 14240 27872
rect 14188 27829 14197 27863
rect 14197 27829 14231 27863
rect 14231 27829 14240 27863
rect 14188 27820 14240 27829
rect 2663 27718 2715 27770
rect 2727 27718 2779 27770
rect 2791 27718 2843 27770
rect 2855 27718 2907 27770
rect 2919 27718 2971 27770
rect 6090 27718 6142 27770
rect 6154 27718 6206 27770
rect 6218 27718 6270 27770
rect 6282 27718 6334 27770
rect 6346 27718 6398 27770
rect 9517 27718 9569 27770
rect 9581 27718 9633 27770
rect 9645 27718 9697 27770
rect 9709 27718 9761 27770
rect 9773 27718 9825 27770
rect 12944 27718 12996 27770
rect 13008 27718 13060 27770
rect 13072 27718 13124 27770
rect 13136 27718 13188 27770
rect 13200 27718 13252 27770
rect 13544 27616 13596 27668
rect 6000 27412 6052 27464
rect 8208 27412 8260 27464
rect 10876 27412 10928 27464
rect 11796 27455 11848 27464
rect 11796 27421 11805 27455
rect 11805 27421 11839 27455
rect 11839 27421 11848 27455
rect 11796 27412 11848 27421
rect 9680 27344 9732 27396
rect 12072 27455 12124 27464
rect 12072 27421 12081 27455
rect 12081 27421 12115 27455
rect 12115 27421 12124 27455
rect 12072 27412 12124 27421
rect 12348 27455 12400 27464
rect 12348 27421 12357 27455
rect 12357 27421 12391 27455
rect 12391 27421 12400 27455
rect 12348 27412 12400 27421
rect 13084 27455 13136 27464
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 13452 27412 13504 27464
rect 14096 27412 14148 27464
rect 6460 27276 6512 27328
rect 7196 27276 7248 27328
rect 8576 27276 8628 27328
rect 9772 27276 9824 27328
rect 11980 27276 12032 27328
rect 13636 27344 13688 27396
rect 13912 27387 13964 27396
rect 13912 27353 13921 27387
rect 13921 27353 13955 27387
rect 13955 27353 13964 27387
rect 13912 27344 13964 27353
rect 12624 27319 12676 27328
rect 12624 27285 12633 27319
rect 12633 27285 12667 27319
rect 12667 27285 12676 27319
rect 12624 27276 12676 27285
rect 12900 27319 12952 27328
rect 12900 27285 12909 27319
rect 12909 27285 12943 27319
rect 12943 27285 12952 27319
rect 12900 27276 12952 27285
rect 13728 27276 13780 27328
rect 4376 27174 4428 27226
rect 4440 27174 4492 27226
rect 4504 27174 4556 27226
rect 4568 27174 4620 27226
rect 4632 27174 4684 27226
rect 7803 27174 7855 27226
rect 7867 27174 7919 27226
rect 7931 27174 7983 27226
rect 7995 27174 8047 27226
rect 8059 27174 8111 27226
rect 11230 27174 11282 27226
rect 11294 27174 11346 27226
rect 11358 27174 11410 27226
rect 11422 27174 11474 27226
rect 11486 27174 11538 27226
rect 14657 27174 14709 27226
rect 14721 27174 14773 27226
rect 14785 27174 14837 27226
rect 14849 27174 14901 27226
rect 14913 27174 14965 27226
rect 5540 27072 5592 27124
rect 8300 27072 8352 27124
rect 9680 27072 9732 27124
rect 11060 27072 11112 27124
rect 11980 27072 12032 27124
rect 12348 27072 12400 27124
rect 12624 27072 12676 27124
rect 12900 27072 12952 27124
rect 756 26936 808 26988
rect 6736 26936 6788 26988
rect 1860 26732 1912 26784
rect 7196 26868 7248 26920
rect 7564 26911 7616 26920
rect 7564 26877 7573 26911
rect 7573 26877 7607 26911
rect 7607 26877 7616 26911
rect 7564 26868 7616 26877
rect 7748 26868 7800 26920
rect 7840 26911 7892 26920
rect 7840 26877 7849 26911
rect 7849 26877 7883 26911
rect 7883 26877 7892 26911
rect 7840 26868 7892 26877
rect 8760 26911 8812 26920
rect 8760 26877 8769 26911
rect 8769 26877 8803 26911
rect 8803 26877 8812 26911
rect 8760 26868 8812 26877
rect 9772 26979 9824 26988
rect 9772 26945 9781 26979
rect 9781 26945 9815 26979
rect 9815 26945 9824 26979
rect 9772 26936 9824 26945
rect 9036 26800 9088 26852
rect 9220 26911 9272 26920
rect 9220 26877 9229 26911
rect 9229 26877 9263 26911
rect 9263 26877 9272 26911
rect 9220 26868 9272 26877
rect 9588 26911 9640 26920
rect 9588 26877 9622 26911
rect 9622 26877 9640 26911
rect 12164 26936 12216 26988
rect 13084 27072 13136 27124
rect 14924 27072 14976 27124
rect 13452 27004 13504 27056
rect 14464 27004 14516 27056
rect 9588 26868 9640 26877
rect 12348 26868 12400 26920
rect 14004 26936 14056 26988
rect 6828 26732 6880 26784
rect 7656 26732 7708 26784
rect 7748 26732 7800 26784
rect 8944 26732 8996 26784
rect 9588 26732 9640 26784
rect 12348 26732 12400 26784
rect 13268 26775 13320 26784
rect 13268 26741 13277 26775
rect 13277 26741 13311 26775
rect 13311 26741 13320 26775
rect 13268 26732 13320 26741
rect 13820 26775 13872 26784
rect 13820 26741 13829 26775
rect 13829 26741 13863 26775
rect 13863 26741 13872 26775
rect 13820 26732 13872 26741
rect 15292 26732 15344 26784
rect 2663 26630 2715 26682
rect 2727 26630 2779 26682
rect 2791 26630 2843 26682
rect 2855 26630 2907 26682
rect 2919 26630 2971 26682
rect 6090 26630 6142 26682
rect 6154 26630 6206 26682
rect 6218 26630 6270 26682
rect 6282 26630 6334 26682
rect 6346 26630 6398 26682
rect 9517 26630 9569 26682
rect 9581 26630 9633 26682
rect 9645 26630 9697 26682
rect 9709 26630 9761 26682
rect 9773 26630 9825 26682
rect 12944 26630 12996 26682
rect 13008 26630 13060 26682
rect 13072 26630 13124 26682
rect 13136 26630 13188 26682
rect 13200 26630 13252 26682
rect 7840 26528 7892 26580
rect 9956 26528 10008 26580
rect 7564 26460 7616 26512
rect 8852 26460 8904 26512
rect 11152 26460 11204 26512
rect 11704 26528 11756 26580
rect 13728 26528 13780 26580
rect 1860 26324 1912 26376
rect 5448 26324 5500 26376
rect 6000 26324 6052 26376
rect 6368 26324 6420 26376
rect 6736 26367 6788 26376
rect 1492 26299 1544 26308
rect 1492 26265 1501 26299
rect 1501 26265 1535 26299
rect 1535 26265 1544 26299
rect 1492 26256 1544 26265
rect 6736 26333 6745 26367
rect 6745 26333 6788 26367
rect 6736 26324 6788 26333
rect 10048 26324 10100 26376
rect 7564 26256 7616 26308
rect 8576 26256 8628 26308
rect 13544 26324 13596 26376
rect 4068 26188 4120 26240
rect 8484 26188 8536 26240
rect 10968 26188 11020 26240
rect 12716 26188 12768 26240
rect 13636 26231 13688 26240
rect 13636 26197 13645 26231
rect 13645 26197 13679 26231
rect 13679 26197 13688 26231
rect 13636 26188 13688 26197
rect 14372 26231 14424 26240
rect 14372 26197 14381 26231
rect 14381 26197 14415 26231
rect 14415 26197 14424 26231
rect 14372 26188 14424 26197
rect 4376 26086 4428 26138
rect 4440 26086 4492 26138
rect 4504 26086 4556 26138
rect 4568 26086 4620 26138
rect 4632 26086 4684 26138
rect 7803 26086 7855 26138
rect 7867 26086 7919 26138
rect 7931 26086 7983 26138
rect 7995 26086 8047 26138
rect 8059 26086 8111 26138
rect 11230 26086 11282 26138
rect 11294 26086 11346 26138
rect 11358 26086 11410 26138
rect 11422 26086 11474 26138
rect 11486 26086 11538 26138
rect 14657 26086 14709 26138
rect 14721 26086 14773 26138
rect 14785 26086 14837 26138
rect 14849 26086 14901 26138
rect 14913 26086 14965 26138
rect 6644 25984 6696 26036
rect 7196 25848 7248 25900
rect 8208 25984 8260 26036
rect 9956 25984 10008 26036
rect 12440 25984 12492 26036
rect 8300 25891 8352 25900
rect 8300 25857 8307 25891
rect 8307 25857 8341 25891
rect 8341 25857 8352 25891
rect 9864 25916 9916 25968
rect 10140 25916 10192 25968
rect 8300 25848 8352 25857
rect 11704 25916 11756 25968
rect 13452 25916 13504 25968
rect 10692 25848 10744 25900
rect 6368 25823 6420 25832
rect 6368 25789 6377 25823
rect 6377 25789 6411 25823
rect 6411 25789 6420 25823
rect 6368 25780 6420 25789
rect 11152 25780 11204 25832
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 13360 25848 13412 25900
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 12440 25780 12492 25789
rect 12532 25823 12584 25832
rect 12532 25789 12566 25823
rect 12566 25789 12584 25823
rect 12532 25780 12584 25789
rect 15108 25780 15160 25832
rect 6644 25644 6696 25696
rect 7380 25687 7432 25696
rect 7380 25653 7389 25687
rect 7389 25653 7423 25687
rect 7423 25653 7432 25687
rect 7380 25644 7432 25653
rect 9220 25644 9272 25696
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 11980 25644 12032 25696
rect 12532 25644 12584 25696
rect 13820 25687 13872 25696
rect 13820 25653 13829 25687
rect 13829 25653 13863 25687
rect 13863 25653 13872 25687
rect 13820 25644 13872 25653
rect 15108 25644 15160 25696
rect 2663 25542 2715 25594
rect 2727 25542 2779 25594
rect 2791 25542 2843 25594
rect 2855 25542 2907 25594
rect 2919 25542 2971 25594
rect 6090 25542 6142 25594
rect 6154 25542 6206 25594
rect 6218 25542 6270 25594
rect 6282 25542 6334 25594
rect 6346 25542 6398 25594
rect 9517 25542 9569 25594
rect 9581 25542 9633 25594
rect 9645 25542 9697 25594
rect 9709 25542 9761 25594
rect 9773 25542 9825 25594
rect 12944 25542 12996 25594
rect 13008 25542 13060 25594
rect 13072 25542 13124 25594
rect 13136 25542 13188 25594
rect 13200 25542 13252 25594
rect 15292 25508 15344 25560
rect 6368 25440 6420 25492
rect 7380 25440 7432 25492
rect 9956 25440 10008 25492
rect 11060 25440 11112 25492
rect 12440 25440 12492 25492
rect 12808 25440 12860 25492
rect 756 25236 808 25288
rect 5448 25236 5500 25288
rect 5724 25236 5776 25288
rect 5816 25279 5868 25288
rect 5816 25245 5825 25279
rect 5825 25245 5859 25279
rect 5859 25245 5868 25279
rect 5816 25236 5868 25245
rect 6552 25279 6604 25288
rect 6552 25245 6561 25279
rect 6561 25245 6595 25279
rect 6595 25245 6604 25279
rect 6552 25236 6604 25245
rect 6736 25236 6788 25288
rect 9956 25236 10008 25288
rect 10508 25236 10560 25288
rect 10968 25236 11020 25288
rect 11704 25236 11756 25288
rect 11980 25236 12032 25288
rect 13636 25304 13688 25356
rect 7380 25168 7432 25220
rect 8668 25168 8720 25220
rect 12900 25279 12952 25288
rect 12900 25245 12934 25279
rect 12934 25245 12952 25279
rect 12900 25236 12952 25245
rect 13728 25236 13780 25288
rect 13820 25168 13872 25220
rect 15568 25168 15620 25220
rect 6644 25100 6696 25152
rect 6736 25100 6788 25152
rect 10692 25100 10744 25152
rect 10876 25100 10928 25152
rect 14372 25143 14424 25152
rect 14372 25109 14381 25143
rect 14381 25109 14415 25143
rect 14415 25109 14424 25143
rect 14372 25100 14424 25109
rect 4376 24998 4428 25050
rect 4440 24998 4492 25050
rect 4504 24998 4556 25050
rect 4568 24998 4620 25050
rect 4632 24998 4684 25050
rect 7803 24998 7855 25050
rect 7867 24998 7919 25050
rect 7931 24998 7983 25050
rect 7995 24998 8047 25050
rect 8059 24998 8111 25050
rect 11230 24998 11282 25050
rect 11294 24998 11346 25050
rect 11358 24998 11410 25050
rect 11422 24998 11474 25050
rect 11486 24998 11538 25050
rect 14657 24998 14709 25050
rect 14721 24998 14773 25050
rect 14785 24998 14837 25050
rect 14849 24998 14901 25050
rect 14913 24998 14965 25050
rect 10140 24896 10192 24948
rect 7564 24828 7616 24880
rect 756 24760 808 24812
rect 7380 24760 7432 24812
rect 6000 24692 6052 24744
rect 7564 24692 7616 24744
rect 9220 24803 9272 24812
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 8576 24692 8628 24744
rect 9128 24692 9180 24744
rect 9404 24692 9456 24744
rect 9772 24692 9824 24744
rect 8760 24624 8812 24676
rect 12072 24803 12124 24812
rect 12072 24769 12081 24803
rect 12081 24769 12115 24803
rect 12115 24769 12124 24803
rect 12072 24760 12124 24769
rect 12440 24803 12492 24812
rect 12440 24769 12447 24803
rect 12447 24769 12481 24803
rect 12481 24769 12492 24803
rect 12440 24760 12492 24769
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 8484 24556 8536 24608
rect 9128 24556 9180 24608
rect 9220 24556 9272 24608
rect 10876 24556 10928 24608
rect 11152 24556 11204 24608
rect 11520 24556 11572 24608
rect 13268 24556 13320 24608
rect 13360 24556 13412 24608
rect 15660 24760 15712 24812
rect 14280 24692 14332 24744
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 2663 24454 2715 24506
rect 2727 24454 2779 24506
rect 2791 24454 2843 24506
rect 2855 24454 2907 24506
rect 2919 24454 2971 24506
rect 6090 24454 6142 24506
rect 6154 24454 6206 24506
rect 6218 24454 6270 24506
rect 6282 24454 6334 24506
rect 6346 24454 6398 24506
rect 9517 24454 9569 24506
rect 9581 24454 9633 24506
rect 9645 24454 9697 24506
rect 9709 24454 9761 24506
rect 9773 24454 9825 24506
rect 12944 24454 12996 24506
rect 13008 24454 13060 24506
rect 13072 24454 13124 24506
rect 13136 24454 13188 24506
rect 13200 24454 13252 24506
rect 6000 24352 6052 24404
rect 7196 24352 7248 24404
rect 9956 24352 10008 24404
rect 10140 24352 10192 24404
rect 10416 24352 10468 24404
rect 8760 24284 8812 24336
rect 9220 24284 9272 24336
rect 9772 24284 9824 24336
rect 6368 24216 6420 24268
rect 6644 24216 6696 24268
rect 6920 24216 6972 24268
rect 7104 24216 7156 24268
rect 6828 24148 6880 24200
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 10416 24216 10468 24268
rect 10692 24259 10744 24268
rect 10692 24225 10726 24259
rect 10726 24225 10744 24259
rect 10692 24216 10744 24225
rect 10876 24259 10928 24268
rect 10876 24225 10885 24259
rect 10885 24225 10919 24259
rect 10919 24225 10928 24259
rect 10876 24216 10928 24225
rect 11888 24352 11940 24404
rect 13452 24284 13504 24336
rect 8668 24080 8720 24132
rect 6644 24012 6696 24064
rect 8852 24012 8904 24064
rect 9772 24148 9824 24200
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 10600 24148 10652 24157
rect 11520 24216 11572 24268
rect 13636 24216 13688 24268
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11940 24191
rect 11888 24148 11940 24157
rect 13820 24148 13872 24200
rect 13728 24080 13780 24132
rect 15108 24080 15160 24132
rect 10968 24012 11020 24064
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 14372 24055 14424 24064
rect 14372 24021 14381 24055
rect 14381 24021 14415 24055
rect 14415 24021 14424 24055
rect 14372 24012 14424 24021
rect 4376 23910 4428 23962
rect 4440 23910 4492 23962
rect 4504 23910 4556 23962
rect 4568 23910 4620 23962
rect 4632 23910 4684 23962
rect 7803 23910 7855 23962
rect 7867 23910 7919 23962
rect 7931 23910 7983 23962
rect 7995 23910 8047 23962
rect 8059 23910 8111 23962
rect 11230 23910 11282 23962
rect 11294 23910 11346 23962
rect 11358 23910 11410 23962
rect 11422 23910 11474 23962
rect 11486 23910 11538 23962
rect 14657 23910 14709 23962
rect 14721 23910 14773 23962
rect 14785 23910 14837 23962
rect 14849 23910 14901 23962
rect 14913 23910 14965 23962
rect 4988 23808 5040 23860
rect 9864 23808 9916 23860
rect 10324 23808 10376 23860
rect 10692 23808 10744 23860
rect 12348 23808 12400 23860
rect 8116 23740 8168 23792
rect 8576 23740 8628 23792
rect 6460 23672 6512 23724
rect 756 23604 808 23656
rect 6920 23647 6972 23656
rect 6920 23613 6929 23647
rect 6929 23613 6963 23647
rect 6963 23613 6972 23647
rect 6920 23604 6972 23613
rect 13728 23740 13780 23792
rect 9128 23647 9180 23656
rect 9128 23613 9137 23647
rect 9137 23613 9171 23647
rect 9171 23613 9180 23647
rect 9128 23604 9180 23613
rect 9956 23604 10008 23656
rect 11980 23715 12032 23724
rect 11980 23681 11989 23715
rect 11989 23681 12023 23715
rect 12023 23681 12032 23715
rect 11980 23672 12032 23681
rect 13176 23715 13228 23724
rect 13176 23681 13185 23715
rect 13185 23681 13219 23715
rect 13219 23681 13228 23715
rect 13176 23672 13228 23681
rect 11704 23604 11756 23656
rect 12348 23604 12400 23656
rect 12624 23647 12676 23656
rect 12624 23613 12633 23647
rect 12633 23613 12667 23647
rect 12667 23613 12676 23647
rect 12624 23604 12676 23613
rect 12992 23647 13044 23656
rect 12992 23613 13026 23647
rect 13026 23613 13044 23647
rect 12992 23604 13044 23613
rect 7196 23468 7248 23520
rect 8208 23468 8260 23520
rect 9404 23468 9456 23520
rect 10876 23468 10928 23520
rect 13268 23468 13320 23520
rect 13360 23468 13412 23520
rect 14372 23511 14424 23520
rect 14372 23477 14381 23511
rect 14381 23477 14415 23511
rect 14415 23477 14424 23511
rect 14372 23468 14424 23477
rect 2663 23366 2715 23418
rect 2727 23366 2779 23418
rect 2791 23366 2843 23418
rect 2855 23366 2907 23418
rect 2919 23366 2971 23418
rect 6090 23366 6142 23418
rect 6154 23366 6206 23418
rect 6218 23366 6270 23418
rect 6282 23366 6334 23418
rect 6346 23366 6398 23418
rect 9517 23366 9569 23418
rect 9581 23366 9633 23418
rect 9645 23366 9697 23418
rect 9709 23366 9761 23418
rect 9773 23366 9825 23418
rect 12944 23366 12996 23418
rect 13008 23366 13060 23418
rect 13072 23366 13124 23418
rect 13136 23366 13188 23418
rect 13200 23366 13252 23418
rect 5448 23264 5500 23316
rect 6920 23264 6972 23316
rect 9128 23264 9180 23316
rect 9956 23264 10008 23316
rect 8484 23196 8536 23248
rect 6552 23171 6604 23180
rect 6552 23137 6561 23171
rect 6561 23137 6595 23171
rect 6595 23137 6604 23171
rect 6552 23128 6604 23137
rect 6736 23128 6788 23180
rect 4252 23103 4304 23112
rect 4252 23069 4261 23103
rect 4261 23069 4295 23103
rect 4295 23069 4304 23103
rect 4252 23060 4304 23069
rect 5172 23060 5224 23112
rect 756 22992 808 23044
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 5724 23060 5776 23112
rect 5816 23103 5868 23112
rect 5816 23069 5825 23103
rect 5825 23069 5859 23103
rect 5859 23069 5868 23103
rect 5816 23060 5868 23069
rect 6828 23103 6880 23112
rect 6828 23069 6837 23103
rect 6837 23069 6871 23103
rect 6871 23069 6880 23103
rect 6828 23060 6880 23069
rect 11152 23264 11204 23316
rect 13728 23264 13780 23316
rect 13636 23196 13688 23248
rect 14372 23239 14424 23248
rect 14372 23205 14381 23239
rect 14381 23205 14415 23239
rect 14415 23205 14424 23239
rect 14372 23196 14424 23205
rect 9128 23060 9180 23112
rect 9772 23093 9824 23112
rect 9772 23060 9779 23093
rect 9779 23060 9813 23093
rect 9813 23060 9824 23093
rect 11152 23103 11204 23112
rect 11152 23069 11159 23103
rect 11159 23069 11193 23103
rect 11193 23069 11204 23103
rect 11152 23060 11204 23069
rect 11796 23060 11848 23112
rect 12808 23060 12860 23112
rect 13360 23060 13412 23112
rect 13452 23060 13504 23112
rect 13636 23103 13688 23112
rect 13636 23069 13645 23103
rect 13645 23069 13679 23103
rect 13679 23069 13688 23103
rect 13636 23060 13688 23069
rect 14280 23060 14332 23112
rect 8484 22992 8536 23044
rect 10048 22992 10100 23044
rect 13912 22992 13964 23044
rect 15936 22992 15988 23044
rect 6920 22924 6972 22976
rect 8116 22924 8168 22976
rect 9588 22924 9640 22976
rect 10876 22924 10928 22976
rect 11888 22967 11940 22976
rect 11888 22933 11897 22967
rect 11897 22933 11931 22967
rect 11931 22933 11940 22967
rect 11888 22924 11940 22933
rect 15108 22924 15160 22976
rect 4376 22822 4428 22874
rect 4440 22822 4492 22874
rect 4504 22822 4556 22874
rect 4568 22822 4620 22874
rect 4632 22822 4684 22874
rect 7803 22822 7855 22874
rect 7867 22822 7919 22874
rect 7931 22822 7983 22874
rect 7995 22822 8047 22874
rect 8059 22822 8111 22874
rect 11230 22822 11282 22874
rect 11294 22822 11346 22874
rect 11358 22822 11410 22874
rect 11422 22822 11474 22874
rect 11486 22822 11538 22874
rect 14657 22822 14709 22874
rect 14721 22822 14773 22874
rect 14785 22822 14837 22874
rect 14849 22822 14901 22874
rect 14913 22822 14965 22874
rect 1584 22720 1636 22772
rect 10692 22720 10744 22772
rect 11152 22720 11204 22772
rect 13636 22720 13688 22772
rect 14280 22720 14332 22772
rect 5080 22584 5132 22636
rect 6000 22584 6052 22636
rect 7196 22584 7248 22636
rect 7564 22584 7616 22636
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 14096 22652 14148 22704
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 13728 22627 13780 22636
rect 13728 22593 13737 22627
rect 13737 22593 13771 22627
rect 13771 22593 13780 22627
rect 13728 22584 13780 22593
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 6644 22448 6696 22500
rect 8208 22516 8260 22568
rect 8576 22559 8628 22568
rect 8576 22525 8585 22559
rect 8585 22525 8619 22559
rect 8619 22525 8628 22559
rect 8576 22516 8628 22525
rect 8668 22559 8720 22568
rect 8668 22525 8702 22559
rect 8702 22525 8720 22559
rect 8668 22516 8720 22525
rect 14004 22516 14056 22568
rect 13360 22448 13412 22500
rect 5816 22380 5868 22432
rect 12624 22380 12676 22432
rect 14004 22380 14056 22432
rect 14924 22380 14976 22432
rect 2663 22278 2715 22330
rect 2727 22278 2779 22330
rect 2791 22278 2843 22330
rect 2855 22278 2907 22330
rect 2919 22278 2971 22330
rect 6090 22278 6142 22330
rect 6154 22278 6206 22330
rect 6218 22278 6270 22330
rect 6282 22278 6334 22330
rect 6346 22278 6398 22330
rect 9517 22278 9569 22330
rect 9581 22278 9633 22330
rect 9645 22278 9697 22330
rect 9709 22278 9761 22330
rect 9773 22278 9825 22330
rect 12944 22278 12996 22330
rect 13008 22278 13060 22330
rect 13072 22278 13124 22330
rect 13136 22278 13188 22330
rect 13200 22278 13252 22330
rect 6828 22176 6880 22228
rect 6920 22176 6972 22228
rect 9588 22176 9640 22228
rect 9956 22176 10008 22228
rect 10232 22108 10284 22160
rect 4252 22040 4304 22092
rect 5448 22083 5500 22092
rect 5448 22049 5457 22083
rect 5457 22049 5491 22083
rect 5491 22049 5500 22083
rect 5448 22040 5500 22049
rect 9680 22040 9732 22092
rect 10692 22176 10744 22228
rect 756 21904 808 21956
rect 3148 22015 3200 22024
rect 3148 21981 3157 22015
rect 3157 21981 3191 22015
rect 3191 21981 3200 22015
rect 3148 21972 3200 21981
rect 5632 21972 5684 22024
rect 6276 21972 6328 22024
rect 6460 21972 6512 22024
rect 6828 22015 6880 22024
rect 6828 21981 6837 22015
rect 6837 21981 6871 22015
rect 6871 21981 6880 22015
rect 6828 21972 6880 21981
rect 7012 21972 7064 22024
rect 9956 21972 10008 22024
rect 10048 21972 10100 22024
rect 9496 21904 9548 21956
rect 12072 22040 12124 22092
rect 13176 22176 13228 22228
rect 13544 22176 13596 22228
rect 14464 22176 14516 22228
rect 11704 21972 11756 22024
rect 11796 22015 11848 22024
rect 11796 21981 11805 22015
rect 11805 21981 11839 22015
rect 11839 21981 11848 22015
rect 11796 21972 11848 21981
rect 12900 21972 12952 22024
rect 12992 22015 13044 22024
rect 12992 21981 13001 22015
rect 13001 21981 13035 22015
rect 13035 21981 13044 22015
rect 12992 21972 13044 21981
rect 14096 22040 14148 22092
rect 15200 22040 15252 22092
rect 15292 22040 15344 22092
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 14004 21972 14056 22024
rect 15108 21904 15160 21956
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 8208 21836 8260 21888
rect 9588 21836 9640 21888
rect 12900 21836 12952 21888
rect 13084 21836 13136 21888
rect 14004 21836 14056 21888
rect 15844 21836 15896 21888
rect 4376 21734 4428 21786
rect 4440 21734 4492 21786
rect 4504 21734 4556 21786
rect 4568 21734 4620 21786
rect 4632 21734 4684 21786
rect 7803 21734 7855 21786
rect 7867 21734 7919 21786
rect 7931 21734 7983 21786
rect 7995 21734 8047 21786
rect 8059 21734 8111 21786
rect 11230 21734 11282 21786
rect 11294 21734 11346 21786
rect 11358 21734 11410 21786
rect 11422 21734 11474 21786
rect 11486 21734 11538 21786
rect 14657 21734 14709 21786
rect 14721 21734 14773 21786
rect 14785 21734 14837 21786
rect 14849 21734 14901 21786
rect 14913 21734 14965 21786
rect 15384 21700 15436 21752
rect 2688 21675 2740 21684
rect 2688 21641 2697 21675
rect 2697 21641 2731 21675
rect 2731 21641 2740 21675
rect 2688 21632 2740 21641
rect 3148 21632 3200 21684
rect 5080 21632 5132 21684
rect 5540 21632 5592 21684
rect 6552 21632 6604 21684
rect 8392 21632 8444 21684
rect 8484 21632 8536 21684
rect 4160 21564 4212 21616
rect 7196 21564 7248 21616
rect 7380 21564 7432 21616
rect 9404 21632 9456 21684
rect 9864 21632 9916 21684
rect 10140 21675 10192 21684
rect 10140 21641 10149 21675
rect 10149 21641 10183 21675
rect 10183 21641 10192 21675
rect 10140 21632 10192 21641
rect 12992 21632 13044 21684
rect 14280 21632 14332 21684
rect 14464 21632 14516 21684
rect 5632 21496 5684 21548
rect 6276 21428 6328 21480
rect 6828 21428 6880 21480
rect 2136 21360 2188 21412
rect 7380 21360 7432 21412
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 8484 21539 8536 21548
rect 8484 21505 8518 21539
rect 8518 21505 8536 21539
rect 8484 21496 8536 21505
rect 8668 21539 8720 21548
rect 8668 21505 8677 21539
rect 8677 21505 8711 21539
rect 8711 21505 8720 21539
rect 8668 21496 8720 21505
rect 9404 21496 9456 21548
rect 7564 21428 7616 21480
rect 8116 21471 8168 21480
rect 8116 21437 8125 21471
rect 8125 21437 8159 21471
rect 8159 21437 8168 21471
rect 8116 21428 8168 21437
rect 9956 21496 10008 21548
rect 10600 21496 10652 21548
rect 10692 21496 10744 21548
rect 12348 21496 12400 21548
rect 13084 21539 13136 21548
rect 13084 21505 13093 21539
rect 13093 21505 13127 21539
rect 13127 21505 13136 21539
rect 13084 21496 13136 21505
rect 13360 21496 13412 21548
rect 14096 21539 14148 21548
rect 14096 21505 14105 21539
rect 14105 21505 14139 21539
rect 14139 21505 14148 21539
rect 14096 21496 14148 21505
rect 14188 21428 14240 21480
rect 5448 21292 5500 21344
rect 9680 21292 9732 21344
rect 9864 21335 9916 21344
rect 9864 21301 9873 21335
rect 9873 21301 9907 21335
rect 9907 21301 9916 21335
rect 9864 21292 9916 21301
rect 11244 21292 11296 21344
rect 11704 21292 11756 21344
rect 12072 21292 12124 21344
rect 13820 21335 13872 21344
rect 13820 21301 13829 21335
rect 13829 21301 13863 21335
rect 13863 21301 13872 21335
rect 13820 21292 13872 21301
rect 2663 21190 2715 21242
rect 2727 21190 2779 21242
rect 2791 21190 2843 21242
rect 2855 21190 2907 21242
rect 2919 21190 2971 21242
rect 6090 21190 6142 21242
rect 6154 21190 6206 21242
rect 6218 21190 6270 21242
rect 6282 21190 6334 21242
rect 6346 21190 6398 21242
rect 9517 21190 9569 21242
rect 9581 21190 9633 21242
rect 9645 21190 9697 21242
rect 9709 21190 9761 21242
rect 9773 21190 9825 21242
rect 12944 21190 12996 21242
rect 13008 21190 13060 21242
rect 13072 21190 13124 21242
rect 13136 21190 13188 21242
rect 13200 21190 13252 21242
rect 5448 21088 5500 21140
rect 8668 21088 8720 21140
rect 9404 21020 9456 21072
rect 4160 20952 4212 21004
rect 5632 20952 5684 21004
rect 6920 20952 6972 21004
rect 756 20884 808 20936
rect 5816 20884 5868 20936
rect 7012 20884 7064 20936
rect 4252 20816 4304 20868
rect 6460 20816 6512 20868
rect 6644 20816 6696 20868
rect 9772 21088 9824 21140
rect 9864 21088 9916 21140
rect 10140 21020 10192 21072
rect 10876 21020 10928 21072
rect 11888 20952 11940 21004
rect 7380 20884 7432 20936
rect 8668 20816 8720 20868
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 9864 20927 9916 20936
rect 9864 20893 9873 20927
rect 9873 20893 9907 20927
rect 9907 20893 9916 20927
rect 9864 20884 9916 20893
rect 6736 20748 6788 20800
rect 7472 20748 7524 20800
rect 10324 20927 10376 20936
rect 10324 20893 10333 20927
rect 10333 20893 10367 20927
rect 10367 20893 10376 20927
rect 10324 20884 10376 20893
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 11244 20884 11296 20936
rect 12440 20927 12492 20936
rect 12440 20893 12449 20927
rect 12449 20893 12483 20927
rect 12483 20893 12492 20927
rect 12440 20884 12492 20893
rect 12624 20884 12676 20936
rect 15108 21088 15160 21140
rect 10876 20748 10928 20800
rect 11244 20748 11296 20800
rect 11888 20748 11940 20800
rect 13544 20748 13596 20800
rect 14188 20748 14240 20800
rect 4376 20646 4428 20698
rect 4440 20646 4492 20698
rect 4504 20646 4556 20698
rect 4568 20646 4620 20698
rect 4632 20646 4684 20698
rect 7803 20646 7855 20698
rect 7867 20646 7919 20698
rect 7931 20646 7983 20698
rect 7995 20646 8047 20698
rect 8059 20646 8111 20698
rect 11230 20646 11282 20698
rect 11294 20646 11346 20698
rect 11358 20646 11410 20698
rect 11422 20646 11474 20698
rect 11486 20646 11538 20698
rect 14657 20646 14709 20698
rect 14721 20646 14773 20698
rect 14785 20646 14837 20698
rect 14849 20646 14901 20698
rect 14913 20646 14965 20698
rect 6552 20544 6604 20596
rect 7104 20544 7156 20596
rect 7380 20544 7432 20596
rect 8668 20544 8720 20596
rect 9864 20544 9916 20596
rect 13360 20544 13412 20596
rect 14096 20544 14148 20596
rect 756 20408 808 20460
rect 4252 20408 4304 20460
rect 5632 20408 5684 20460
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 6736 20476 6788 20528
rect 11520 20476 11572 20528
rect 12440 20476 12492 20528
rect 7288 20408 7340 20460
rect 6828 20383 6880 20392
rect 6828 20349 6837 20383
rect 6837 20349 6871 20383
rect 6871 20349 6880 20383
rect 6828 20340 6880 20349
rect 7012 20272 7064 20324
rect 11244 20408 11296 20460
rect 12164 20451 12216 20460
rect 12164 20417 12173 20451
rect 12173 20417 12207 20451
rect 12207 20417 12216 20451
rect 12164 20408 12216 20417
rect 12256 20408 12308 20460
rect 11980 20340 12032 20392
rect 12440 20340 12492 20392
rect 12072 20272 12124 20324
rect 7564 20204 7616 20256
rect 12440 20204 12492 20256
rect 12716 20408 12768 20460
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 14464 20451 14516 20460
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 13360 20383 13412 20392
rect 13360 20349 13394 20383
rect 13394 20349 13412 20383
rect 13360 20340 13412 20349
rect 12716 20272 12768 20324
rect 2663 20102 2715 20154
rect 2727 20102 2779 20154
rect 2791 20102 2843 20154
rect 2855 20102 2907 20154
rect 2919 20102 2971 20154
rect 6090 20102 6142 20154
rect 6154 20102 6206 20154
rect 6218 20102 6270 20154
rect 6282 20102 6334 20154
rect 6346 20102 6398 20154
rect 9517 20102 9569 20154
rect 9581 20102 9633 20154
rect 9645 20102 9697 20154
rect 9709 20102 9761 20154
rect 9773 20102 9825 20154
rect 12944 20102 12996 20154
rect 13008 20102 13060 20154
rect 13072 20102 13124 20154
rect 13136 20102 13188 20154
rect 13200 20102 13252 20154
rect 6000 20000 6052 20052
rect 6368 20043 6420 20052
rect 6368 20009 6377 20043
rect 6377 20009 6411 20043
rect 6411 20009 6420 20043
rect 6368 20000 6420 20009
rect 6828 20000 6880 20052
rect 7012 20000 7064 20052
rect 756 19728 808 19780
rect 5724 19796 5776 19848
rect 6092 19796 6144 19848
rect 6368 19796 6420 19848
rect 6552 19839 6604 19848
rect 6552 19805 6553 19839
rect 6553 19805 6587 19839
rect 6587 19805 6604 19839
rect 6552 19796 6604 19805
rect 6736 19796 6788 19848
rect 7104 19796 7156 19848
rect 9128 20000 9180 20052
rect 9772 20000 9824 20052
rect 9312 19809 9364 19848
rect 9312 19796 9337 19809
rect 9337 19796 9364 19809
rect 3332 19660 3384 19712
rect 5632 19660 5684 19712
rect 6000 19660 6052 19712
rect 7104 19660 7156 19712
rect 8668 19660 8720 19712
rect 8944 19660 8996 19712
rect 11796 20000 11848 20052
rect 11520 19864 11572 19916
rect 12440 20000 12492 20052
rect 12716 20043 12768 20052
rect 12716 20009 12725 20043
rect 12725 20009 12759 20043
rect 12759 20009 12768 20043
rect 12716 20000 12768 20009
rect 13728 20000 13780 20052
rect 15108 20000 15160 20052
rect 15568 20000 15620 20052
rect 13820 19932 13872 19984
rect 14004 19932 14056 19984
rect 13268 19864 13320 19916
rect 11888 19796 11940 19848
rect 12348 19796 12400 19848
rect 14004 19796 14056 19848
rect 14188 19839 14240 19848
rect 14188 19805 14197 19839
rect 14197 19805 14231 19839
rect 14231 19805 14240 19839
rect 14188 19796 14240 19805
rect 14648 19728 14700 19780
rect 10048 19703 10100 19712
rect 10048 19669 10057 19703
rect 10057 19669 10091 19703
rect 10091 19669 10100 19703
rect 10048 19660 10100 19669
rect 14188 19660 14240 19712
rect 14464 19660 14516 19712
rect 4376 19558 4428 19610
rect 4440 19558 4492 19610
rect 4504 19558 4556 19610
rect 4568 19558 4620 19610
rect 4632 19558 4684 19610
rect 7803 19558 7855 19610
rect 7867 19558 7919 19610
rect 7931 19558 7983 19610
rect 7995 19558 8047 19610
rect 8059 19558 8111 19610
rect 11230 19558 11282 19610
rect 11294 19558 11346 19610
rect 11358 19558 11410 19610
rect 11422 19558 11474 19610
rect 11486 19558 11538 19610
rect 14657 19558 14709 19610
rect 14721 19558 14773 19610
rect 14785 19558 14837 19610
rect 14849 19558 14901 19610
rect 14913 19558 14965 19610
rect 5172 19456 5224 19508
rect 6920 19456 6972 19508
rect 9312 19456 9364 19508
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 5724 19320 5776 19372
rect 4068 19252 4120 19304
rect 5540 19252 5592 19304
rect 6092 19363 6144 19372
rect 6092 19329 6101 19363
rect 6101 19329 6135 19363
rect 6135 19329 6144 19363
rect 6092 19320 6144 19329
rect 8392 19388 8444 19440
rect 8760 19388 8812 19440
rect 12164 19456 12216 19508
rect 14096 19456 14148 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 9128 19320 9180 19372
rect 9864 19320 9916 19372
rect 13636 19388 13688 19440
rect 6644 19252 6696 19304
rect 6828 19252 6880 19304
rect 7748 19252 7800 19304
rect 3424 19116 3476 19168
rect 4252 19116 4304 19168
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 9680 19184 9732 19236
rect 8208 19116 8260 19168
rect 9036 19116 9088 19168
rect 10048 19252 10100 19304
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 10508 19295 10560 19304
rect 10508 19261 10542 19295
rect 10542 19261 10560 19295
rect 10508 19252 10560 19261
rect 10692 19295 10744 19304
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 10508 19116 10560 19168
rect 11428 19116 11480 19168
rect 12440 19320 12492 19372
rect 12348 19252 12400 19304
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12624 19116 12676 19125
rect 14464 19184 14516 19236
rect 2663 19014 2715 19066
rect 2727 19014 2779 19066
rect 2791 19014 2843 19066
rect 2855 19014 2907 19066
rect 2919 19014 2971 19066
rect 6090 19014 6142 19066
rect 6154 19014 6206 19066
rect 6218 19014 6270 19066
rect 6282 19014 6334 19066
rect 6346 19014 6398 19066
rect 9517 19014 9569 19066
rect 9581 19014 9633 19066
rect 9645 19014 9697 19066
rect 9709 19014 9761 19066
rect 9773 19014 9825 19066
rect 12944 19014 12996 19066
rect 13008 19014 13060 19066
rect 13072 19014 13124 19066
rect 13136 19014 13188 19066
rect 13200 19014 13252 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 5724 18912 5776 18964
rect 7564 18912 7616 18964
rect 5632 18844 5684 18896
rect 756 18708 808 18760
rect 10692 18912 10744 18964
rect 11152 18912 11204 18964
rect 11796 18912 11848 18964
rect 12256 18912 12308 18964
rect 13636 18844 13688 18896
rect 13912 18844 13964 18896
rect 5816 18751 5868 18760
rect 5816 18717 5825 18751
rect 5825 18717 5859 18751
rect 5859 18717 5868 18751
rect 5816 18708 5868 18717
rect 4804 18640 4856 18692
rect 6184 18640 6236 18692
rect 5632 18572 5684 18624
rect 6000 18615 6052 18624
rect 6000 18581 6009 18615
rect 6009 18581 6043 18615
rect 6043 18581 6052 18615
rect 6000 18572 6052 18581
rect 6092 18572 6144 18624
rect 6828 18708 6880 18760
rect 7380 18708 7432 18760
rect 9864 18776 9916 18828
rect 11428 18776 11480 18828
rect 7656 18708 7708 18760
rect 9036 18708 9088 18760
rect 9312 18751 9364 18760
rect 9312 18717 9321 18751
rect 9321 18717 9355 18751
rect 9355 18717 9364 18751
rect 9312 18708 9364 18717
rect 10140 18708 10192 18760
rect 7380 18572 7432 18624
rect 7748 18572 7800 18624
rect 8944 18572 8996 18624
rect 10048 18572 10100 18624
rect 10600 18572 10652 18624
rect 12072 18708 12124 18760
rect 12716 18708 12768 18760
rect 13912 18751 13964 18760
rect 13912 18717 13921 18751
rect 13921 18717 13955 18751
rect 13955 18717 13964 18751
rect 13912 18708 13964 18717
rect 14464 18640 14516 18692
rect 15108 18640 15160 18692
rect 10784 18572 10836 18624
rect 13268 18572 13320 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 4376 18470 4428 18522
rect 4440 18470 4492 18522
rect 4504 18470 4556 18522
rect 4568 18470 4620 18522
rect 4632 18470 4684 18522
rect 7803 18470 7855 18522
rect 7867 18470 7919 18522
rect 7931 18470 7983 18522
rect 7995 18470 8047 18522
rect 8059 18470 8111 18522
rect 11230 18470 11282 18522
rect 11294 18470 11346 18522
rect 11358 18470 11410 18522
rect 11422 18470 11474 18522
rect 11486 18470 11538 18522
rect 14657 18470 14709 18522
rect 14721 18470 14773 18522
rect 14785 18470 14837 18522
rect 14849 18470 14901 18522
rect 14913 18470 14965 18522
rect 5540 18411 5592 18420
rect 5540 18377 5549 18411
rect 5549 18377 5583 18411
rect 5583 18377 5592 18411
rect 5540 18368 5592 18377
rect 5816 18411 5868 18420
rect 5816 18377 5825 18411
rect 5825 18377 5859 18411
rect 5859 18377 5868 18411
rect 5816 18368 5868 18377
rect 6000 18368 6052 18420
rect 6828 18368 6880 18420
rect 8760 18368 8812 18420
rect 9312 18368 9364 18420
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 4160 18275 4212 18284
rect 4160 18241 4169 18275
rect 4169 18241 4203 18275
rect 4203 18241 4212 18275
rect 4160 18232 4212 18241
rect 4436 18275 4488 18284
rect 4436 18241 4470 18275
rect 4470 18241 4488 18275
rect 4436 18232 4488 18241
rect 6736 18300 6788 18352
rect 7656 18300 7708 18352
rect 572 18164 624 18216
rect 2504 18096 2556 18148
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 9036 18275 9088 18284
rect 9036 18241 9045 18275
rect 9045 18241 9079 18275
rect 9079 18241 9088 18275
rect 9036 18232 9088 18241
rect 7380 18164 7432 18216
rect 7012 18096 7064 18148
rect 8208 18164 8260 18216
rect 10692 18300 10744 18352
rect 10784 18300 10836 18352
rect 10876 18300 10928 18352
rect 13360 18368 13412 18420
rect 14372 18368 14424 18420
rect 14648 18368 14700 18420
rect 15292 18368 15344 18420
rect 12164 18300 12216 18352
rect 13452 18300 13504 18352
rect 13820 18300 13872 18352
rect 9680 18275 9732 18284
rect 9680 18241 9689 18275
rect 9689 18241 9723 18275
rect 9723 18241 9732 18275
rect 9680 18232 9732 18241
rect 11244 18232 11296 18284
rect 11796 18275 11848 18284
rect 11796 18241 11803 18275
rect 11803 18241 11837 18275
rect 11837 18241 11848 18275
rect 11796 18232 11848 18241
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 14372 18232 14424 18284
rect 10784 18164 10836 18216
rect 10968 18096 11020 18148
rect 8208 18028 8260 18080
rect 10508 18028 10560 18080
rect 12440 18028 12492 18080
rect 12716 18028 12768 18080
rect 12808 18028 12860 18080
rect 13452 18028 13504 18080
rect 14188 18028 14240 18080
rect 2663 17926 2715 17978
rect 2727 17926 2779 17978
rect 2791 17926 2843 17978
rect 2855 17926 2907 17978
rect 2919 17926 2971 17978
rect 6090 17926 6142 17978
rect 6154 17926 6206 17978
rect 6218 17926 6270 17978
rect 6282 17926 6334 17978
rect 6346 17926 6398 17978
rect 9517 17926 9569 17978
rect 9581 17926 9633 17978
rect 9645 17926 9697 17978
rect 9709 17926 9761 17978
rect 9773 17926 9825 17978
rect 12944 17926 12996 17978
rect 13008 17926 13060 17978
rect 13072 17926 13124 17978
rect 13136 17926 13188 17978
rect 13200 17926 13252 17978
rect 10600 17824 10652 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 12532 17867 12584 17876
rect 12532 17833 12541 17867
rect 12541 17833 12575 17867
rect 12575 17833 12584 17867
rect 12532 17824 12584 17833
rect 13360 17824 13412 17876
rect 15108 17824 15160 17876
rect 15568 17824 15620 17876
rect 4896 17688 4948 17740
rect 5448 17688 5500 17740
rect 6184 17688 6236 17740
rect 3976 17620 4028 17672
rect 9772 17688 9824 17740
rect 10784 17731 10836 17740
rect 10784 17697 10793 17731
rect 10793 17697 10827 17731
rect 10827 17697 10836 17731
rect 10784 17688 10836 17697
rect 12072 17688 12124 17740
rect 12440 17688 12492 17740
rect 9312 17620 9364 17672
rect 9864 17620 9916 17672
rect 11060 17663 11112 17672
rect 4160 17552 4212 17604
rect 4436 17552 4488 17604
rect 5908 17595 5960 17604
rect 5908 17561 5917 17595
rect 5917 17561 5951 17595
rect 5951 17561 5960 17595
rect 5908 17552 5960 17561
rect 6552 17552 6604 17604
rect 6644 17595 6696 17604
rect 6644 17561 6653 17595
rect 6653 17561 6687 17595
rect 6687 17561 6696 17595
rect 6644 17552 6696 17561
rect 6828 17552 6880 17604
rect 11060 17629 11067 17663
rect 11067 17629 11101 17663
rect 11101 17629 11112 17663
rect 11060 17620 11112 17629
rect 13728 17756 13780 17808
rect 14280 17688 14332 17740
rect 12808 17620 12860 17672
rect 13084 17620 13136 17672
rect 11428 17552 11480 17604
rect 7012 17527 7064 17536
rect 7012 17493 7021 17527
rect 7021 17493 7055 17527
rect 7055 17493 7064 17527
rect 7012 17484 7064 17493
rect 9036 17484 9088 17536
rect 11060 17484 11112 17536
rect 11888 17552 11940 17604
rect 12072 17552 12124 17604
rect 14096 17620 14148 17672
rect 15844 17620 15896 17672
rect 14648 17552 14700 17604
rect 12164 17484 12216 17536
rect 4376 17382 4428 17434
rect 4440 17382 4492 17434
rect 4504 17382 4556 17434
rect 4568 17382 4620 17434
rect 4632 17382 4684 17434
rect 7803 17382 7855 17434
rect 7867 17382 7919 17434
rect 7931 17382 7983 17434
rect 7995 17382 8047 17434
rect 8059 17382 8111 17434
rect 11230 17382 11282 17434
rect 11294 17382 11346 17434
rect 11358 17382 11410 17434
rect 11422 17382 11474 17434
rect 11486 17382 11538 17434
rect 14657 17382 14709 17434
rect 14721 17382 14773 17434
rect 14785 17382 14837 17434
rect 14849 17382 14901 17434
rect 14913 17382 14965 17434
rect 756 17144 808 17196
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 5908 17280 5960 17332
rect 7564 17280 7616 17332
rect 7748 17280 7800 17332
rect 8668 17280 8720 17332
rect 5264 17144 5316 17196
rect 9036 17144 9088 17196
rect 9220 17144 9272 17196
rect 11980 17280 12032 17332
rect 15200 17280 15252 17332
rect 15292 17212 15344 17264
rect 15568 17212 15620 17264
rect 5632 17076 5684 17128
rect 6184 17076 6236 17128
rect 8852 17076 8904 17128
rect 4896 16940 4948 16992
rect 8300 17008 8352 17060
rect 7564 16940 7616 16992
rect 10140 17076 10192 17128
rect 10508 17076 10560 17128
rect 10600 17119 10652 17128
rect 10600 17085 10609 17119
rect 10609 17085 10643 17119
rect 10643 17085 10652 17119
rect 10600 17076 10652 17085
rect 11612 17076 11664 17128
rect 10048 17051 10100 17060
rect 10048 17017 10057 17051
rect 10057 17017 10091 17051
rect 10091 17017 10100 17051
rect 10048 17008 10100 17017
rect 10784 16940 10836 16992
rect 11244 16983 11296 16992
rect 11244 16949 11253 16983
rect 11253 16949 11287 16983
rect 11287 16949 11296 16983
rect 11244 16940 11296 16949
rect 12440 17187 12492 17196
rect 12440 17153 12449 17187
rect 12449 17153 12483 17187
rect 12483 17153 12492 17187
rect 12440 17144 12492 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 13544 17187 13596 17196
rect 13544 17153 13553 17187
rect 13553 17153 13587 17187
rect 13587 17153 13596 17187
rect 13544 17144 13596 17153
rect 13636 17144 13688 17196
rect 12164 17119 12216 17128
rect 12164 17085 12173 17119
rect 12173 17085 12207 17119
rect 12207 17085 12216 17119
rect 12164 17076 12216 17085
rect 12532 17076 12584 17128
rect 13084 17076 13136 17128
rect 11888 16940 11940 16992
rect 2663 16838 2715 16890
rect 2727 16838 2779 16890
rect 2791 16838 2843 16890
rect 2855 16838 2907 16890
rect 2919 16838 2971 16890
rect 6090 16838 6142 16890
rect 6154 16838 6206 16890
rect 6218 16838 6270 16890
rect 6282 16838 6334 16890
rect 6346 16838 6398 16890
rect 9517 16838 9569 16890
rect 9581 16838 9633 16890
rect 9645 16838 9697 16890
rect 9709 16838 9761 16890
rect 9773 16838 9825 16890
rect 12944 16838 12996 16890
rect 13008 16838 13060 16890
rect 13072 16838 13124 16890
rect 13136 16838 13188 16890
rect 13200 16838 13252 16890
rect 4896 16736 4948 16788
rect 6552 16779 6604 16788
rect 6552 16745 6561 16779
rect 6561 16745 6595 16779
rect 6595 16745 6604 16779
rect 6552 16736 6604 16745
rect 8300 16736 8352 16788
rect 9680 16736 9732 16788
rect 10600 16736 10652 16788
rect 12072 16736 12124 16788
rect 12716 16736 12768 16788
rect 8668 16668 8720 16720
rect 14188 16668 14240 16720
rect 5448 16600 5500 16652
rect 2504 16532 2556 16584
rect 5172 16532 5224 16584
rect 11888 16600 11940 16652
rect 12624 16600 12676 16652
rect 13084 16643 13136 16652
rect 13084 16609 13118 16643
rect 13118 16609 13136 16643
rect 13084 16600 13136 16609
rect 13268 16643 13320 16652
rect 13268 16609 13277 16643
rect 13277 16609 13311 16643
rect 13311 16609 13320 16643
rect 13268 16600 13320 16609
rect 756 16464 808 16516
rect 5632 16464 5684 16516
rect 6552 16532 6604 16584
rect 7104 16522 7156 16574
rect 9312 16532 9364 16584
rect 9680 16575 9732 16584
rect 9680 16541 9687 16575
rect 9687 16541 9721 16575
rect 9721 16541 9732 16575
rect 9680 16532 9732 16541
rect 11244 16532 11296 16584
rect 7748 16464 7800 16516
rect 10140 16464 10192 16516
rect 7104 16396 7156 16448
rect 9588 16396 9640 16448
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 12808 16396 12860 16448
rect 13820 16396 13872 16448
rect 4376 16294 4428 16346
rect 4440 16294 4492 16346
rect 4504 16294 4556 16346
rect 4568 16294 4620 16346
rect 4632 16294 4684 16346
rect 7803 16294 7855 16346
rect 7867 16294 7919 16346
rect 7931 16294 7983 16346
rect 7995 16294 8047 16346
rect 8059 16294 8111 16346
rect 11230 16294 11282 16346
rect 11294 16294 11346 16346
rect 11358 16294 11410 16346
rect 11422 16294 11474 16346
rect 11486 16294 11538 16346
rect 14657 16294 14709 16346
rect 14721 16294 14773 16346
rect 14785 16294 14837 16346
rect 14849 16294 14901 16346
rect 14913 16294 14965 16346
rect 7840 16192 7892 16244
rect 7104 16124 7156 16176
rect 9864 16124 9916 16176
rect 10048 16192 10100 16244
rect 12348 16235 12400 16244
rect 12348 16201 12357 16235
rect 12357 16201 12391 16235
rect 12391 16201 12400 16235
rect 12348 16192 12400 16201
rect 848 16056 900 16108
rect 7288 16056 7340 16108
rect 7564 15988 7616 16040
rect 7748 15988 7800 16040
rect 8392 16099 8444 16108
rect 8392 16065 8401 16099
rect 8401 16065 8435 16099
rect 8435 16065 8444 16099
rect 8392 16056 8444 16065
rect 8576 16056 8628 16108
rect 8668 16099 8720 16108
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 9588 16056 9640 16108
rect 8208 15988 8260 16040
rect 9312 15988 9364 16040
rect 12716 16056 12768 16108
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 2504 15852 2556 15904
rect 12808 15920 12860 15972
rect 13636 16031 13688 16040
rect 13636 15997 13670 16031
rect 13670 15997 13688 16031
rect 13636 15988 13688 15997
rect 9864 15852 9916 15904
rect 11612 15852 11664 15904
rect 13084 15852 13136 15904
rect 2663 15750 2715 15802
rect 2727 15750 2779 15802
rect 2791 15750 2843 15802
rect 2855 15750 2907 15802
rect 2919 15750 2971 15802
rect 6090 15750 6142 15802
rect 6154 15750 6206 15802
rect 6218 15750 6270 15802
rect 6282 15750 6334 15802
rect 6346 15750 6398 15802
rect 9517 15750 9569 15802
rect 9581 15750 9633 15802
rect 9645 15750 9697 15802
rect 9709 15750 9761 15802
rect 9773 15750 9825 15802
rect 12944 15750 12996 15802
rect 13008 15750 13060 15802
rect 13072 15750 13124 15802
rect 13136 15750 13188 15802
rect 13200 15750 13252 15802
rect 1308 15444 1360 15496
rect 2044 15444 2096 15496
rect 2504 15444 2556 15496
rect 5172 15444 5224 15496
rect 5448 15444 5500 15496
rect 5632 15648 5684 15700
rect 8392 15648 8444 15700
rect 11612 15580 11664 15632
rect 13268 15691 13320 15700
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 11796 15512 11848 15564
rect 6920 15444 6972 15496
rect 7288 15444 7340 15496
rect 8944 15444 8996 15496
rect 9312 15444 9364 15496
rect 9864 15444 9916 15496
rect 11980 15512 12032 15564
rect 2504 15308 2556 15360
rect 7196 15308 7248 15360
rect 8576 15376 8628 15428
rect 11796 15376 11848 15428
rect 10416 15308 10468 15360
rect 10692 15308 10744 15360
rect 10876 15308 10928 15360
rect 14832 15444 14884 15496
rect 12348 15376 12400 15428
rect 15108 15376 15160 15428
rect 13176 15308 13228 15360
rect 4376 15206 4428 15258
rect 4440 15206 4492 15258
rect 4504 15206 4556 15258
rect 4568 15206 4620 15258
rect 4632 15206 4684 15258
rect 7803 15206 7855 15258
rect 7867 15206 7919 15258
rect 7931 15206 7983 15258
rect 7995 15206 8047 15258
rect 8059 15206 8111 15258
rect 11230 15206 11282 15258
rect 11294 15206 11346 15258
rect 11358 15206 11410 15258
rect 11422 15206 11474 15258
rect 11486 15206 11538 15258
rect 14657 15206 14709 15258
rect 14721 15206 14773 15258
rect 14785 15206 14837 15258
rect 14849 15206 14901 15258
rect 14913 15206 14965 15258
rect 2044 14968 2096 15020
rect 1308 14900 1360 14952
rect 8576 15104 8628 15156
rect 7840 15011 7892 15020
rect 7840 14977 7849 15011
rect 7849 14977 7883 15011
rect 7883 14977 7892 15011
rect 7840 14968 7892 14977
rect 7196 14900 7248 14952
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 2412 14807 2464 14816
rect 2412 14773 2421 14807
rect 2421 14773 2455 14807
rect 2455 14773 2464 14807
rect 2412 14764 2464 14773
rect 7472 14832 7524 14884
rect 9312 14832 9364 14884
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10232 14900 10284 14952
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 13360 15104 13412 15156
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 11704 14968 11756 15020
rect 12348 14968 12400 15020
rect 12716 14968 12768 15020
rect 13728 15036 13780 15088
rect 14188 14968 14240 15020
rect 10508 14943 10560 14952
rect 10508 14909 10542 14943
rect 10542 14909 10560 14943
rect 10508 14900 10560 14909
rect 11980 14900 12032 14952
rect 10140 14875 10192 14884
rect 10140 14841 10149 14875
rect 10149 14841 10183 14875
rect 10183 14841 10192 14875
rect 10140 14832 10192 14841
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9220 14764 9272 14816
rect 12348 14764 12400 14816
rect 12900 14764 12952 14816
rect 2663 14662 2715 14714
rect 2727 14662 2779 14714
rect 2791 14662 2843 14714
rect 2855 14662 2907 14714
rect 2919 14662 2971 14714
rect 6090 14662 6142 14714
rect 6154 14662 6206 14714
rect 6218 14662 6270 14714
rect 6282 14662 6334 14714
rect 6346 14662 6398 14714
rect 9517 14662 9569 14714
rect 9581 14662 9633 14714
rect 9645 14662 9697 14714
rect 9709 14662 9761 14714
rect 9773 14662 9825 14714
rect 12944 14662 12996 14714
rect 13008 14662 13060 14714
rect 13072 14662 13124 14714
rect 13136 14662 13188 14714
rect 13200 14662 13252 14714
rect 848 14560 900 14612
rect 2412 14560 2464 14612
rect 3608 14560 3660 14612
rect 8116 14560 8168 14612
rect 8300 14560 8352 14612
rect 8576 14560 8628 14612
rect 8668 14492 8720 14544
rect 10140 14560 10192 14612
rect 12256 14560 12308 14612
rect 14004 14560 14056 14612
rect 13544 14492 13596 14544
rect 7840 14424 7892 14476
rect 13176 14424 13228 14476
rect 13636 14424 13688 14476
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 6368 14356 6420 14408
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 7196 14288 7248 14340
rect 7656 14288 7708 14340
rect 8392 14356 8444 14408
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 9220 14399 9272 14408
rect 8944 14356 8996 14365
rect 8576 14288 8628 14340
rect 9036 14288 9088 14340
rect 9220 14365 9229 14399
rect 9229 14365 9272 14399
rect 9220 14356 9272 14365
rect 10232 14356 10284 14408
rect 10048 14288 10100 14340
rect 10784 14220 10836 14272
rect 10968 14288 11020 14340
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12124 14399
rect 12072 14356 12124 14365
rect 11152 14288 11204 14340
rect 14832 14356 14884 14408
rect 14280 14331 14332 14340
rect 14280 14297 14289 14331
rect 14289 14297 14323 14331
rect 14323 14297 14332 14331
rect 14280 14288 14332 14297
rect 11704 14220 11756 14272
rect 12716 14220 12768 14272
rect 13452 14220 13504 14272
rect 13636 14220 13688 14272
rect 4376 14118 4428 14170
rect 4440 14118 4492 14170
rect 4504 14118 4556 14170
rect 4568 14118 4620 14170
rect 4632 14118 4684 14170
rect 7803 14118 7855 14170
rect 7867 14118 7919 14170
rect 7931 14118 7983 14170
rect 7995 14118 8047 14170
rect 8059 14118 8111 14170
rect 11230 14118 11282 14170
rect 11294 14118 11346 14170
rect 11358 14118 11410 14170
rect 11422 14118 11474 14170
rect 11486 14118 11538 14170
rect 14657 14118 14709 14170
rect 14721 14118 14773 14170
rect 14785 14118 14837 14170
rect 14849 14118 14901 14170
rect 14913 14118 14965 14170
rect 2044 14016 2096 14068
rect 6460 13948 6512 14000
rect 1860 13923 1912 13932
rect 1860 13889 1869 13923
rect 1869 13889 1903 13923
rect 1903 13889 1912 13923
rect 1860 13880 1912 13889
rect 5448 13880 5500 13932
rect 6368 13923 6420 13932
rect 6368 13889 6377 13923
rect 6377 13889 6411 13923
rect 6411 13889 6420 13923
rect 6368 13880 6420 13889
rect 6644 13923 6696 13932
rect 6644 13889 6651 13923
rect 6651 13889 6685 13923
rect 6685 13889 6696 13923
rect 6644 13880 6696 13889
rect 7104 13880 7156 13932
rect 7472 14016 7524 14068
rect 9220 14016 9272 14068
rect 11152 14016 11204 14068
rect 11704 14016 11756 14068
rect 12164 14016 12216 14068
rect 9956 13948 10008 14000
rect 7656 13812 7708 13864
rect 8208 13855 8260 13864
rect 8208 13821 8217 13855
rect 8217 13821 8251 13855
rect 8251 13821 8260 13855
rect 8208 13812 8260 13821
rect 8300 13812 8352 13864
rect 9036 13923 9088 13932
rect 9036 13889 9070 13923
rect 9070 13889 9088 13923
rect 9036 13880 9088 13889
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 10416 13880 10468 13932
rect 8944 13855 8996 13864
rect 8944 13821 8953 13855
rect 8953 13821 8987 13855
rect 8987 13821 8996 13855
rect 8944 13812 8996 13821
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10048 13812 10100 13821
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 13636 13948 13688 14000
rect 11704 13855 11756 13864
rect 11704 13821 11713 13855
rect 11713 13821 11747 13855
rect 11747 13821 11756 13855
rect 11704 13812 11756 13821
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 12256 13812 12308 13864
rect 12532 13855 12584 13864
rect 12532 13821 12566 13855
rect 12566 13821 12584 13855
rect 12532 13812 12584 13821
rect 13636 13855 13688 13864
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 13728 13812 13780 13864
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 2504 13719 2556 13728
rect 2504 13685 2513 13719
rect 2513 13685 2547 13719
rect 2547 13685 2556 13719
rect 2504 13676 2556 13685
rect 9036 13676 9088 13728
rect 11980 13744 12032 13796
rect 11428 13676 11480 13728
rect 13176 13676 13228 13728
rect 13360 13676 13412 13728
rect 2663 13574 2715 13626
rect 2727 13574 2779 13626
rect 2791 13574 2843 13626
rect 2855 13574 2907 13626
rect 2919 13574 2971 13626
rect 6090 13574 6142 13626
rect 6154 13574 6206 13626
rect 6218 13574 6270 13626
rect 6282 13574 6334 13626
rect 6346 13574 6398 13626
rect 9517 13574 9569 13626
rect 9581 13574 9633 13626
rect 9645 13574 9697 13626
rect 9709 13574 9761 13626
rect 9773 13574 9825 13626
rect 12944 13574 12996 13626
rect 13008 13574 13060 13626
rect 13072 13574 13124 13626
rect 13136 13574 13188 13626
rect 13200 13574 13252 13626
rect 1308 13268 1360 13320
rect 5448 13472 5500 13524
rect 7472 13472 7524 13524
rect 8392 13472 8444 13524
rect 8760 13472 8812 13524
rect 13912 13515 13964 13524
rect 13912 13481 13921 13515
rect 13921 13481 13955 13515
rect 13955 13481 13964 13515
rect 13912 13472 13964 13481
rect 14372 13472 14424 13524
rect 1676 13311 1728 13320
rect 1676 13277 1683 13311
rect 1683 13277 1717 13311
rect 1717 13277 1728 13311
rect 1676 13268 1728 13277
rect 2136 13268 2188 13320
rect 4252 13268 4304 13320
rect 5632 13268 5684 13320
rect 6092 13311 6144 13320
rect 6092 13277 6101 13311
rect 6101 13277 6135 13311
rect 6135 13277 6144 13311
rect 6092 13268 6144 13277
rect 6460 13268 6512 13320
rect 2504 13132 2556 13184
rect 6736 13200 6788 13252
rect 9496 13268 9548 13320
rect 10416 13268 10468 13320
rect 10232 13200 10284 13252
rect 7104 13175 7156 13184
rect 7104 13141 7113 13175
rect 7113 13141 7147 13175
rect 7147 13141 7156 13175
rect 7104 13132 7156 13141
rect 8760 13132 8812 13184
rect 10140 13132 10192 13184
rect 11520 13336 11572 13388
rect 12716 13379 12768 13388
rect 12716 13345 12725 13379
rect 12725 13345 12759 13379
rect 12759 13345 12768 13379
rect 12716 13336 12768 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 13084 13379 13136 13388
rect 13084 13345 13118 13379
rect 13118 13345 13136 13379
rect 13084 13336 13136 13345
rect 11796 13268 11848 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 12072 13268 12124 13277
rect 12164 13268 12216 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 15292 13336 15344 13388
rect 15844 13336 15896 13388
rect 10692 13175 10744 13184
rect 10692 13141 10701 13175
rect 10701 13141 10735 13175
rect 10735 13141 10744 13175
rect 10692 13132 10744 13141
rect 14464 13200 14516 13252
rect 4376 13030 4428 13082
rect 4440 13030 4492 13082
rect 4504 13030 4556 13082
rect 4568 13030 4620 13082
rect 4632 13030 4684 13082
rect 7803 13030 7855 13082
rect 7867 13030 7919 13082
rect 7931 13030 7983 13082
rect 7995 13030 8047 13082
rect 8059 13030 8111 13082
rect 11230 13030 11282 13082
rect 11294 13030 11346 13082
rect 11358 13030 11410 13082
rect 11422 13030 11474 13082
rect 11486 13030 11538 13082
rect 14657 13030 14709 13082
rect 14721 13030 14773 13082
rect 14785 13030 14837 13082
rect 14849 13030 14901 13082
rect 14913 13030 14965 13082
rect 1768 12928 1820 12980
rect 6736 12928 6788 12980
rect 7104 12928 7156 12980
rect 7564 12928 7616 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 1308 12724 1360 12776
rect 7656 12724 7708 12776
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8576 12835 8628 12844
rect 8576 12801 8610 12835
rect 8610 12801 8628 12835
rect 8576 12792 8628 12801
rect 8760 12835 8812 12844
rect 8760 12801 8769 12835
rect 8769 12801 8803 12835
rect 8803 12801 8812 12835
rect 8760 12792 8812 12801
rect 9772 12835 9824 12844
rect 9772 12801 9779 12835
rect 9779 12801 9813 12835
rect 9813 12801 9824 12835
rect 9772 12792 9824 12801
rect 11796 12835 11848 12844
rect 11796 12801 11805 12835
rect 11805 12801 11839 12835
rect 11839 12801 11848 12835
rect 11796 12792 11848 12801
rect 12440 12928 12492 12980
rect 12716 12928 12768 12980
rect 12348 12860 12400 12912
rect 13176 12860 13228 12912
rect 14464 12971 14516 12980
rect 14464 12937 14473 12971
rect 14473 12937 14507 12971
rect 14507 12937 14516 12971
rect 14464 12928 14516 12937
rect 7472 12656 7524 12708
rect 9404 12724 9456 12776
rect 11980 12724 12032 12776
rect 13912 12792 13964 12844
rect 14004 12835 14056 12844
rect 14004 12801 14013 12835
rect 14013 12801 14047 12835
rect 14047 12801 14056 12835
rect 14004 12792 14056 12801
rect 15108 12792 15160 12844
rect 14188 12724 14240 12776
rect 13544 12656 13596 12708
rect 13820 12656 13872 12708
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 7012 12588 7064 12640
rect 7656 12588 7708 12640
rect 7932 12588 7984 12640
rect 9956 12588 10008 12640
rect 10508 12631 10560 12640
rect 10508 12597 10517 12631
rect 10517 12597 10551 12631
rect 10551 12597 10560 12631
rect 10508 12588 10560 12597
rect 10600 12588 10652 12640
rect 2663 12486 2715 12538
rect 2727 12486 2779 12538
rect 2791 12486 2843 12538
rect 2855 12486 2907 12538
rect 2919 12486 2971 12538
rect 6090 12486 6142 12538
rect 6154 12486 6206 12538
rect 6218 12486 6270 12538
rect 6282 12486 6334 12538
rect 6346 12486 6398 12538
rect 9517 12486 9569 12538
rect 9581 12486 9633 12538
rect 9645 12486 9697 12538
rect 9709 12486 9761 12538
rect 9773 12486 9825 12538
rect 12944 12486 12996 12538
rect 13008 12486 13060 12538
rect 13072 12486 13124 12538
rect 13136 12486 13188 12538
rect 13200 12486 13252 12538
rect 1860 12384 1912 12436
rect 4988 12384 5040 12436
rect 9680 12384 9732 12436
rect 11612 12384 11664 12436
rect 7380 12316 7432 12368
rect 14096 12384 14148 12436
rect 15936 12384 15988 12436
rect 7564 12291 7616 12300
rect 7564 12257 7573 12291
rect 7573 12257 7607 12291
rect 7607 12257 7616 12291
rect 7564 12248 7616 12257
rect 7932 12291 7984 12300
rect 7932 12257 7966 12291
rect 7966 12257 7984 12291
rect 7932 12248 7984 12257
rect 10324 12248 10376 12300
rect 10876 12248 10928 12300
rect 2412 12180 2464 12232
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 6736 12180 6788 12232
rect 7012 12180 7064 12232
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 11612 12291 11664 12300
rect 11612 12257 11621 12291
rect 11621 12257 11655 12291
rect 11655 12257 11664 12291
rect 11612 12248 11664 12257
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 13360 12248 13412 12300
rect 13452 12248 13504 12300
rect 848 12044 900 12096
rect 7840 12044 7892 12096
rect 8392 12044 8444 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 9956 12044 10008 12096
rect 10416 12112 10468 12164
rect 10784 12112 10836 12164
rect 10692 12044 10744 12096
rect 10876 12087 10928 12096
rect 10876 12053 10885 12087
rect 10885 12053 10919 12087
rect 10919 12053 10928 12087
rect 10876 12044 10928 12053
rect 12622 12223 12674 12232
rect 12622 12189 12658 12223
rect 12658 12189 12674 12223
rect 12622 12180 12674 12189
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 14280 12223 14332 12232
rect 14280 12189 14289 12223
rect 14289 12189 14323 12223
rect 14323 12189 14332 12223
rect 14280 12180 14332 12189
rect 13820 12044 13872 12096
rect 4376 11942 4428 11994
rect 4440 11942 4492 11994
rect 4504 11942 4556 11994
rect 4568 11942 4620 11994
rect 4632 11942 4684 11994
rect 7803 11942 7855 11994
rect 7867 11942 7919 11994
rect 7931 11942 7983 11994
rect 7995 11942 8047 11994
rect 8059 11942 8111 11994
rect 11230 11942 11282 11994
rect 11294 11942 11346 11994
rect 11358 11942 11410 11994
rect 11422 11942 11474 11994
rect 11486 11942 11538 11994
rect 14657 11942 14709 11994
rect 14721 11942 14773 11994
rect 14785 11942 14837 11994
rect 14849 11942 14901 11994
rect 14913 11942 14965 11994
rect 5540 11840 5592 11892
rect 3792 11772 3844 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 6920 11704 6972 11756
rect 8208 11840 8260 11892
rect 8392 11840 8444 11892
rect 10140 11840 10192 11892
rect 10784 11840 10836 11892
rect 11152 11840 11204 11892
rect 11612 11840 11664 11892
rect 13360 11840 13412 11892
rect 15568 11840 15620 11892
rect 7288 11772 7340 11824
rect 8852 11747 8904 11756
rect 8852 11713 8861 11747
rect 8861 11713 8895 11747
rect 8895 11713 8904 11747
rect 8852 11704 8904 11713
rect 10876 11772 10928 11824
rect 9864 11704 9916 11756
rect 10692 11704 10744 11756
rect 12348 11704 12400 11756
rect 5632 11636 5684 11688
rect 9772 11636 9824 11688
rect 10876 11636 10928 11688
rect 11152 11636 11204 11688
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 6736 11568 6788 11620
rect 13544 11679 13596 11688
rect 13544 11645 13578 11679
rect 13578 11645 13596 11679
rect 13544 11636 13596 11645
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 848 11500 900 11552
rect 12716 11568 12768 11620
rect 13268 11568 13320 11620
rect 10600 11500 10652 11552
rect 12072 11500 12124 11552
rect 12900 11500 12952 11552
rect 13452 11500 13504 11552
rect 2663 11398 2715 11450
rect 2727 11398 2779 11450
rect 2791 11398 2843 11450
rect 2855 11398 2907 11450
rect 2919 11398 2971 11450
rect 6090 11398 6142 11450
rect 6154 11398 6206 11450
rect 6218 11398 6270 11450
rect 6282 11398 6334 11450
rect 6346 11398 6398 11450
rect 9517 11398 9569 11450
rect 9581 11398 9633 11450
rect 9645 11398 9697 11450
rect 9709 11398 9761 11450
rect 9773 11398 9825 11450
rect 12944 11398 12996 11450
rect 13008 11398 13060 11450
rect 13072 11398 13124 11450
rect 13136 11398 13188 11450
rect 13200 11398 13252 11450
rect 5724 11296 5776 11348
rect 7564 11296 7616 11348
rect 8852 11296 8904 11348
rect 9680 11296 9732 11348
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 6460 11160 6512 11212
rect 10692 11296 10744 11348
rect 11244 11296 11296 11348
rect 12256 11296 12308 11348
rect 12808 11296 12860 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 13544 11228 13596 11280
rect 3884 11092 3936 11144
rect 5816 11092 5868 11144
rect 10416 11092 10468 11144
rect 11244 11135 11296 11144
rect 11244 11101 11251 11135
rect 11251 11101 11285 11135
rect 11285 11101 11296 11135
rect 11244 11092 11296 11101
rect 12072 11092 12124 11144
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12676 11135
rect 12624 11092 12676 11101
rect 8576 11024 8628 11076
rect 13820 11160 13872 11212
rect 14096 11092 14148 11144
rect 15200 11092 15252 11144
rect 11704 10956 11756 11008
rect 12348 10956 12400 11008
rect 12716 10956 12768 11008
rect 13912 10956 13964 11008
rect 4376 10854 4428 10906
rect 4440 10854 4492 10906
rect 4504 10854 4556 10906
rect 4568 10854 4620 10906
rect 4632 10854 4684 10906
rect 7803 10854 7855 10906
rect 7867 10854 7919 10906
rect 7931 10854 7983 10906
rect 7995 10854 8047 10906
rect 8059 10854 8111 10906
rect 11230 10854 11282 10906
rect 11294 10854 11346 10906
rect 11358 10854 11410 10906
rect 11422 10854 11474 10906
rect 11486 10854 11538 10906
rect 14657 10854 14709 10906
rect 14721 10854 14773 10906
rect 14785 10854 14837 10906
rect 14849 10854 14901 10906
rect 14913 10854 14965 10906
rect 1492 10752 1544 10804
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 12624 10752 12676 10804
rect 13728 10752 13780 10804
rect 15844 10752 15896 10804
rect 4252 10684 4304 10736
rect 5356 10684 5408 10736
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6880 10659
rect 6828 10616 6880 10625
rect 6368 10548 6420 10600
rect 848 10412 900 10464
rect 5540 10480 5592 10532
rect 7840 10548 7892 10600
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 5448 10412 5500 10464
rect 9680 10548 9732 10600
rect 14188 10684 14240 10736
rect 12532 10616 12584 10668
rect 15108 10616 15160 10668
rect 11980 10548 12032 10600
rect 12256 10480 12308 10532
rect 6368 10412 6420 10464
rect 7380 10412 7432 10464
rect 8116 10412 8168 10464
rect 8484 10412 8536 10464
rect 11612 10412 11664 10464
rect 12072 10412 12124 10464
rect 2663 10310 2715 10362
rect 2727 10310 2779 10362
rect 2791 10310 2843 10362
rect 2855 10310 2907 10362
rect 2919 10310 2971 10362
rect 6090 10310 6142 10362
rect 6154 10310 6206 10362
rect 6218 10310 6270 10362
rect 6282 10310 6334 10362
rect 6346 10310 6398 10362
rect 9517 10310 9569 10362
rect 9581 10310 9633 10362
rect 9645 10310 9697 10362
rect 9709 10310 9761 10362
rect 9773 10310 9825 10362
rect 12944 10310 12996 10362
rect 13008 10310 13060 10362
rect 13072 10310 13124 10362
rect 13136 10310 13188 10362
rect 13200 10310 13252 10362
rect 1308 10004 1360 10056
rect 1584 10004 1636 10056
rect 8484 10208 8536 10260
rect 9404 10208 9456 10260
rect 5264 10140 5316 10192
rect 5448 10140 5500 10192
rect 7656 10140 7708 10192
rect 5080 10072 5132 10124
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 7472 10072 7524 10124
rect 7840 10115 7892 10124
rect 7840 10081 7849 10115
rect 7849 10081 7883 10115
rect 7883 10081 7892 10115
rect 7840 10072 7892 10081
rect 12072 10208 12124 10260
rect 13268 10208 13320 10260
rect 13360 10208 13412 10260
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 14096 10208 14148 10260
rect 10416 10140 10468 10192
rect 6552 10004 6604 10056
rect 5632 9936 5684 9988
rect 5908 9936 5960 9988
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 9220 10004 9272 10056
rect 10508 10004 10560 10056
rect 11060 10004 11112 10056
rect 12256 10004 12308 10056
rect 13820 10140 13872 10192
rect 14648 10072 14700 10124
rect 15200 10004 15252 10056
rect 1584 9868 1636 9920
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 5264 9868 5316 9920
rect 5356 9911 5408 9920
rect 5356 9877 5365 9911
rect 5365 9877 5399 9911
rect 5399 9877 5408 9911
rect 5356 9868 5408 9877
rect 7472 9868 7524 9920
rect 15108 9936 15160 9988
rect 13268 9868 13320 9920
rect 4376 9766 4428 9818
rect 4440 9766 4492 9818
rect 4504 9766 4556 9818
rect 4568 9766 4620 9818
rect 4632 9766 4684 9818
rect 7803 9766 7855 9818
rect 7867 9766 7919 9818
rect 7931 9766 7983 9818
rect 7995 9766 8047 9818
rect 8059 9766 8111 9818
rect 11230 9766 11282 9818
rect 11294 9766 11346 9818
rect 11358 9766 11410 9818
rect 11422 9766 11474 9818
rect 11486 9766 11538 9818
rect 14657 9766 14709 9818
rect 14721 9766 14773 9818
rect 14785 9766 14837 9818
rect 14849 9766 14901 9818
rect 14913 9766 14965 9818
rect 1492 9664 1544 9716
rect 940 9596 992 9648
rect 5080 9664 5132 9716
rect 5632 9664 5684 9716
rect 4160 9596 4212 9648
rect 2412 9528 2464 9580
rect 5356 9596 5408 9648
rect 7472 9664 7524 9716
rect 9956 9664 10008 9716
rect 10416 9664 10468 9716
rect 10692 9664 10744 9716
rect 11520 9664 11572 9716
rect 12440 9664 12492 9716
rect 13544 9664 13596 9716
rect 14096 9664 14148 9716
rect 15384 9664 15436 9716
rect 5264 9460 5316 9512
rect 6552 9392 6604 9444
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 3976 9324 4028 9376
rect 7380 9460 7432 9512
rect 7288 9324 7340 9376
rect 8300 9571 8352 9580
rect 8300 9537 8309 9571
rect 8309 9537 8343 9571
rect 8343 9537 8352 9571
rect 8300 9528 8352 9537
rect 9864 9528 9916 9580
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 11336 9571 11388 9580
rect 11336 9537 11345 9571
rect 11345 9537 11379 9571
rect 11379 9537 11388 9571
rect 11336 9528 11388 9537
rect 7656 9460 7708 9512
rect 8024 9503 8076 9512
rect 8024 9469 8033 9503
rect 8033 9469 8067 9503
rect 8067 9469 8076 9503
rect 8024 9460 8076 9469
rect 8208 9460 8260 9512
rect 9128 9460 9180 9512
rect 9404 9460 9456 9512
rect 10232 9460 10284 9512
rect 10508 9503 10560 9512
rect 10508 9469 10542 9503
rect 10542 9469 10560 9503
rect 10508 9460 10560 9469
rect 7840 9392 7892 9444
rect 10140 9435 10192 9444
rect 10140 9401 10149 9435
rect 10149 9401 10183 9435
rect 10183 9401 10192 9435
rect 10140 9392 10192 9401
rect 11152 9392 11204 9444
rect 11704 9392 11756 9444
rect 11980 9528 12032 9580
rect 12716 9596 12768 9648
rect 14372 9596 14424 9648
rect 12532 9528 12584 9580
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 12808 9460 12860 9512
rect 12072 9392 12124 9444
rect 10508 9324 10560 9376
rect 12440 9324 12492 9376
rect 13820 9324 13872 9376
rect 2663 9222 2715 9274
rect 2727 9222 2779 9274
rect 2791 9222 2843 9274
rect 2855 9222 2907 9274
rect 2919 9222 2971 9274
rect 6090 9222 6142 9274
rect 6154 9222 6206 9274
rect 6218 9222 6270 9274
rect 6282 9222 6334 9274
rect 6346 9222 6398 9274
rect 9517 9222 9569 9274
rect 9581 9222 9633 9274
rect 9645 9222 9697 9274
rect 9709 9222 9761 9274
rect 9773 9222 9825 9274
rect 12944 9222 12996 9274
rect 13008 9222 13060 9274
rect 13072 9222 13124 9274
rect 13136 9222 13188 9274
rect 13200 9222 13252 9274
rect 1492 9120 1544 9172
rect 10140 9120 10192 9172
rect 12072 9120 12124 9172
rect 15108 9120 15160 9172
rect 12992 9052 13044 9104
rect 7288 8984 7340 9036
rect 8392 8984 8444 9036
rect 9864 9027 9916 9036
rect 9864 8993 9873 9027
rect 9873 8993 9907 9027
rect 9907 8993 9916 9027
rect 9864 8984 9916 8993
rect 10324 8984 10376 9036
rect 10692 8984 10744 9036
rect 1400 8848 1452 8900
rect 7472 8916 7524 8968
rect 8024 8916 8076 8968
rect 8852 8916 8904 8968
rect 7840 8848 7892 8900
rect 9036 8848 9088 8900
rect 9956 8959 10008 8968
rect 9956 8925 9990 8959
rect 9990 8925 10008 8959
rect 10968 8984 11020 9036
rect 12440 8984 12492 9036
rect 9956 8916 10008 8925
rect 11244 8916 11296 8968
rect 11980 8916 12032 8968
rect 12072 8959 12124 8968
rect 12072 8925 12081 8959
rect 12081 8925 12115 8959
rect 12115 8925 12124 8959
rect 12072 8916 12124 8925
rect 14372 8984 14424 9036
rect 14464 8984 14516 9036
rect 10692 8848 10744 8900
rect 10876 8848 10928 8900
rect 12900 8848 12952 8900
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 9312 8780 9364 8832
rect 9956 8780 10008 8832
rect 10232 8780 10284 8832
rect 12532 8780 12584 8832
rect 13452 8780 13504 8832
rect 4376 8678 4428 8730
rect 4440 8678 4492 8730
rect 4504 8678 4556 8730
rect 4568 8678 4620 8730
rect 4632 8678 4684 8730
rect 7803 8678 7855 8730
rect 7867 8678 7919 8730
rect 7931 8678 7983 8730
rect 7995 8678 8047 8730
rect 8059 8678 8111 8730
rect 11230 8678 11282 8730
rect 11294 8678 11346 8730
rect 11358 8678 11410 8730
rect 11422 8678 11474 8730
rect 11486 8678 11538 8730
rect 14657 8678 14709 8730
rect 14721 8678 14773 8730
rect 14785 8678 14837 8730
rect 14849 8678 14901 8730
rect 14913 8678 14965 8730
rect 2136 8576 2188 8628
rect 2412 8576 2464 8628
rect 4988 8508 5040 8560
rect 6460 8576 6512 8628
rect 6552 8576 6604 8628
rect 9956 8576 10008 8628
rect 10232 8576 10284 8628
rect 10876 8576 10928 8628
rect 12716 8576 12768 8628
rect 13544 8576 13596 8628
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 7564 8440 7616 8492
rect 9496 8440 9548 8492
rect 9772 8440 9824 8492
rect 10416 8483 10468 8492
rect 10416 8449 10450 8483
rect 10450 8449 10468 8483
rect 10416 8440 10468 8449
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 11428 8440 11480 8492
rect 8576 8415 8628 8424
rect 8576 8381 8585 8415
rect 8585 8381 8619 8415
rect 8619 8381 8628 8415
rect 8576 8372 8628 8381
rect 7472 8304 7524 8356
rect 9680 8372 9732 8424
rect 11612 8372 11664 8424
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 12532 8483 12584 8492
rect 12532 8449 12566 8483
rect 12566 8449 12584 8483
rect 12532 8440 12584 8449
rect 13728 8440 13780 8492
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 10048 8347 10100 8356
rect 10048 8313 10063 8347
rect 10063 8313 10097 8347
rect 10097 8313 10100 8347
rect 10048 8304 10100 8313
rect 11428 8304 11480 8356
rect 2136 8279 2188 8288
rect 2136 8245 2145 8279
rect 2145 8245 2179 8279
rect 2179 8245 2188 8279
rect 2136 8236 2188 8245
rect 7932 8236 7984 8288
rect 10416 8236 10468 8288
rect 11152 8236 11204 8288
rect 11612 8236 11664 8288
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 13544 8372 13596 8424
rect 14096 8372 14148 8424
rect 12900 8236 12952 8288
rect 13360 8236 13412 8288
rect 2663 8134 2715 8186
rect 2727 8134 2779 8186
rect 2791 8134 2843 8186
rect 2855 8134 2907 8186
rect 2919 8134 2971 8186
rect 6090 8134 6142 8186
rect 6154 8134 6206 8186
rect 6218 8134 6270 8186
rect 6282 8134 6334 8186
rect 6346 8134 6398 8186
rect 9517 8134 9569 8186
rect 9581 8134 9633 8186
rect 9645 8134 9697 8186
rect 9709 8134 9761 8186
rect 9773 8134 9825 8186
rect 12944 8134 12996 8186
rect 13008 8134 13060 8186
rect 13072 8134 13124 8186
rect 13136 8134 13188 8186
rect 13200 8134 13252 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 6736 8032 6788 8084
rect 7196 8032 7248 8084
rect 7012 7896 7064 7948
rect 2136 7828 2188 7880
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 7472 7896 7524 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 8576 8032 8628 8084
rect 9128 8032 9180 8084
rect 7932 7939 7984 7948
rect 11796 8032 11848 8084
rect 9956 7964 10008 8016
rect 7932 7905 7966 7939
rect 7966 7905 7984 7939
rect 7932 7896 7984 7905
rect 9772 7896 9824 7948
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 11244 7964 11296 8016
rect 10600 7939 10652 7948
rect 10600 7905 10609 7939
rect 10609 7905 10643 7939
rect 10643 7905 10652 7939
rect 10600 7896 10652 7905
rect 11152 7896 11204 7948
rect 4804 7692 4856 7744
rect 6736 7692 6788 7744
rect 9128 7828 9180 7880
rect 9404 7871 9456 7880
rect 9404 7837 9413 7871
rect 9413 7837 9447 7871
rect 9447 7837 9456 7871
rect 9404 7828 9456 7837
rect 10416 7871 10468 7880
rect 10416 7837 10450 7871
rect 10450 7837 10468 7871
rect 10416 7828 10468 7837
rect 12716 8032 12768 8084
rect 12900 7964 12952 8016
rect 12716 7896 12768 7948
rect 12072 7828 12124 7880
rect 9036 7760 9088 7812
rect 14188 7828 14240 7880
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 14556 7760 14608 7812
rect 12624 7692 12676 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 4376 7590 4428 7642
rect 4440 7590 4492 7642
rect 4504 7590 4556 7642
rect 4568 7590 4620 7642
rect 4632 7590 4684 7642
rect 7803 7590 7855 7642
rect 7867 7590 7919 7642
rect 7931 7590 7983 7642
rect 7995 7590 8047 7642
rect 8059 7590 8111 7642
rect 11230 7590 11282 7642
rect 11294 7590 11346 7642
rect 11358 7590 11410 7642
rect 11422 7590 11474 7642
rect 11486 7590 11538 7642
rect 14657 7590 14709 7642
rect 14721 7590 14773 7642
rect 14785 7590 14837 7642
rect 14849 7590 14901 7642
rect 14913 7590 14965 7642
rect 6000 7488 6052 7540
rect 6828 7488 6880 7540
rect 7564 7531 7616 7540
rect 7564 7497 7573 7531
rect 7573 7497 7607 7531
rect 7607 7497 7616 7531
rect 7564 7488 7616 7497
rect 9588 7488 9640 7540
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 5724 7352 5776 7404
rect 7196 7420 7248 7472
rect 6828 7395 6880 7404
rect 6828 7361 6835 7395
rect 6835 7361 6869 7395
rect 6869 7361 6880 7395
rect 6828 7352 6880 7361
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 9036 7352 9088 7404
rect 11888 7488 11940 7540
rect 12348 7488 12400 7540
rect 13268 7488 13320 7540
rect 15660 7488 15712 7540
rect 9956 7420 10008 7472
rect 10600 7420 10652 7472
rect 10784 7352 10836 7404
rect 8208 7216 8260 7268
rect 848 7148 900 7200
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 11888 7284 11940 7336
rect 12256 7352 12308 7404
rect 12808 7395 12860 7404
rect 12808 7361 12817 7395
rect 12817 7361 12851 7395
rect 12851 7361 12860 7395
rect 12808 7352 12860 7361
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13728 7352 13780 7404
rect 12716 7284 12768 7336
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 10416 7148 10468 7200
rect 12532 7148 12584 7200
rect 14372 7148 14424 7200
rect 2663 7046 2715 7098
rect 2727 7046 2779 7098
rect 2791 7046 2843 7098
rect 2855 7046 2907 7098
rect 2919 7046 2971 7098
rect 6090 7046 6142 7098
rect 6154 7046 6206 7098
rect 6218 7046 6270 7098
rect 6282 7046 6334 7098
rect 6346 7046 6398 7098
rect 9517 7046 9569 7098
rect 9581 7046 9633 7098
rect 9645 7046 9697 7098
rect 9709 7046 9761 7098
rect 9773 7046 9825 7098
rect 12944 7046 12996 7098
rect 13008 7046 13060 7098
rect 13072 7046 13124 7098
rect 13136 7046 13188 7098
rect 13200 7046 13252 7098
rect 2136 6944 2188 6996
rect 6828 6944 6880 6996
rect 9956 6944 10008 6996
rect 8116 6876 8168 6928
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 6920 6740 6972 6792
rect 9404 6808 9456 6860
rect 10048 6876 10100 6928
rect 10876 6944 10928 6996
rect 14372 6987 14424 6996
rect 14372 6953 14381 6987
rect 14381 6953 14415 6987
rect 14415 6953 14424 6987
rect 14372 6944 14424 6953
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 9864 6740 9916 6792
rect 9680 6672 9732 6724
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11612 6808 11664 6860
rect 12256 6808 12308 6860
rect 13360 6808 13412 6860
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11796 6740 11848 6792
rect 12808 6783 12860 6792
rect 12808 6749 12817 6783
rect 12817 6749 12851 6783
rect 12851 6749 12860 6783
rect 12808 6740 12860 6749
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 14004 6740 14056 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 9956 6604 10008 6656
rect 12072 6604 12124 6656
rect 12532 6715 12584 6724
rect 12532 6681 12541 6715
rect 12541 6681 12575 6715
rect 12575 6681 12584 6715
rect 12532 6672 12584 6681
rect 12716 6672 12768 6724
rect 13912 6604 13964 6656
rect 4376 6502 4428 6554
rect 4440 6502 4492 6554
rect 4504 6502 4556 6554
rect 4568 6502 4620 6554
rect 4632 6502 4684 6554
rect 7803 6502 7855 6554
rect 7867 6502 7919 6554
rect 7931 6502 7983 6554
rect 7995 6502 8047 6554
rect 8059 6502 8111 6554
rect 11230 6502 11282 6554
rect 11294 6502 11346 6554
rect 11358 6502 11410 6554
rect 11422 6502 11474 6554
rect 11486 6502 11538 6554
rect 14657 6502 14709 6554
rect 14721 6502 14773 6554
rect 14785 6502 14837 6554
rect 14849 6502 14901 6554
rect 14913 6502 14965 6554
rect 848 6400 900 6452
rect 8300 6332 8352 6384
rect 11980 6400 12032 6452
rect 10692 6332 10744 6384
rect 12164 6332 12216 6384
rect 13176 6400 13228 6452
rect 13268 6332 13320 6384
rect 14464 6400 14516 6452
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 6920 6264 6972 6316
rect 7196 6196 7248 6248
rect 8852 6264 8904 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 10968 6264 11020 6316
rect 12808 6264 12860 6316
rect 12992 6264 13044 6316
rect 9312 6196 9364 6248
rect 12348 6196 12400 6248
rect 9404 6171 9456 6180
rect 9404 6137 9413 6171
rect 9413 6137 9447 6171
rect 9447 6137 9456 6171
rect 9404 6128 9456 6137
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 10324 6060 10376 6112
rect 10968 6128 11020 6180
rect 13912 6264 13964 6316
rect 15108 6264 15160 6316
rect 11152 6060 11204 6112
rect 2663 5958 2715 6010
rect 2727 5958 2779 6010
rect 2791 5958 2843 6010
rect 2855 5958 2907 6010
rect 2919 5958 2971 6010
rect 6090 5958 6142 6010
rect 6154 5958 6206 6010
rect 6218 5958 6270 6010
rect 6282 5958 6334 6010
rect 6346 5958 6398 6010
rect 9517 5958 9569 6010
rect 9581 5958 9633 6010
rect 9645 5958 9697 6010
rect 9709 5958 9761 6010
rect 9773 5958 9825 6010
rect 12944 5958 12996 6010
rect 13008 5958 13060 6010
rect 13072 5958 13124 6010
rect 13136 5958 13188 6010
rect 13200 5958 13252 6010
rect 2504 5856 2556 5908
rect 9128 5856 9180 5908
rect 11152 5856 11204 5908
rect 7196 5720 7248 5772
rect 9772 5763 9824 5772
rect 9772 5729 9781 5763
rect 9781 5729 9815 5763
rect 9815 5729 9824 5763
rect 9772 5720 9824 5729
rect 9956 5763 10008 5772
rect 9956 5729 9965 5763
rect 9965 5729 9999 5763
rect 9999 5729 10008 5763
rect 9956 5720 10008 5729
rect 10140 5720 10192 5772
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 10968 5763 11020 5772
rect 10968 5729 10977 5763
rect 10977 5729 11011 5763
rect 11011 5729 11020 5763
rect 10968 5720 11020 5729
rect 13544 5899 13596 5908
rect 13544 5865 13553 5899
rect 13553 5865 13587 5899
rect 13587 5865 13596 5899
rect 13544 5856 13596 5865
rect 14372 5899 14424 5908
rect 14372 5865 14381 5899
rect 14381 5865 14415 5899
rect 14415 5865 14424 5899
rect 14372 5856 14424 5865
rect 15292 5856 15344 5908
rect 12072 5788 12124 5840
rect 12256 5788 12308 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 6736 5652 6788 5704
rect 8208 5652 8260 5704
rect 9312 5652 9364 5704
rect 10876 5652 10928 5704
rect 11980 5720 12032 5772
rect 12716 5763 12768 5772
rect 12716 5729 12750 5763
rect 12750 5729 12768 5763
rect 12716 5720 12768 5729
rect 12900 5695 12952 5704
rect 12900 5661 12909 5695
rect 12909 5661 12943 5695
rect 12943 5661 12952 5695
rect 12900 5652 12952 5661
rect 14832 5652 14884 5704
rect 1584 5516 1636 5568
rect 5816 5516 5868 5568
rect 8300 5516 8352 5568
rect 11796 5584 11848 5636
rect 14280 5627 14332 5636
rect 14280 5593 14289 5627
rect 14289 5593 14323 5627
rect 14323 5593 14332 5627
rect 14280 5584 14332 5593
rect 11704 5516 11756 5568
rect 4376 5414 4428 5466
rect 4440 5414 4492 5466
rect 4504 5414 4556 5466
rect 4568 5414 4620 5466
rect 4632 5414 4684 5466
rect 7803 5414 7855 5466
rect 7867 5414 7919 5466
rect 7931 5414 7983 5466
rect 7995 5414 8047 5466
rect 8059 5414 8111 5466
rect 11230 5414 11282 5466
rect 11294 5414 11346 5466
rect 11358 5414 11410 5466
rect 11422 5414 11474 5466
rect 11486 5414 11538 5466
rect 14657 5414 14709 5466
rect 14721 5414 14773 5466
rect 14785 5414 14837 5466
rect 14849 5414 14901 5466
rect 14913 5414 14965 5466
rect 7656 5312 7708 5364
rect 8300 5249 8352 5296
rect 3976 5176 4028 5228
rect 7196 5176 7248 5228
rect 8300 5244 8325 5249
rect 8325 5244 8352 5249
rect 10140 5312 10192 5364
rect 13360 5312 13412 5364
rect 940 4972 992 5024
rect 8944 5176 8996 5228
rect 15108 5244 15160 5296
rect 8300 4972 8352 5024
rect 10784 5108 10836 5160
rect 13728 5176 13780 5228
rect 14004 5176 14056 5228
rect 12072 5040 12124 5092
rect 12532 4972 12584 5024
rect 2663 4870 2715 4922
rect 2727 4870 2779 4922
rect 2791 4870 2843 4922
rect 2855 4870 2907 4922
rect 2919 4870 2971 4922
rect 6090 4870 6142 4922
rect 6154 4870 6206 4922
rect 6218 4870 6270 4922
rect 6282 4870 6334 4922
rect 6346 4870 6398 4922
rect 9517 4870 9569 4922
rect 9581 4870 9633 4922
rect 9645 4870 9697 4922
rect 9709 4870 9761 4922
rect 9773 4870 9825 4922
rect 12944 4870 12996 4922
rect 13008 4870 13060 4922
rect 13072 4870 13124 4922
rect 13136 4870 13188 4922
rect 13200 4870 13252 4922
rect 848 4768 900 4820
rect 8300 4632 8352 4684
rect 11980 4768 12032 4820
rect 12072 4768 12124 4820
rect 12716 4768 12768 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 13912 4768 13964 4820
rect 11152 4632 11204 4684
rect 2044 4564 2096 4616
rect 7288 4496 7340 4548
rect 11060 4564 11112 4616
rect 12624 4496 12676 4548
rect 15200 4564 15252 4616
rect 4376 4326 4428 4378
rect 4440 4326 4492 4378
rect 4504 4326 4556 4378
rect 4568 4326 4620 4378
rect 4632 4326 4684 4378
rect 7803 4326 7855 4378
rect 7867 4326 7919 4378
rect 7931 4326 7983 4378
rect 7995 4326 8047 4378
rect 8059 4326 8111 4378
rect 11230 4326 11282 4378
rect 11294 4326 11346 4378
rect 11358 4326 11410 4378
rect 11422 4326 11474 4378
rect 11486 4326 11538 4378
rect 14657 4326 14709 4378
rect 14721 4326 14773 4378
rect 14785 4326 14837 4378
rect 14849 4326 14901 4378
rect 14913 4326 14965 4378
rect 12624 4224 12676 4276
rect 10600 4156 10652 4208
rect 756 4088 808 4140
rect 8760 4131 8812 4140
rect 8760 4097 8767 4131
rect 8767 4097 8801 4131
rect 8801 4097 8812 4131
rect 8760 4088 8812 4097
rect 11152 4088 11204 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11940 4131
rect 11888 4088 11940 4097
rect 8300 4020 8352 4072
rect 9404 3952 9456 4004
rect 3424 3884 3476 3936
rect 12532 4020 12584 4072
rect 12072 3884 12124 3936
rect 12348 3884 12400 3936
rect 13820 3884 13872 3936
rect 2663 3782 2715 3834
rect 2727 3782 2779 3834
rect 2791 3782 2843 3834
rect 2855 3782 2907 3834
rect 2919 3782 2971 3834
rect 6090 3782 6142 3834
rect 6154 3782 6206 3834
rect 6218 3782 6270 3834
rect 6282 3782 6334 3834
rect 6346 3782 6398 3834
rect 9517 3782 9569 3834
rect 9581 3782 9633 3834
rect 9645 3782 9697 3834
rect 9709 3782 9761 3834
rect 9773 3782 9825 3834
rect 12944 3782 12996 3834
rect 13008 3782 13060 3834
rect 13072 3782 13124 3834
rect 13136 3782 13188 3834
rect 13200 3782 13252 3834
rect 13268 3680 13320 3732
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 12072 3587 12124 3596
rect 12072 3553 12081 3587
rect 12081 3553 12115 3587
rect 12115 3553 12124 3587
rect 12072 3544 12124 3553
rect 11152 3476 11204 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 4376 3238 4428 3290
rect 4440 3238 4492 3290
rect 4504 3238 4556 3290
rect 4568 3238 4620 3290
rect 4632 3238 4684 3290
rect 7803 3238 7855 3290
rect 7867 3238 7919 3290
rect 7931 3238 7983 3290
rect 7995 3238 8047 3290
rect 8059 3238 8111 3290
rect 11230 3238 11282 3290
rect 11294 3238 11346 3290
rect 11358 3238 11410 3290
rect 11422 3238 11474 3290
rect 11486 3238 11538 3290
rect 14657 3238 14709 3290
rect 14721 3238 14773 3290
rect 14785 3238 14837 3290
rect 14849 3238 14901 3290
rect 14913 3238 14965 3290
rect 2663 2694 2715 2746
rect 2727 2694 2779 2746
rect 2791 2694 2843 2746
rect 2855 2694 2907 2746
rect 2919 2694 2971 2746
rect 6090 2694 6142 2746
rect 6154 2694 6206 2746
rect 6218 2694 6270 2746
rect 6282 2694 6334 2746
rect 6346 2694 6398 2746
rect 9517 2694 9569 2746
rect 9581 2694 9633 2746
rect 9645 2694 9697 2746
rect 9709 2694 9761 2746
rect 9773 2694 9825 2746
rect 12944 2694 12996 2746
rect 13008 2694 13060 2746
rect 13072 2694 13124 2746
rect 13136 2694 13188 2746
rect 13200 2694 13252 2746
rect 1216 2592 1268 2644
rect 4068 2320 4120 2372
rect 4376 2150 4428 2202
rect 4440 2150 4492 2202
rect 4504 2150 4556 2202
rect 4568 2150 4620 2202
rect 4632 2150 4684 2202
rect 7803 2150 7855 2202
rect 7867 2150 7919 2202
rect 7931 2150 7983 2202
rect 7995 2150 8047 2202
rect 8059 2150 8111 2202
rect 11230 2150 11282 2202
rect 11294 2150 11346 2202
rect 11358 2150 11410 2202
rect 11422 2150 11474 2202
rect 11486 2150 11538 2202
rect 14657 2150 14709 2202
rect 14721 2150 14773 2202
rect 14785 2150 14837 2202
rect 14849 2150 14901 2202
rect 14913 2150 14965 2202
rect 4068 2091 4120 2100
rect 4068 2057 4077 2091
rect 4077 2057 4111 2091
rect 4111 2057 4120 2091
rect 4068 2048 4120 2057
rect 2228 1980 2280 2032
rect 5816 2091 5868 2100
rect 5816 2057 5825 2091
rect 5825 2057 5859 2091
rect 5859 2057 5868 2091
rect 5816 2048 5868 2057
rect 6644 2048 6696 2100
rect 7196 2091 7248 2100
rect 7196 2057 7205 2091
rect 7205 2057 7239 2091
rect 7239 2057 7248 2091
rect 7196 2048 7248 2057
rect 7656 2048 7708 2100
rect 8668 2091 8720 2100
rect 8668 2057 8677 2091
rect 8677 2057 8711 2091
rect 8711 2057 8720 2091
rect 8668 2048 8720 2057
rect 10876 2091 10928 2100
rect 10876 2057 10885 2091
rect 10885 2057 10919 2091
rect 10919 2057 10928 2091
rect 10876 2048 10928 2057
rect 12440 2048 12492 2100
rect 13360 2048 13412 2100
rect 15752 2048 15804 2100
rect 2136 1955 2188 1964
rect 2136 1921 2145 1955
rect 2145 1921 2179 1955
rect 2179 1921 2188 1955
rect 2136 1912 2188 1921
rect 4252 1955 4304 1964
rect 4252 1921 4261 1955
rect 4261 1921 4295 1955
rect 4295 1921 4304 1955
rect 4252 1912 4304 1921
rect 4988 1955 5040 1964
rect 4988 1921 4997 1955
rect 4997 1921 5031 1955
rect 5031 1921 5040 1955
rect 4988 1912 5040 1921
rect 5724 1955 5776 1964
rect 5724 1921 5733 1955
rect 5733 1921 5767 1955
rect 5767 1921 5776 1955
rect 5724 1912 5776 1921
rect 6460 1955 6512 1964
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 12072 1980 12124 2032
rect 13452 1980 13504 2032
rect 15016 1980 15068 2032
rect 7104 1955 7156 1964
rect 7104 1921 7113 1955
rect 7113 1921 7147 1955
rect 7147 1921 7156 1955
rect 7104 1912 7156 1921
rect 7840 1955 7892 1964
rect 7840 1921 7849 1955
rect 7849 1921 7883 1955
rect 7883 1921 7892 1955
rect 7840 1912 7892 1921
rect 8576 1955 8628 1964
rect 8576 1921 8585 1955
rect 8585 1921 8619 1955
rect 8619 1921 8628 1955
rect 8576 1912 8628 1921
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 10048 1955 10100 1964
rect 10048 1921 10057 1955
rect 10057 1921 10091 1955
rect 10091 1921 10100 1955
rect 10048 1912 10100 1921
rect 10784 1955 10836 1964
rect 10784 1921 10793 1955
rect 10793 1921 10827 1955
rect 10827 1921 10836 1955
rect 10784 1912 10836 1921
rect 11612 1955 11664 1964
rect 11612 1921 11621 1955
rect 11621 1921 11655 1955
rect 11655 1921 11664 1955
rect 11612 1912 11664 1921
rect 12256 1955 12308 1964
rect 12256 1921 12265 1955
rect 12265 1921 12299 1955
rect 12299 1921 12308 1955
rect 12256 1912 12308 1921
rect 13268 1912 13320 1964
rect 13728 1955 13780 1964
rect 13728 1921 13737 1955
rect 13737 1921 13771 1955
rect 13771 1921 13780 1955
rect 13728 1912 13780 1921
rect 3240 1776 3292 1828
rect 2412 1708 2464 1760
rect 11704 1751 11756 1760
rect 11704 1717 11713 1751
rect 11713 1717 11747 1751
rect 11747 1717 11756 1751
rect 11704 1708 11756 1717
rect 2663 1606 2715 1658
rect 2727 1606 2779 1658
rect 2791 1606 2843 1658
rect 2855 1606 2907 1658
rect 2919 1606 2971 1658
rect 6090 1606 6142 1658
rect 6154 1606 6206 1658
rect 6218 1606 6270 1658
rect 6282 1606 6334 1658
rect 6346 1606 6398 1658
rect 9517 1606 9569 1658
rect 9581 1606 9633 1658
rect 9645 1606 9697 1658
rect 9709 1606 9761 1658
rect 9773 1606 9825 1658
rect 12944 1606 12996 1658
rect 13008 1606 13060 1658
rect 13072 1606 13124 1658
rect 13136 1606 13188 1658
rect 13200 1606 13252 1658
rect 4252 1504 4304 1556
rect 4988 1504 5040 1556
rect 5724 1504 5776 1556
rect 6460 1504 6512 1556
rect 7104 1504 7156 1556
rect 7840 1504 7892 1556
rect 8576 1504 8628 1556
rect 9312 1504 9364 1556
rect 10048 1504 10100 1556
rect 10784 1504 10836 1556
rect 11612 1504 11664 1556
rect 12256 1504 12308 1556
rect 13268 1504 13320 1556
rect 13452 1547 13504 1556
rect 13452 1513 13461 1547
rect 13461 1513 13495 1547
rect 13495 1513 13504 1547
rect 13452 1504 13504 1513
rect 13728 1547 13780 1556
rect 13728 1513 13737 1547
rect 13737 1513 13771 1547
rect 13771 1513 13780 1547
rect 13728 1504 13780 1513
rect 1308 1300 1360 1352
rect 1584 1300 1636 1352
rect 2228 1275 2280 1284
rect 2228 1241 2237 1275
rect 2237 1241 2271 1275
rect 2271 1241 2280 1275
rect 2228 1232 2280 1241
rect 2780 1300 2832 1352
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4252 1300 4304 1352
rect 4988 1300 5040 1352
rect 5724 1300 5776 1352
rect 6460 1300 6512 1352
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8668 1300 8720 1352
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 10416 1343 10468 1352
rect 10416 1309 10425 1343
rect 10425 1309 10459 1343
rect 10459 1309 10468 1343
rect 10416 1300 10468 1309
rect 10876 1300 10928 1352
rect 11612 1300 11664 1352
rect 12348 1300 12400 1352
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 13360 1343 13412 1352
rect 13360 1309 13369 1343
rect 13369 1309 13403 1343
rect 13403 1309 13412 1343
rect 13360 1300 13412 1309
rect 13912 1343 13964 1352
rect 13912 1309 13921 1343
rect 13921 1309 13955 1343
rect 13955 1309 13964 1343
rect 13912 1300 13964 1309
rect 14556 1300 14608 1352
rect 15476 1300 15528 1352
rect 12532 1232 12584 1284
rect 4376 1062 4428 1114
rect 4440 1062 4492 1114
rect 4504 1062 4556 1114
rect 4568 1062 4620 1114
rect 4632 1062 4684 1114
rect 7803 1062 7855 1114
rect 7867 1062 7919 1114
rect 7931 1062 7983 1114
rect 7995 1062 8047 1114
rect 8059 1062 8111 1114
rect 11230 1062 11282 1114
rect 11294 1062 11346 1114
rect 11358 1062 11410 1114
rect 11422 1062 11474 1114
rect 11486 1062 11538 1114
rect 14657 1062 14709 1114
rect 14721 1062 14773 1114
rect 14785 1062 14837 1114
rect 14849 1062 14901 1114
rect 14913 1062 14965 1114
rect 2228 960 2280 1012
rect 8392 960 8444 1012
rect 13084 960 13136 1012
rect 15292 960 15344 1012
<< metal2 >>
rect 570 44463 626 44623
rect 1306 44463 1362 44623
rect 2042 44463 2098 44623
rect 2778 44463 2834 44623
rect 3514 44463 3570 44623
rect 4250 44463 4306 44623
rect 4986 44463 5042 44623
rect 5722 44463 5778 44623
rect 6458 44463 6514 44623
rect 7194 44463 7250 44623
rect 7930 44463 7986 44623
rect 8036 44526 8248 44554
rect 584 43450 612 44463
rect 572 43444 624 43450
rect 572 43386 624 43392
rect 1320 43058 1348 44463
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1400 43104 1452 43110
rect 1320 43052 1400 43058
rect 1320 43046 1452 43052
rect 1320 43030 1440 43046
rect 1216 42628 1268 42634
rect 1216 42570 1268 42576
rect 756 41132 808 41138
rect 756 41074 808 41080
rect 768 40633 796 41074
rect 754 40624 810 40633
rect 754 40559 810 40568
rect 756 39432 808 39438
rect 756 39374 808 39380
rect 768 39001 796 39374
rect 754 38992 810 39001
rect 754 38927 810 38936
rect 756 38344 808 38350
rect 756 38286 808 38292
rect 768 38185 796 38286
rect 754 38176 810 38185
rect 754 38111 810 38120
rect 756 37868 808 37874
rect 756 37810 808 37816
rect 768 37369 796 37810
rect 754 37360 810 37369
rect 754 37295 810 37304
rect 756 36780 808 36786
rect 756 36722 808 36728
rect 768 36553 796 36722
rect 754 36544 810 36553
rect 754 36479 810 36488
rect 756 35080 808 35086
rect 756 35022 808 35028
rect 768 34921 796 35022
rect 754 34912 810 34921
rect 754 34847 810 34856
rect 756 33516 808 33522
rect 756 33458 808 33464
rect 768 33289 796 33458
rect 754 33280 810 33289
rect 754 33215 810 33224
rect 756 32904 808 32910
rect 756 32846 808 32852
rect 768 32473 796 32846
rect 754 32464 810 32473
rect 754 32399 810 32408
rect 756 31340 808 31346
rect 756 31282 808 31288
rect 768 30841 796 31282
rect 754 30832 810 30841
rect 754 30767 810 30776
rect 756 30252 808 30258
rect 756 30194 808 30200
rect 768 30025 796 30194
rect 754 30016 810 30025
rect 754 29951 810 29960
rect 756 29640 808 29646
rect 756 29582 808 29588
rect 768 29209 796 29582
rect 754 29200 810 29209
rect 754 29135 810 29144
rect 756 28552 808 28558
rect 756 28494 808 28500
rect 768 28393 796 28494
rect 754 28384 810 28393
rect 754 28319 810 28328
rect 756 26988 808 26994
rect 756 26930 808 26936
rect 768 26761 796 26930
rect 754 26752 810 26761
rect 754 26687 810 26696
rect 756 25288 808 25294
rect 756 25230 808 25236
rect 768 25129 796 25230
rect 754 25120 810 25129
rect 754 25055 810 25064
rect 756 24812 808 24818
rect 756 24754 808 24760
rect 768 24313 796 24754
rect 754 24304 810 24313
rect 754 24239 810 24248
rect 756 23656 808 23662
rect 756 23598 808 23604
rect 768 23497 796 23598
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 756 23044 808 23050
rect 756 22986 808 22992
rect 768 22681 796 22986
rect 754 22672 810 22681
rect 754 22607 810 22616
rect 756 21956 808 21962
rect 756 21898 808 21904
rect 768 21865 796 21898
rect 754 21856 810 21865
rect 754 21791 810 21800
rect 754 21040 810 21049
rect 754 20975 810 20984
rect 768 20942 796 20975
rect 756 20936 808 20942
rect 756 20878 808 20884
rect 756 20460 808 20466
rect 756 20402 808 20408
rect 768 20233 796 20402
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 756 19780 808 19786
rect 756 19722 808 19728
rect 768 19417 796 19722
rect 754 19408 810 19417
rect 754 19343 810 19352
rect 756 18760 808 18766
rect 756 18702 808 18708
rect 768 18601 796 18702
rect 754 18592 810 18601
rect 754 18527 810 18536
rect 572 18216 624 18222
rect 572 18158 624 18164
rect 584 160 612 18158
rect 756 17196 808 17202
rect 756 17138 808 17144
rect 768 16969 796 17138
rect 754 16960 810 16969
rect 754 16895 810 16904
rect 756 16516 808 16522
rect 756 16458 808 16464
rect 768 16153 796 16458
rect 754 16144 810 16153
rect 754 16079 810 16088
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15337 888 16050
rect 846 15328 902 15337
rect 846 15263 902 15272
rect 848 14612 900 14618
rect 848 14554 900 14560
rect 860 14521 888 14554
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 848 12096 900 12102
rect 846 12064 848 12073
rect 900 12064 902 12073
rect 846 11999 902 12008
rect 848 11552 900 11558
rect 848 11494 900 11500
rect 860 11257 888 11494
rect 846 11248 902 11257
rect 846 11183 902 11192
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 900 10432 902 10441
rect 846 10367 902 10376
rect 940 9648 992 9654
rect 938 9616 940 9625
rect 992 9616 994 9625
rect 938 9551 994 9560
rect 848 7200 900 7206
rect 846 7168 848 7177
rect 900 7168 902 7177
rect 846 7103 902 7112
rect 848 6452 900 6458
rect 848 6394 900 6400
rect 860 6361 888 6394
rect 846 6352 902 6361
rect 846 6287 902 6296
rect 846 5536 902 5545
rect 846 5471 902 5480
rect 860 4826 888 5471
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 848 4820 900 4826
rect 848 4762 900 4768
rect 952 4729 980 4966
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 756 4140 808 4146
rect 756 4082 808 4088
rect 768 3913 796 4082
rect 754 3904 810 3913
rect 754 3839 810 3848
rect 1228 2650 1256 42570
rect 1400 40044 1452 40050
rect 1400 39986 1452 39992
rect 1412 39953 1440 39986
rect 1398 39944 1454 39953
rect 1398 39879 1454 39888
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 35873 1440 36110
rect 1398 35864 1454 35873
rect 1398 35799 1454 35808
rect 1780 35290 1808 43250
rect 2056 43178 2084 44463
rect 2792 43450 2820 44463
rect 3528 43450 3556 44463
rect 4264 43450 4292 44463
rect 4376 43548 4684 43557
rect 4376 43546 4382 43548
rect 4438 43546 4462 43548
rect 4518 43546 4542 43548
rect 4598 43546 4622 43548
rect 4678 43546 4684 43548
rect 4438 43494 4440 43546
rect 4620 43494 4622 43546
rect 4376 43492 4382 43494
rect 4438 43492 4462 43494
rect 4518 43492 4542 43494
rect 4598 43492 4622 43494
rect 4678 43492 4684 43494
rect 4376 43483 4684 43492
rect 5000 43450 5028 44463
rect 5736 43450 5764 44463
rect 6472 43450 6500 44463
rect 7208 43450 7236 44463
rect 7944 44418 7972 44463
rect 8036 44418 8064 44526
rect 7944 44390 8064 44418
rect 7803 43548 8111 43557
rect 7803 43546 7809 43548
rect 7865 43546 7889 43548
rect 7945 43546 7969 43548
rect 8025 43546 8049 43548
rect 8105 43546 8111 43548
rect 7865 43494 7867 43546
rect 8047 43494 8049 43546
rect 7803 43492 7809 43494
rect 7865 43492 7889 43494
rect 7945 43492 7969 43494
rect 8025 43492 8049 43494
rect 8105 43492 8111 43494
rect 7803 43483 8111 43492
rect 8220 43450 8248 44526
rect 8666 44463 8722 44623
rect 9402 44463 9458 44623
rect 10138 44463 10194 44623
rect 10874 44463 10930 44623
rect 11610 44463 11666 44623
rect 12346 44463 12402 44623
rect 13082 44463 13138 44623
rect 13818 44463 13874 44623
rect 14554 44463 14610 44623
rect 15290 44463 15346 44623
rect 8680 43450 8708 44463
rect 9416 43450 9444 44463
rect 10152 43450 10180 44463
rect 10888 43450 10916 44463
rect 11230 43548 11538 43557
rect 11230 43546 11236 43548
rect 11292 43546 11316 43548
rect 11372 43546 11396 43548
rect 11452 43546 11476 43548
rect 11532 43546 11538 43548
rect 11292 43494 11294 43546
rect 11474 43494 11476 43546
rect 11230 43492 11236 43494
rect 11292 43492 11316 43494
rect 11372 43492 11396 43494
rect 11452 43492 11476 43494
rect 11532 43492 11538 43494
rect 11230 43483 11538 43492
rect 11624 43466 11652 44463
rect 2780 43444 2832 43450
rect 2780 43386 2832 43392
rect 3516 43444 3568 43450
rect 3516 43386 3568 43392
rect 4252 43444 4304 43450
rect 4252 43386 4304 43392
rect 4988 43444 5040 43450
rect 4988 43386 5040 43392
rect 5724 43444 5776 43450
rect 5724 43386 5776 43392
rect 6460 43444 6512 43450
rect 6460 43386 6512 43392
rect 7196 43444 7248 43450
rect 7196 43386 7248 43392
rect 8208 43444 8260 43450
rect 8208 43386 8260 43392
rect 8668 43444 8720 43450
rect 8668 43386 8720 43392
rect 9404 43444 9456 43450
rect 9404 43386 9456 43392
rect 10140 43444 10192 43450
rect 10140 43386 10192 43392
rect 10876 43444 10928 43450
rect 11624 43438 11744 43466
rect 12360 43450 12388 44463
rect 13096 43450 13124 44463
rect 13832 43450 13860 44463
rect 10876 43386 10928 43392
rect 2136 43308 2188 43314
rect 2136 43250 2188 43256
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 3792 43308 3844 43314
rect 3792 43250 3844 43256
rect 4344 43308 4396 43314
rect 4344 43250 4396 43256
rect 5080 43308 5132 43314
rect 5080 43250 5132 43256
rect 5816 43308 5868 43314
rect 5816 43250 5868 43256
rect 6552 43308 6604 43314
rect 6552 43250 6604 43256
rect 7288 43308 7340 43314
rect 7288 43250 7340 43256
rect 8024 43308 8076 43314
rect 8024 43250 8076 43256
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 9312 43308 9364 43314
rect 9312 43250 9364 43256
rect 10232 43308 10284 43314
rect 10232 43250 10284 43256
rect 11612 43308 11664 43314
rect 11612 43250 11664 43256
rect 2044 43172 2096 43178
rect 2044 43114 2096 43120
rect 2148 42906 2176 43250
rect 2136 42900 2188 42906
rect 2136 42842 2188 42848
rect 2228 42696 2280 42702
rect 2228 42638 2280 42644
rect 2240 42362 2268 42638
rect 2228 42356 2280 42362
rect 2228 42298 2280 42304
rect 2412 42288 2464 42294
rect 2412 42230 2464 42236
rect 2228 42220 2280 42226
rect 2228 42162 2280 42168
rect 2136 38344 2188 38350
rect 2136 38286 2188 38292
rect 2148 35894 2176 38286
rect 2240 36922 2268 42162
rect 2424 39012 2452 42230
rect 2332 38984 2452 39012
rect 2228 36916 2280 36922
rect 2228 36858 2280 36864
rect 2148 35866 2268 35894
rect 1768 35284 1820 35290
rect 1768 35226 1820 35232
rect 1952 35080 2004 35086
rect 1952 35022 2004 35028
rect 1964 34746 1992 35022
rect 1952 34740 2004 34746
rect 1952 34682 2004 34688
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 1412 34513 1440 34546
rect 1398 34504 1454 34513
rect 1398 34439 1454 34448
rect 1964 34202 1992 34546
rect 1952 34196 2004 34202
rect 1952 34138 2004 34144
rect 1676 32768 1728 32774
rect 1676 32710 1728 32716
rect 1688 32570 1716 32710
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31657 1440 31758
rect 1398 31648 1454 31657
rect 1398 31583 1454 31592
rect 1584 31136 1636 31142
rect 1584 31078 1636 31084
rect 1596 30938 1624 31078
rect 1584 30932 1636 30938
rect 1584 30874 1636 30880
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1596 28218 1624 28358
rect 1584 28212 1636 28218
rect 1584 28154 1636 28160
rect 1688 28098 1716 32506
rect 1768 32020 1820 32026
rect 1768 31962 1820 31968
rect 1492 28076 1544 28082
rect 1492 28018 1544 28024
rect 1596 28070 1716 28098
rect 1504 27577 1532 28018
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 1492 26308 1544 26314
rect 1492 26250 1544 26256
rect 1504 26217 1532 26250
rect 1596 26234 1624 28070
rect 1676 27872 1728 27878
rect 1676 27814 1728 27820
rect 1688 27713 1716 27814
rect 1674 27704 1730 27713
rect 1674 27639 1730 27648
rect 1490 26208 1546 26217
rect 1596 26206 1716 26234
rect 1490 26143 1546 26152
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1596 22778 1624 22918
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 1582 21448 1638 21457
rect 1582 21383 1638 21392
rect 1596 18970 1624 21383
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17921 1532 18226
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 1688 16574 1716 26206
rect 1412 16546 1716 16574
rect 1308 15496 1360 15502
rect 1308 15438 1360 15444
rect 1320 14958 1348 15438
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1320 13326 1348 14894
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 12782 1348 13262
rect 1308 12776 1360 12782
rect 1308 12718 1360 12724
rect 1320 10062 1348 12718
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1412 9081 1440 16546
rect 1780 14362 1808 31962
rect 2044 29844 2096 29850
rect 2044 29786 2096 29792
rect 1952 28212 2004 28218
rect 1952 28154 2004 28160
rect 1860 26784 1912 26790
rect 1860 26726 1912 26732
rect 1872 26382 1900 26726
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1596 14334 1808 14362
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 10810 1532 11698
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 9722 1532 10610
rect 1596 10062 1624 14334
rect 1674 14104 1730 14113
rect 1872 14056 1900 26318
rect 1964 15008 1992 28154
rect 2056 15502 2084 29786
rect 2136 21412 2188 21418
rect 2136 21354 2188 21360
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2044 15020 2096 15026
rect 1964 14980 2044 15008
rect 2044 14962 2096 14968
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 14074 2084 14214
rect 1674 14039 1730 14048
rect 1688 13326 1716 14039
rect 1780 14028 1900 14056
rect 2044 14068 2096 14074
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1780 12986 1808 14028
rect 2044 14010 2096 14016
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1872 12442 1900 13874
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13025 1992 13670
rect 2148 13326 2176 21354
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 1950 13016 2006 13025
rect 1950 12951 2006 12960
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1492 9172 1544 9178
rect 1596 9160 1624 9862
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1544 9132 1624 9160
rect 1492 9114 1544 9120
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1412 8906 1440 9007
rect 1400 8900 1452 8906
rect 1400 8842 1452 8848
rect 1504 6914 1532 9114
rect 2148 8634 2176 9318
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1582 8392 1638 8401
rect 1582 8327 1638 8336
rect 1860 8356 1912 8362
rect 1596 8090 1624 8327
rect 1860 8298 1912 8304
rect 1872 8265 1900 8298
rect 2136 8288 2188 8294
rect 1858 8256 1914 8265
rect 2136 8230 2188 8236
rect 1858 8191 1914 8200
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 2148 7886 2176 8230
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 7002 2176 7346
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 1412 6886 1532 6914
rect 1412 6798 1440 6886
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5710 1440 6734
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1216 2644 1268 2650
rect 1216 2586 1268 2592
rect 1596 1358 1624 5510
rect 2056 4622 2084 6054
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2240 2038 2268 35866
rect 2332 6914 2360 38984
rect 2412 30048 2464 30054
rect 2412 29990 2464 29996
rect 2424 29850 2452 29990
rect 2412 29844 2464 29850
rect 2412 29786 2464 29792
rect 2516 22114 2544 43250
rect 2663 43004 2971 43013
rect 2663 43002 2669 43004
rect 2725 43002 2749 43004
rect 2805 43002 2829 43004
rect 2885 43002 2909 43004
rect 2965 43002 2971 43004
rect 2725 42950 2727 43002
rect 2907 42950 2909 43002
rect 2663 42948 2669 42950
rect 2725 42948 2749 42950
rect 2805 42948 2829 42950
rect 2885 42948 2909 42950
rect 2965 42948 2971 42950
rect 2663 42939 2971 42948
rect 3068 42906 3096 43250
rect 3804 42906 3832 43250
rect 4356 42906 4384 43250
rect 3056 42900 3108 42906
rect 3056 42842 3108 42848
rect 3792 42900 3844 42906
rect 3792 42842 3844 42848
rect 4344 42900 4396 42906
rect 4344 42842 4396 42848
rect 2964 42696 3016 42702
rect 2964 42638 3016 42644
rect 3516 42696 3568 42702
rect 3516 42638 3568 42644
rect 2976 42362 3004 42638
rect 2964 42356 3016 42362
rect 2964 42298 3016 42304
rect 3056 42220 3108 42226
rect 3056 42162 3108 42168
rect 2663 41916 2971 41925
rect 2663 41914 2669 41916
rect 2725 41914 2749 41916
rect 2805 41914 2829 41916
rect 2885 41914 2909 41916
rect 2965 41914 2971 41916
rect 2725 41862 2727 41914
rect 2907 41862 2909 41914
rect 2663 41860 2669 41862
rect 2725 41860 2749 41862
rect 2805 41860 2829 41862
rect 2885 41860 2909 41862
rect 2965 41860 2971 41862
rect 2663 41851 2971 41860
rect 3068 41818 3096 42162
rect 3240 42084 3292 42090
rect 3240 42026 3292 42032
rect 3056 41812 3108 41818
rect 3056 41754 3108 41760
rect 2663 40828 2971 40837
rect 2663 40826 2669 40828
rect 2725 40826 2749 40828
rect 2805 40826 2829 40828
rect 2885 40826 2909 40828
rect 2965 40826 2971 40828
rect 2725 40774 2727 40826
rect 2907 40774 2909 40826
rect 2663 40772 2669 40774
rect 2725 40772 2749 40774
rect 2805 40772 2829 40774
rect 2885 40772 2909 40774
rect 2965 40772 2971 40774
rect 2663 40763 2971 40772
rect 2663 39740 2971 39749
rect 2663 39738 2669 39740
rect 2725 39738 2749 39740
rect 2805 39738 2829 39740
rect 2885 39738 2909 39740
rect 2965 39738 2971 39740
rect 2725 39686 2727 39738
rect 2907 39686 2909 39738
rect 2663 39684 2669 39686
rect 2725 39684 2749 39686
rect 2805 39684 2829 39686
rect 2885 39684 2909 39686
rect 2965 39684 2971 39686
rect 2663 39675 2971 39684
rect 2663 38652 2971 38661
rect 2663 38650 2669 38652
rect 2725 38650 2749 38652
rect 2805 38650 2829 38652
rect 2885 38650 2909 38652
rect 2965 38650 2971 38652
rect 2725 38598 2727 38650
rect 2907 38598 2909 38650
rect 2663 38596 2669 38598
rect 2725 38596 2749 38598
rect 2805 38596 2829 38598
rect 2885 38596 2909 38598
rect 2965 38596 2971 38598
rect 2663 38587 2971 38596
rect 2663 37564 2971 37573
rect 2663 37562 2669 37564
rect 2725 37562 2749 37564
rect 2805 37562 2829 37564
rect 2885 37562 2909 37564
rect 2965 37562 2971 37564
rect 2725 37510 2727 37562
rect 2907 37510 2909 37562
rect 2663 37508 2669 37510
rect 2725 37508 2749 37510
rect 2805 37508 2829 37510
rect 2885 37508 2909 37510
rect 2965 37508 2971 37510
rect 2663 37499 2971 37508
rect 2663 36476 2971 36485
rect 2663 36474 2669 36476
rect 2725 36474 2749 36476
rect 2805 36474 2829 36476
rect 2885 36474 2909 36476
rect 2965 36474 2971 36476
rect 2725 36422 2727 36474
rect 2907 36422 2909 36474
rect 2663 36420 2669 36422
rect 2725 36420 2749 36422
rect 2805 36420 2829 36422
rect 2885 36420 2909 36422
rect 2965 36420 2971 36422
rect 2663 36411 2971 36420
rect 2663 35388 2971 35397
rect 2663 35386 2669 35388
rect 2725 35386 2749 35388
rect 2805 35386 2829 35388
rect 2885 35386 2909 35388
rect 2965 35386 2971 35388
rect 2725 35334 2727 35386
rect 2907 35334 2909 35386
rect 2663 35332 2669 35334
rect 2725 35332 2749 35334
rect 2805 35332 2829 35334
rect 2885 35332 2909 35334
rect 2965 35332 2971 35334
rect 2663 35323 2971 35332
rect 2663 34300 2971 34309
rect 2663 34298 2669 34300
rect 2725 34298 2749 34300
rect 2805 34298 2829 34300
rect 2885 34298 2909 34300
rect 2965 34298 2971 34300
rect 2725 34246 2727 34298
rect 2907 34246 2909 34298
rect 2663 34244 2669 34246
rect 2725 34244 2749 34246
rect 2805 34244 2829 34246
rect 2885 34244 2909 34246
rect 2965 34244 2971 34246
rect 2663 34235 2971 34244
rect 2663 33212 2971 33221
rect 2663 33210 2669 33212
rect 2725 33210 2749 33212
rect 2805 33210 2829 33212
rect 2885 33210 2909 33212
rect 2965 33210 2971 33212
rect 2725 33158 2727 33210
rect 2907 33158 2909 33210
rect 2663 33156 2669 33158
rect 2725 33156 2749 33158
rect 2805 33156 2829 33158
rect 2885 33156 2909 33158
rect 2965 33156 2971 33158
rect 2663 33147 2971 33156
rect 2663 32124 2971 32133
rect 2663 32122 2669 32124
rect 2725 32122 2749 32124
rect 2805 32122 2829 32124
rect 2885 32122 2909 32124
rect 2965 32122 2971 32124
rect 2725 32070 2727 32122
rect 2907 32070 2909 32122
rect 2663 32068 2669 32070
rect 2725 32068 2749 32070
rect 2805 32068 2829 32070
rect 2885 32068 2909 32070
rect 2965 32068 2971 32070
rect 2663 32059 2971 32068
rect 2663 31036 2971 31045
rect 2663 31034 2669 31036
rect 2725 31034 2749 31036
rect 2805 31034 2829 31036
rect 2885 31034 2909 31036
rect 2965 31034 2971 31036
rect 2725 30982 2727 31034
rect 2907 30982 2909 31034
rect 2663 30980 2669 30982
rect 2725 30980 2749 30982
rect 2805 30980 2829 30982
rect 2885 30980 2909 30982
rect 2965 30980 2971 30982
rect 2663 30971 2971 30980
rect 2663 29948 2971 29957
rect 2663 29946 2669 29948
rect 2725 29946 2749 29948
rect 2805 29946 2829 29948
rect 2885 29946 2909 29948
rect 2965 29946 2971 29948
rect 2725 29894 2727 29946
rect 2907 29894 2909 29946
rect 2663 29892 2669 29894
rect 2725 29892 2749 29894
rect 2805 29892 2829 29894
rect 2885 29892 2909 29894
rect 2965 29892 2971 29894
rect 2663 29883 2971 29892
rect 2663 28860 2971 28869
rect 2663 28858 2669 28860
rect 2725 28858 2749 28860
rect 2805 28858 2829 28860
rect 2885 28858 2909 28860
rect 2965 28858 2971 28860
rect 2725 28806 2727 28858
rect 2907 28806 2909 28858
rect 2663 28804 2669 28806
rect 2725 28804 2749 28806
rect 2805 28804 2829 28806
rect 2885 28804 2909 28806
rect 2965 28804 2971 28806
rect 2663 28795 2971 28804
rect 2663 27772 2971 27781
rect 2663 27770 2669 27772
rect 2725 27770 2749 27772
rect 2805 27770 2829 27772
rect 2885 27770 2909 27772
rect 2965 27770 2971 27772
rect 2725 27718 2727 27770
rect 2907 27718 2909 27770
rect 2663 27716 2669 27718
rect 2725 27716 2749 27718
rect 2805 27716 2829 27718
rect 2885 27716 2909 27718
rect 2965 27716 2971 27718
rect 2663 27707 2971 27716
rect 2663 26684 2971 26693
rect 2663 26682 2669 26684
rect 2725 26682 2749 26684
rect 2805 26682 2829 26684
rect 2885 26682 2909 26684
rect 2965 26682 2971 26684
rect 2725 26630 2727 26682
rect 2907 26630 2909 26682
rect 2663 26628 2669 26630
rect 2725 26628 2749 26630
rect 2805 26628 2829 26630
rect 2885 26628 2909 26630
rect 2965 26628 2971 26630
rect 2663 26619 2971 26628
rect 2663 25596 2971 25605
rect 2663 25594 2669 25596
rect 2725 25594 2749 25596
rect 2805 25594 2829 25596
rect 2885 25594 2909 25596
rect 2965 25594 2971 25596
rect 2725 25542 2727 25594
rect 2907 25542 2909 25594
rect 2663 25540 2669 25542
rect 2725 25540 2749 25542
rect 2805 25540 2829 25542
rect 2885 25540 2909 25542
rect 2965 25540 2971 25542
rect 2663 25531 2971 25540
rect 2663 24508 2971 24517
rect 2663 24506 2669 24508
rect 2725 24506 2749 24508
rect 2805 24506 2829 24508
rect 2885 24506 2909 24508
rect 2965 24506 2971 24508
rect 2725 24454 2727 24506
rect 2907 24454 2909 24506
rect 2663 24452 2669 24454
rect 2725 24452 2749 24454
rect 2805 24452 2829 24454
rect 2885 24452 2909 24454
rect 2965 24452 2971 24454
rect 2663 24443 2971 24452
rect 2663 23420 2971 23429
rect 2663 23418 2669 23420
rect 2725 23418 2749 23420
rect 2805 23418 2829 23420
rect 2885 23418 2909 23420
rect 2965 23418 2971 23420
rect 2725 23366 2727 23418
rect 2907 23366 2909 23418
rect 2663 23364 2669 23366
rect 2725 23364 2749 23366
rect 2805 23364 2829 23366
rect 2885 23364 2909 23366
rect 2965 23364 2971 23366
rect 2663 23355 2971 23364
rect 2663 22332 2971 22341
rect 2663 22330 2669 22332
rect 2725 22330 2749 22332
rect 2805 22330 2829 22332
rect 2885 22330 2909 22332
rect 2965 22330 2971 22332
rect 2725 22278 2727 22330
rect 2907 22278 2909 22330
rect 2663 22276 2669 22278
rect 2725 22276 2749 22278
rect 2805 22276 2829 22278
rect 2885 22276 2909 22278
rect 2965 22276 2971 22278
rect 2663 22267 2971 22276
rect 2516 22086 2728 22114
rect 2700 21690 2728 22086
rect 3148 22024 3200 22030
rect 3148 21966 3200 21972
rect 3160 21690 3188 21966
rect 2688 21684 2740 21690
rect 2688 21626 2740 21632
rect 3148 21684 3200 21690
rect 3148 21626 3200 21632
rect 2663 21244 2971 21253
rect 2663 21242 2669 21244
rect 2725 21242 2749 21244
rect 2805 21242 2829 21244
rect 2885 21242 2909 21244
rect 2965 21242 2971 21244
rect 2725 21190 2727 21242
rect 2907 21190 2909 21242
rect 2663 21188 2669 21190
rect 2725 21188 2749 21190
rect 2805 21188 2829 21190
rect 2885 21188 2909 21190
rect 2965 21188 2971 21190
rect 2663 21179 2971 21188
rect 2663 20156 2971 20165
rect 2663 20154 2669 20156
rect 2725 20154 2749 20156
rect 2805 20154 2829 20156
rect 2885 20154 2909 20156
rect 2965 20154 2971 20156
rect 2725 20102 2727 20154
rect 2907 20102 2909 20154
rect 2663 20100 2669 20102
rect 2725 20100 2749 20102
rect 2805 20100 2829 20102
rect 2885 20100 2909 20102
rect 2965 20100 2971 20102
rect 2663 20091 2971 20100
rect 2663 19068 2971 19077
rect 2663 19066 2669 19068
rect 2725 19066 2749 19068
rect 2805 19066 2829 19068
rect 2885 19066 2909 19068
rect 2965 19066 2971 19068
rect 2725 19014 2727 19066
rect 2907 19014 2909 19066
rect 2663 19012 2669 19014
rect 2725 19012 2749 19014
rect 2805 19012 2829 19014
rect 2885 19012 2909 19014
rect 2965 19012 2971 19014
rect 2663 19003 2971 19012
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 16590 2544 18090
rect 2663 17980 2971 17989
rect 2663 17978 2669 17980
rect 2725 17978 2749 17980
rect 2805 17978 2829 17980
rect 2885 17978 2909 17980
rect 2965 17978 2971 17980
rect 2725 17926 2727 17978
rect 2907 17926 2909 17978
rect 2663 17924 2669 17926
rect 2725 17924 2749 17926
rect 2805 17924 2829 17926
rect 2885 17924 2909 17926
rect 2965 17924 2971 17926
rect 2663 17915 2971 17924
rect 2663 16892 2971 16901
rect 2663 16890 2669 16892
rect 2725 16890 2749 16892
rect 2805 16890 2829 16892
rect 2885 16890 2909 16892
rect 2965 16890 2971 16892
rect 2725 16838 2727 16890
rect 2907 16838 2909 16890
rect 2663 16836 2669 16838
rect 2725 16836 2749 16838
rect 2805 16836 2829 16838
rect 2885 16836 2909 16838
rect 2965 16836 2971 16838
rect 2663 16827 2971 16836
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2516 15502 2544 15846
rect 2663 15804 2971 15813
rect 2663 15802 2669 15804
rect 2725 15802 2749 15804
rect 2805 15802 2829 15804
rect 2885 15802 2909 15804
rect 2965 15802 2971 15804
rect 2725 15750 2727 15802
rect 2907 15750 2909 15802
rect 2663 15748 2669 15750
rect 2725 15748 2749 15750
rect 2805 15748 2829 15750
rect 2885 15748 2909 15750
rect 2965 15748 2971 15750
rect 2663 15739 2971 15748
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2504 15360 2556 15366
rect 2504 15302 2556 15308
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 14618 2452 14758
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2516 14414 2544 15302
rect 2663 14716 2971 14725
rect 2663 14714 2669 14716
rect 2725 14714 2749 14716
rect 2805 14714 2829 14716
rect 2885 14714 2909 14716
rect 2965 14714 2971 14716
rect 2725 14662 2727 14714
rect 2907 14662 2909 14714
rect 2663 14660 2669 14662
rect 2725 14660 2749 14662
rect 2805 14660 2829 14662
rect 2885 14660 2909 14662
rect 2965 14660 2971 14662
rect 2663 14651 2971 14660
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 2504 13728 2556 13734
rect 2502 13696 2504 13705
rect 2556 13696 2558 13705
rect 2502 13631 2558 13640
rect 2663 13628 2971 13637
rect 2663 13626 2669 13628
rect 2725 13626 2749 13628
rect 2805 13626 2829 13628
rect 2885 13626 2909 13628
rect 2965 13626 2971 13628
rect 2725 13574 2727 13626
rect 2907 13574 2909 13626
rect 2663 13572 2669 13574
rect 2725 13572 2749 13574
rect 2805 13572 2829 13574
rect 2885 13572 2909 13574
rect 2965 13572 2971 13574
rect 2663 13563 2971 13572
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12238 2452 12582
rect 2516 12238 2544 13126
rect 2663 12540 2971 12549
rect 2663 12538 2669 12540
rect 2725 12538 2749 12540
rect 2805 12538 2829 12540
rect 2885 12538 2909 12540
rect 2965 12538 2971 12540
rect 2725 12486 2727 12538
rect 2907 12486 2909 12538
rect 2663 12484 2669 12486
rect 2725 12484 2749 12486
rect 2805 12484 2829 12486
rect 2885 12484 2909 12486
rect 2965 12484 2971 12486
rect 2663 12475 2971 12484
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2663 11452 2971 11461
rect 2663 11450 2669 11452
rect 2725 11450 2749 11452
rect 2805 11450 2829 11452
rect 2885 11450 2909 11452
rect 2965 11450 2971 11452
rect 2725 11398 2727 11450
rect 2907 11398 2909 11450
rect 2663 11396 2669 11398
rect 2725 11396 2749 11398
rect 2805 11396 2829 11398
rect 2885 11396 2909 11398
rect 2965 11396 2971 11398
rect 2663 11387 2971 11396
rect 2663 10364 2971 10373
rect 2663 10362 2669 10364
rect 2725 10362 2749 10364
rect 2805 10362 2829 10364
rect 2885 10362 2909 10364
rect 2965 10362 2971 10364
rect 2725 10310 2727 10362
rect 2907 10310 2909 10362
rect 2663 10308 2669 10310
rect 2725 10308 2749 10310
rect 2805 10308 2829 10310
rect 2885 10308 2909 10310
rect 2965 10308 2971 10310
rect 2663 10299 2971 10308
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9586 2452 9862
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2663 9276 2971 9285
rect 2663 9274 2669 9276
rect 2725 9274 2749 9276
rect 2805 9274 2829 9276
rect 2885 9274 2909 9276
rect 2965 9274 2971 9276
rect 2725 9222 2727 9274
rect 2907 9222 2909 9274
rect 2663 9220 2669 9222
rect 2725 9220 2749 9222
rect 2805 9220 2829 9222
rect 2885 9220 2909 9222
rect 2965 9220 2971 9222
rect 2663 9211 2971 9220
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8634 2452 8774
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2663 8188 2971 8197
rect 2663 8186 2669 8188
rect 2725 8186 2749 8188
rect 2805 8186 2829 8188
rect 2885 8186 2909 8188
rect 2965 8186 2971 8188
rect 2725 8134 2727 8186
rect 2907 8134 2909 8186
rect 2663 8132 2669 8134
rect 2725 8132 2749 8134
rect 2805 8132 2829 8134
rect 2885 8132 2909 8134
rect 2965 8132 2971 8134
rect 2663 8123 2971 8132
rect 2663 7100 2971 7109
rect 2663 7098 2669 7100
rect 2725 7098 2749 7100
rect 2805 7098 2829 7100
rect 2885 7098 2909 7100
rect 2965 7098 2971 7100
rect 2725 7046 2727 7098
rect 2907 7046 2909 7098
rect 2663 7044 2669 7046
rect 2725 7044 2749 7046
rect 2805 7044 2829 7046
rect 2885 7044 2909 7046
rect 2965 7044 2971 7046
rect 2663 7035 2971 7044
rect 2332 6886 2452 6914
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 1308 1352 1360 1358
rect 1308 1294 1360 1300
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 1320 160 1348 1294
rect 570 0 626 160
rect 1306 0 1362 160
rect 2042 82 2098 160
rect 2148 82 2176 1906
rect 2424 1766 2452 6886
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5914 2544 6258
rect 2663 6012 2971 6021
rect 2663 6010 2669 6012
rect 2725 6010 2749 6012
rect 2805 6010 2829 6012
rect 2885 6010 2909 6012
rect 2965 6010 2971 6012
rect 2725 5958 2727 6010
rect 2907 5958 2909 6010
rect 2663 5956 2669 5958
rect 2725 5956 2749 5958
rect 2805 5956 2829 5958
rect 2885 5956 2909 5958
rect 2965 5956 2971 5958
rect 2663 5947 2971 5956
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2663 4924 2971 4933
rect 2663 4922 2669 4924
rect 2725 4922 2749 4924
rect 2805 4922 2829 4924
rect 2885 4922 2909 4924
rect 2965 4922 2971 4924
rect 2725 4870 2727 4922
rect 2907 4870 2909 4922
rect 2663 4868 2669 4870
rect 2725 4868 2749 4870
rect 2805 4868 2829 4870
rect 2885 4868 2909 4870
rect 2965 4868 2971 4870
rect 2663 4859 2971 4868
rect 2663 3836 2971 3845
rect 2663 3834 2669 3836
rect 2725 3834 2749 3836
rect 2805 3834 2829 3836
rect 2885 3834 2909 3836
rect 2965 3834 2971 3836
rect 2725 3782 2727 3834
rect 2907 3782 2909 3834
rect 2663 3780 2669 3782
rect 2725 3780 2749 3782
rect 2805 3780 2829 3782
rect 2885 3780 2909 3782
rect 2965 3780 2971 3782
rect 2663 3771 2971 3780
rect 2663 2748 2971 2757
rect 2663 2746 2669 2748
rect 2725 2746 2749 2748
rect 2805 2746 2829 2748
rect 2885 2746 2909 2748
rect 2965 2746 2971 2748
rect 2725 2694 2727 2746
rect 2907 2694 2909 2746
rect 2663 2692 2669 2694
rect 2725 2692 2749 2694
rect 2805 2692 2829 2694
rect 2885 2692 2909 2694
rect 2965 2692 2971 2694
rect 2663 2683 2971 2692
rect 3252 1834 3280 42026
rect 3528 22094 3556 42638
rect 4376 42460 4684 42469
rect 4376 42458 4382 42460
rect 4438 42458 4462 42460
rect 4518 42458 4542 42460
rect 4598 42458 4622 42460
rect 4678 42458 4684 42460
rect 4438 42406 4440 42458
rect 4620 42406 4622 42458
rect 4376 42404 4382 42406
rect 4438 42404 4462 42406
rect 4518 42404 4542 42406
rect 4598 42404 4622 42406
rect 4678 42404 4684 42406
rect 4376 42395 4684 42404
rect 3608 42152 3660 42158
rect 3608 42094 3660 42100
rect 3344 22066 3556 22094
rect 3344 21894 3372 22066
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3344 6225 3372 19654
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3330 6216 3386 6225
rect 3330 6151 3386 6160
rect 3436 3942 3464 19110
rect 3620 14618 3648 42094
rect 4376 41372 4684 41381
rect 4376 41370 4382 41372
rect 4438 41370 4462 41372
rect 4518 41370 4542 41372
rect 4598 41370 4622 41372
rect 4678 41370 4684 41372
rect 4438 41318 4440 41370
rect 4620 41318 4622 41370
rect 4376 41316 4382 41318
rect 4438 41316 4462 41318
rect 4518 41316 4542 41318
rect 4598 41316 4622 41318
rect 4678 41316 4684 41318
rect 4376 41307 4684 41316
rect 4376 40284 4684 40293
rect 4376 40282 4382 40284
rect 4438 40282 4462 40284
rect 4518 40282 4542 40284
rect 4598 40282 4622 40284
rect 4678 40282 4684 40284
rect 4438 40230 4440 40282
rect 4620 40230 4622 40282
rect 4376 40228 4382 40230
rect 4438 40228 4462 40230
rect 4518 40228 4542 40230
rect 4598 40228 4622 40230
rect 4678 40228 4684 40230
rect 4376 40219 4684 40228
rect 4376 39196 4684 39205
rect 4376 39194 4382 39196
rect 4438 39194 4462 39196
rect 4518 39194 4542 39196
rect 4598 39194 4622 39196
rect 4678 39194 4684 39196
rect 4438 39142 4440 39194
rect 4620 39142 4622 39194
rect 4376 39140 4382 39142
rect 4438 39140 4462 39142
rect 4518 39140 4542 39142
rect 4598 39140 4622 39142
rect 4678 39140 4684 39142
rect 4376 39131 4684 39140
rect 5092 39098 5120 43250
rect 5828 42906 5856 43250
rect 6090 43004 6398 43013
rect 6090 43002 6096 43004
rect 6152 43002 6176 43004
rect 6232 43002 6256 43004
rect 6312 43002 6336 43004
rect 6392 43002 6398 43004
rect 6152 42950 6154 43002
rect 6334 42950 6336 43002
rect 6090 42948 6096 42950
rect 6152 42948 6176 42950
rect 6232 42948 6256 42950
rect 6312 42948 6336 42950
rect 6392 42948 6398 42950
rect 6090 42939 6398 42948
rect 6564 42906 6592 43250
rect 7300 42906 7328 43250
rect 8036 42906 8064 43250
rect 8956 42906 8984 43250
rect 9324 42906 9352 43250
rect 9517 43004 9825 43013
rect 9517 43002 9523 43004
rect 9579 43002 9603 43004
rect 9659 43002 9683 43004
rect 9739 43002 9763 43004
rect 9819 43002 9825 43004
rect 9579 42950 9581 43002
rect 9761 42950 9763 43002
rect 9517 42948 9523 42950
rect 9579 42948 9603 42950
rect 9659 42948 9683 42950
rect 9739 42948 9763 42950
rect 9819 42948 9825 42950
rect 9517 42939 9825 42948
rect 10244 42906 10272 43250
rect 11624 42906 11652 43250
rect 11716 43110 11744 43438
rect 12348 43444 12400 43450
rect 12348 43386 12400 43392
rect 13084 43444 13136 43450
rect 13084 43386 13136 43392
rect 13820 43444 13872 43450
rect 13820 43386 13872 43392
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 12532 43308 12584 43314
rect 12532 43250 12584 43256
rect 13268 43308 13320 43314
rect 13268 43250 13320 43256
rect 13636 43308 13688 43314
rect 13636 43250 13688 43256
rect 14096 43308 14148 43314
rect 14096 43250 14148 43256
rect 11704 43104 11756 43110
rect 11704 43046 11756 43052
rect 12084 42906 12112 43250
rect 12544 42906 12572 43250
rect 12944 43004 13252 43013
rect 12944 43002 12950 43004
rect 13006 43002 13030 43004
rect 13086 43002 13110 43004
rect 13166 43002 13190 43004
rect 13246 43002 13252 43004
rect 13006 42950 13008 43002
rect 13188 42950 13190 43002
rect 12944 42948 12950 42950
rect 13006 42948 13030 42950
rect 13086 42948 13110 42950
rect 13166 42948 13190 42950
rect 13246 42948 13252 42950
rect 12944 42939 13252 42948
rect 13280 42906 13308 43250
rect 13648 42906 13676 43250
rect 14108 42906 14136 43250
rect 14568 43246 14596 44463
rect 14657 43548 14965 43557
rect 14657 43546 14663 43548
rect 14719 43546 14743 43548
rect 14799 43546 14823 43548
rect 14879 43546 14903 43548
rect 14959 43546 14965 43548
rect 14719 43494 14721 43546
rect 14901 43494 14903 43546
rect 14657 43492 14663 43494
rect 14719 43492 14743 43494
rect 14799 43492 14823 43494
rect 14879 43492 14903 43494
rect 14959 43492 14965 43494
rect 14657 43483 14965 43492
rect 14556 43240 14608 43246
rect 14556 43182 14608 43188
rect 5816 42900 5868 42906
rect 5816 42842 5868 42848
rect 6552 42900 6604 42906
rect 6552 42842 6604 42848
rect 7288 42900 7340 42906
rect 7288 42842 7340 42848
rect 8024 42900 8076 42906
rect 8024 42842 8076 42848
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 9312 42900 9364 42906
rect 9312 42842 9364 42848
rect 10232 42900 10284 42906
rect 10232 42842 10284 42848
rect 11612 42900 11664 42906
rect 11612 42842 11664 42848
rect 12072 42900 12124 42906
rect 12072 42842 12124 42848
rect 12532 42900 12584 42906
rect 12532 42842 12584 42848
rect 13268 42900 13320 42906
rect 13268 42842 13320 42848
rect 13636 42900 13688 42906
rect 13636 42842 13688 42848
rect 14096 42900 14148 42906
rect 14096 42842 14148 42848
rect 15304 42770 15332 44463
rect 15292 42764 15344 42770
rect 15292 42706 15344 42712
rect 5908 42696 5960 42702
rect 5908 42638 5960 42644
rect 6644 42696 6696 42702
rect 6644 42638 6696 42644
rect 7288 42696 7340 42702
rect 7288 42638 7340 42644
rect 8208 42696 8260 42702
rect 8208 42638 8260 42644
rect 8760 42696 8812 42702
rect 8760 42638 8812 42644
rect 9496 42696 9548 42702
rect 9496 42638 9548 42644
rect 10232 42696 10284 42702
rect 10232 42638 10284 42644
rect 10968 42696 11020 42702
rect 10968 42638 11020 42644
rect 11704 42696 11756 42702
rect 11704 42638 11756 42644
rect 12440 42696 12492 42702
rect 12440 42638 12492 42644
rect 13176 42696 13228 42702
rect 13176 42638 13228 42644
rect 14096 42696 14148 42702
rect 14096 42638 14148 42644
rect 5920 42362 5948 42638
rect 6656 42362 6684 42638
rect 7300 42362 7328 42638
rect 7803 42460 8111 42469
rect 7803 42458 7809 42460
rect 7865 42458 7889 42460
rect 7945 42458 7969 42460
rect 8025 42458 8049 42460
rect 8105 42458 8111 42460
rect 7865 42406 7867 42458
rect 8047 42406 8049 42458
rect 7803 42404 7809 42406
rect 7865 42404 7889 42406
rect 7945 42404 7969 42406
rect 8025 42404 8049 42406
rect 8105 42404 8111 42406
rect 7803 42395 8111 42404
rect 8220 42362 8248 42638
rect 8772 42362 8800 42638
rect 9508 42362 9536 42638
rect 10244 42362 10272 42638
rect 10980 42362 11008 42638
rect 11230 42460 11538 42469
rect 11230 42458 11236 42460
rect 11292 42458 11316 42460
rect 11372 42458 11396 42460
rect 11452 42458 11476 42460
rect 11532 42458 11538 42460
rect 11292 42406 11294 42458
rect 11474 42406 11476 42458
rect 11230 42404 11236 42406
rect 11292 42404 11316 42406
rect 11372 42404 11396 42406
rect 11452 42404 11476 42406
rect 11532 42404 11538 42406
rect 11230 42395 11538 42404
rect 11716 42362 11744 42638
rect 12452 42362 12480 42638
rect 13188 42362 13216 42638
rect 13544 42628 13596 42634
rect 13544 42570 13596 42576
rect 13556 42362 13584 42570
rect 5908 42356 5960 42362
rect 5908 42298 5960 42304
rect 6644 42356 6696 42362
rect 6644 42298 6696 42304
rect 7288 42356 7340 42362
rect 7288 42298 7340 42304
rect 8208 42356 8260 42362
rect 8208 42298 8260 42304
rect 8760 42356 8812 42362
rect 8760 42298 8812 42304
rect 9496 42356 9548 42362
rect 9496 42298 9548 42304
rect 10232 42356 10284 42362
rect 10232 42298 10284 42304
rect 10968 42356 11020 42362
rect 10968 42298 11020 42304
rect 11704 42356 11756 42362
rect 11704 42298 11756 42304
rect 12440 42356 12492 42362
rect 12440 42298 12492 42304
rect 13176 42356 13228 42362
rect 13176 42298 13228 42304
rect 13544 42356 13596 42362
rect 13544 42298 13596 42304
rect 14108 42294 14136 42638
rect 14280 42560 14332 42566
rect 14280 42502 14332 42508
rect 14292 42362 14320 42502
rect 14657 42460 14965 42469
rect 14657 42458 14663 42460
rect 14719 42458 14743 42460
rect 14799 42458 14823 42460
rect 14879 42458 14903 42460
rect 14959 42458 14965 42460
rect 14719 42406 14721 42458
rect 14901 42406 14903 42458
rect 14657 42404 14663 42406
rect 14719 42404 14743 42406
rect 14799 42404 14823 42406
rect 14879 42404 14903 42406
rect 14959 42404 14965 42406
rect 14657 42395 14965 42404
rect 14280 42356 14332 42362
rect 14280 42298 14332 42304
rect 14096 42288 14148 42294
rect 14096 42230 14148 42236
rect 5724 42220 5776 42226
rect 5724 42162 5776 42168
rect 6552 42220 6604 42226
rect 6552 42162 6604 42168
rect 7288 42220 7340 42226
rect 7288 42162 7340 42168
rect 8116 42220 8168 42226
rect 8116 42162 8168 42168
rect 10968 42220 11020 42226
rect 10968 42162 11020 42168
rect 11704 42220 11756 42226
rect 11704 42162 11756 42168
rect 12440 42220 12492 42226
rect 12440 42162 12492 42168
rect 14004 42220 14056 42226
rect 14004 42162 14056 42168
rect 14188 42220 14240 42226
rect 14188 42162 14240 42168
rect 15752 42220 15804 42226
rect 15752 42162 15804 42168
rect 5736 41857 5764 42162
rect 6090 41916 6398 41925
rect 6090 41914 6096 41916
rect 6152 41914 6176 41916
rect 6232 41914 6256 41916
rect 6312 41914 6336 41916
rect 6392 41914 6398 41916
rect 6152 41862 6154 41914
rect 6334 41862 6336 41914
rect 6090 41860 6096 41862
rect 6152 41860 6176 41862
rect 6232 41860 6256 41862
rect 6312 41860 6336 41862
rect 6392 41860 6398 41862
rect 5722 41848 5778 41857
rect 6090 41851 6398 41860
rect 6564 41857 6592 42162
rect 5722 41783 5778 41792
rect 6550 41848 6606 41857
rect 6550 41783 6606 41792
rect 6920 41608 6972 41614
rect 7300 41585 7328 42162
rect 8128 41857 8156 42162
rect 9517 41916 9825 41925
rect 9517 41914 9523 41916
rect 9579 41914 9603 41916
rect 9659 41914 9683 41916
rect 9739 41914 9763 41916
rect 9819 41914 9825 41916
rect 9579 41862 9581 41914
rect 9761 41862 9763 41914
rect 9517 41860 9523 41862
rect 9579 41860 9603 41862
rect 9659 41860 9683 41862
rect 9739 41860 9763 41862
rect 9819 41860 9825 41862
rect 8114 41848 8170 41857
rect 9517 41851 9825 41860
rect 10980 41857 11008 42162
rect 11716 42129 11744 42162
rect 11702 42120 11758 42129
rect 11702 42055 11758 42064
rect 8114 41783 8170 41792
rect 10966 41848 11022 41857
rect 10966 41783 11022 41792
rect 12452 41585 12480 42162
rect 12944 41916 13252 41925
rect 12944 41914 12950 41916
rect 13006 41914 13030 41916
rect 13086 41914 13110 41916
rect 13166 41914 13190 41916
rect 13246 41914 13252 41916
rect 13006 41862 13008 41914
rect 13188 41862 13190 41914
rect 12944 41860 12950 41862
rect 13006 41860 13030 41862
rect 13086 41860 13110 41862
rect 13166 41860 13190 41862
rect 13246 41860 13252 41862
rect 12944 41851 13252 41860
rect 14016 41682 14044 42162
rect 14200 41818 14228 42162
rect 15108 42016 15160 42022
rect 15108 41958 15160 41964
rect 14188 41812 14240 41818
rect 14188 41754 14240 41760
rect 14004 41676 14056 41682
rect 14004 41618 14056 41624
rect 15016 41676 15068 41682
rect 15016 41618 15068 41624
rect 6920 41550 6972 41556
rect 7286 41576 7342 41585
rect 6090 40828 6398 40837
rect 6090 40826 6096 40828
rect 6152 40826 6176 40828
rect 6232 40826 6256 40828
rect 6312 40826 6336 40828
rect 6392 40826 6398 40828
rect 6152 40774 6154 40826
rect 6334 40774 6336 40826
rect 6090 40772 6096 40774
rect 6152 40772 6176 40774
rect 6232 40772 6256 40774
rect 6312 40772 6336 40774
rect 6392 40772 6398 40774
rect 6090 40763 6398 40772
rect 6090 39740 6398 39749
rect 6090 39738 6096 39740
rect 6152 39738 6176 39740
rect 6232 39738 6256 39740
rect 6312 39738 6336 39740
rect 6392 39738 6398 39740
rect 6152 39686 6154 39738
rect 6334 39686 6336 39738
rect 6090 39684 6096 39686
rect 6152 39684 6176 39686
rect 6232 39684 6256 39686
rect 6312 39684 6336 39686
rect 6392 39684 6398 39686
rect 6090 39675 6398 39684
rect 5080 39092 5132 39098
rect 5080 39034 5132 39040
rect 5172 38956 5224 38962
rect 5172 38898 5224 38904
rect 5184 38554 5212 38898
rect 6090 38652 6398 38661
rect 6090 38650 6096 38652
rect 6152 38650 6176 38652
rect 6232 38650 6256 38652
rect 6312 38650 6336 38652
rect 6392 38650 6398 38652
rect 6152 38598 6154 38650
rect 6334 38598 6336 38650
rect 6090 38596 6096 38598
rect 6152 38596 6176 38598
rect 6232 38596 6256 38598
rect 6312 38596 6336 38598
rect 6392 38596 6398 38598
rect 6090 38587 6398 38596
rect 5172 38548 5224 38554
rect 5172 38490 5224 38496
rect 4376 38108 4684 38117
rect 4376 38106 4382 38108
rect 4438 38106 4462 38108
rect 4518 38106 4542 38108
rect 4598 38106 4622 38108
rect 4678 38106 4684 38108
rect 4438 38054 4440 38106
rect 4620 38054 4622 38106
rect 4376 38052 4382 38054
rect 4438 38052 4462 38054
rect 4518 38052 4542 38054
rect 4598 38052 4622 38054
rect 4678 38052 4684 38054
rect 4376 38043 4684 38052
rect 5724 37664 5776 37670
rect 5724 37606 5776 37612
rect 6552 37664 6604 37670
rect 6552 37606 6604 37612
rect 4376 37020 4684 37029
rect 4376 37018 4382 37020
rect 4438 37018 4462 37020
rect 4518 37018 4542 37020
rect 4598 37018 4622 37020
rect 4678 37018 4684 37020
rect 4438 36966 4440 37018
rect 4620 36966 4622 37018
rect 4376 36964 4382 36966
rect 4438 36964 4462 36966
rect 4518 36964 4542 36966
rect 4598 36964 4622 36966
rect 4678 36964 4684 36966
rect 4376 36955 4684 36964
rect 4252 36780 4304 36786
rect 4252 36722 4304 36728
rect 3700 33652 3752 33658
rect 3700 33594 3752 33600
rect 3712 18737 3740 33594
rect 3792 30592 3844 30598
rect 3792 30534 3844 30540
rect 3804 28422 3832 30534
rect 3884 30116 3936 30122
rect 3884 30058 3936 30064
rect 3896 29578 3924 30058
rect 4264 29714 4292 36722
rect 5172 36712 5224 36718
rect 5172 36654 5224 36660
rect 4376 35932 4684 35941
rect 4376 35930 4382 35932
rect 4438 35930 4462 35932
rect 4518 35930 4542 35932
rect 4598 35930 4622 35932
rect 4678 35930 4684 35932
rect 4438 35878 4440 35930
rect 4620 35878 4622 35930
rect 4376 35876 4382 35878
rect 4438 35876 4462 35878
rect 4518 35876 4542 35878
rect 4598 35876 4622 35878
rect 4678 35876 4684 35878
rect 4376 35867 4684 35876
rect 4376 34844 4684 34853
rect 4376 34842 4382 34844
rect 4438 34842 4462 34844
rect 4518 34842 4542 34844
rect 4598 34842 4622 34844
rect 4678 34842 4684 34844
rect 4438 34790 4440 34842
rect 4620 34790 4622 34842
rect 4376 34788 4382 34790
rect 4438 34788 4462 34790
rect 4518 34788 4542 34790
rect 4598 34788 4622 34790
rect 4678 34788 4684 34790
rect 4376 34779 4684 34788
rect 4804 34672 4856 34678
rect 4804 34614 4856 34620
rect 4376 33756 4684 33765
rect 4376 33754 4382 33756
rect 4438 33754 4462 33756
rect 4518 33754 4542 33756
rect 4598 33754 4622 33756
rect 4678 33754 4684 33756
rect 4438 33702 4440 33754
rect 4620 33702 4622 33754
rect 4376 33700 4382 33702
rect 4438 33700 4462 33702
rect 4518 33700 4542 33702
rect 4598 33700 4622 33702
rect 4678 33700 4684 33702
rect 4376 33691 4684 33700
rect 4376 32668 4684 32677
rect 4376 32666 4382 32668
rect 4438 32666 4462 32668
rect 4518 32666 4542 32668
rect 4598 32666 4622 32668
rect 4678 32666 4684 32668
rect 4438 32614 4440 32666
rect 4620 32614 4622 32666
rect 4376 32612 4382 32614
rect 4438 32612 4462 32614
rect 4518 32612 4542 32614
rect 4598 32612 4622 32614
rect 4678 32612 4684 32614
rect 4376 32603 4684 32612
rect 4376 31580 4684 31589
rect 4376 31578 4382 31580
rect 4438 31578 4462 31580
rect 4518 31578 4542 31580
rect 4598 31578 4622 31580
rect 4678 31578 4684 31580
rect 4438 31526 4440 31578
rect 4620 31526 4622 31578
rect 4376 31524 4382 31526
rect 4438 31524 4462 31526
rect 4518 31524 4542 31526
rect 4598 31524 4622 31526
rect 4678 31524 4684 31526
rect 4376 31515 4684 31524
rect 4376 30492 4684 30501
rect 4376 30490 4382 30492
rect 4438 30490 4462 30492
rect 4518 30490 4542 30492
rect 4598 30490 4622 30492
rect 4678 30490 4684 30492
rect 4438 30438 4440 30490
rect 4620 30438 4622 30490
rect 4376 30436 4382 30438
rect 4438 30436 4462 30438
rect 4518 30436 4542 30438
rect 4598 30436 4622 30438
rect 4678 30436 4684 30438
rect 4376 30427 4684 30436
rect 4252 29708 4304 29714
rect 4252 29650 4304 29656
rect 3884 29572 3936 29578
rect 3884 29514 3936 29520
rect 3792 28416 3844 28422
rect 3792 28358 3844 28364
rect 3698 18728 3754 18737
rect 3698 18663 3754 18672
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3804 11830 3832 28358
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3896 11150 3924 29514
rect 4376 29404 4684 29413
rect 4376 29402 4382 29404
rect 4438 29402 4462 29404
rect 4518 29402 4542 29404
rect 4598 29402 4622 29404
rect 4678 29402 4684 29404
rect 4438 29350 4440 29402
rect 4620 29350 4622 29402
rect 4376 29348 4382 29350
rect 4438 29348 4462 29350
rect 4518 29348 4542 29350
rect 4598 29348 4622 29350
rect 4678 29348 4684 29350
rect 4376 29339 4684 29348
rect 3974 29200 4030 29209
rect 3974 29135 4030 29144
rect 3988 17678 4016 29135
rect 4376 28316 4684 28325
rect 4376 28314 4382 28316
rect 4438 28314 4462 28316
rect 4518 28314 4542 28316
rect 4598 28314 4622 28316
rect 4678 28314 4684 28316
rect 4438 28262 4440 28314
rect 4620 28262 4622 28314
rect 4376 28260 4382 28262
rect 4438 28260 4462 28262
rect 4518 28260 4542 28262
rect 4598 28260 4622 28262
rect 4678 28260 4684 28262
rect 4376 28251 4684 28260
rect 4376 27228 4684 27237
rect 4376 27226 4382 27228
rect 4438 27226 4462 27228
rect 4518 27226 4542 27228
rect 4598 27226 4622 27228
rect 4678 27226 4684 27228
rect 4438 27174 4440 27226
rect 4620 27174 4622 27226
rect 4376 27172 4382 27174
rect 4438 27172 4462 27174
rect 4518 27172 4542 27174
rect 4598 27172 4622 27174
rect 4678 27172 4684 27174
rect 4376 27163 4684 27172
rect 4068 26240 4120 26246
rect 4068 26182 4120 26188
rect 4080 19310 4108 26182
rect 4376 26140 4684 26149
rect 4376 26138 4382 26140
rect 4438 26138 4462 26140
rect 4518 26138 4542 26140
rect 4598 26138 4622 26140
rect 4678 26138 4684 26140
rect 4438 26086 4440 26138
rect 4620 26086 4622 26138
rect 4376 26084 4382 26086
rect 4438 26084 4462 26086
rect 4518 26084 4542 26086
rect 4598 26084 4622 26086
rect 4678 26084 4684 26086
rect 4376 26075 4684 26084
rect 4376 25052 4684 25061
rect 4376 25050 4382 25052
rect 4438 25050 4462 25052
rect 4518 25050 4542 25052
rect 4598 25050 4622 25052
rect 4678 25050 4684 25052
rect 4438 24998 4440 25050
rect 4620 24998 4622 25050
rect 4376 24996 4382 24998
rect 4438 24996 4462 24998
rect 4518 24996 4542 24998
rect 4598 24996 4622 24998
rect 4678 24996 4684 24998
rect 4376 24987 4684 24996
rect 4376 23964 4684 23973
rect 4376 23962 4382 23964
rect 4438 23962 4462 23964
rect 4518 23962 4542 23964
rect 4598 23962 4622 23964
rect 4678 23962 4684 23964
rect 4438 23910 4440 23962
rect 4620 23910 4622 23962
rect 4376 23908 4382 23910
rect 4438 23908 4462 23910
rect 4518 23908 4542 23910
rect 4598 23908 4622 23910
rect 4678 23908 4684 23910
rect 4376 23899 4684 23908
rect 4252 23112 4304 23118
rect 4252 23054 4304 23060
rect 4264 22098 4292 23054
rect 4376 22876 4684 22885
rect 4376 22874 4382 22876
rect 4438 22874 4462 22876
rect 4518 22874 4542 22876
rect 4598 22874 4622 22876
rect 4678 22874 4684 22876
rect 4438 22822 4440 22874
rect 4620 22822 4622 22874
rect 4376 22820 4382 22822
rect 4438 22820 4462 22822
rect 4518 22820 4542 22822
rect 4598 22820 4622 22822
rect 4678 22820 4684 22822
rect 4376 22811 4684 22820
rect 4252 22092 4304 22098
rect 4252 22034 4304 22040
rect 4376 21788 4684 21797
rect 4376 21786 4382 21788
rect 4438 21786 4462 21788
rect 4518 21786 4542 21788
rect 4598 21786 4622 21788
rect 4678 21786 4684 21788
rect 4438 21734 4440 21786
rect 4620 21734 4622 21786
rect 4376 21732 4382 21734
rect 4438 21732 4462 21734
rect 4518 21732 4542 21734
rect 4598 21732 4622 21734
rect 4678 21732 4684 21734
rect 4376 21723 4684 21732
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4172 21010 4200 21558
rect 4160 21004 4212 21010
rect 4160 20946 4212 20952
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4172 18290 4200 20946
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4264 20466 4292 20810
rect 4376 20700 4684 20709
rect 4376 20698 4382 20700
rect 4438 20698 4462 20700
rect 4518 20698 4542 20700
rect 4598 20698 4622 20700
rect 4678 20698 4684 20700
rect 4438 20646 4440 20698
rect 4620 20646 4622 20698
rect 4376 20644 4382 20646
rect 4438 20644 4462 20646
rect 4518 20644 4542 20646
rect 4598 20644 4622 20646
rect 4678 20644 4684 20646
rect 4376 20635 4684 20644
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4264 19174 4292 20402
rect 4376 19612 4684 19621
rect 4376 19610 4382 19612
rect 4438 19610 4462 19612
rect 4518 19610 4542 19612
rect 4598 19610 4622 19612
rect 4678 19610 4684 19612
rect 4438 19558 4440 19610
rect 4620 19558 4622 19610
rect 4376 19556 4382 19558
rect 4438 19556 4462 19558
rect 4518 19556 4542 19558
rect 4598 19556 4622 19558
rect 4678 19556 4684 19558
rect 4376 19547 4684 19556
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4816 18698 4844 34614
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4376 18524 4684 18533
rect 4376 18522 4382 18524
rect 4438 18522 4462 18524
rect 4518 18522 4542 18524
rect 4598 18522 4622 18524
rect 4678 18522 4684 18524
rect 4438 18470 4440 18522
rect 4620 18470 4622 18522
rect 4376 18468 4382 18470
rect 4438 18468 4462 18470
rect 4518 18468 4542 18470
rect 4598 18468 4622 18470
rect 4678 18468 4684 18470
rect 4376 18459 4684 18468
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 4448 17610 4476 18226
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 4172 9654 4200 17546
rect 4376 17436 4684 17445
rect 4376 17434 4382 17436
rect 4438 17434 4462 17436
rect 4518 17434 4542 17436
rect 4598 17434 4622 17436
rect 4678 17434 4684 17436
rect 4438 17382 4440 17434
rect 4620 17382 4622 17434
rect 4376 17380 4382 17382
rect 4438 17380 4462 17382
rect 4518 17380 4542 17382
rect 4598 17380 4622 17382
rect 4678 17380 4684 17382
rect 4376 17371 4684 17380
rect 4376 16348 4684 16357
rect 4376 16346 4382 16348
rect 4438 16346 4462 16348
rect 4518 16346 4542 16348
rect 4598 16346 4622 16348
rect 4678 16346 4684 16348
rect 4438 16294 4440 16346
rect 4620 16294 4622 16346
rect 4376 16292 4382 16294
rect 4438 16292 4462 16294
rect 4518 16292 4542 16294
rect 4598 16292 4622 16294
rect 4678 16292 4684 16294
rect 4376 16283 4684 16292
rect 4376 15260 4684 15269
rect 4376 15258 4382 15260
rect 4438 15258 4462 15260
rect 4518 15258 4542 15260
rect 4598 15258 4622 15260
rect 4678 15258 4684 15260
rect 4438 15206 4440 15258
rect 4620 15206 4622 15258
rect 4376 15204 4382 15206
rect 4438 15204 4462 15206
rect 4518 15204 4542 15206
rect 4598 15204 4622 15206
rect 4678 15204 4684 15206
rect 4376 15195 4684 15204
rect 4376 14172 4684 14181
rect 4376 14170 4382 14172
rect 4438 14170 4462 14172
rect 4518 14170 4542 14172
rect 4598 14170 4622 14172
rect 4678 14170 4684 14172
rect 4438 14118 4440 14170
rect 4620 14118 4622 14170
rect 4376 14116 4382 14118
rect 4438 14116 4462 14118
rect 4518 14116 4542 14118
rect 4598 14116 4622 14118
rect 4678 14116 4684 14118
rect 4376 14107 4684 14116
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 10742 4292 13262
rect 4376 13084 4684 13093
rect 4376 13082 4382 13084
rect 4438 13082 4462 13084
rect 4518 13082 4542 13084
rect 4598 13082 4622 13084
rect 4678 13082 4684 13084
rect 4438 13030 4440 13082
rect 4620 13030 4622 13082
rect 4376 13028 4382 13030
rect 4438 13028 4462 13030
rect 4518 13028 4542 13030
rect 4598 13028 4622 13030
rect 4678 13028 4684 13030
rect 4376 13019 4684 13028
rect 4376 11996 4684 12005
rect 4376 11994 4382 11996
rect 4438 11994 4462 11996
rect 4518 11994 4542 11996
rect 4598 11994 4622 11996
rect 4678 11994 4684 11996
rect 4438 11942 4440 11994
rect 4620 11942 4622 11994
rect 4376 11940 4382 11942
rect 4438 11940 4462 11942
rect 4518 11940 4542 11942
rect 4598 11940 4622 11942
rect 4678 11940 4684 11942
rect 4376 11931 4684 11940
rect 4376 10908 4684 10917
rect 4376 10906 4382 10908
rect 4438 10906 4462 10908
rect 4518 10906 4542 10908
rect 4598 10906 4622 10908
rect 4678 10906 4684 10908
rect 4438 10854 4440 10906
rect 4620 10854 4622 10906
rect 4376 10852 4382 10854
rect 4438 10852 4462 10854
rect 4518 10852 4542 10854
rect 4598 10852 4622 10854
rect 4678 10852 4684 10854
rect 4376 10843 4684 10852
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4376 9820 4684 9829
rect 4376 9818 4382 9820
rect 4438 9818 4462 9820
rect 4518 9818 4542 9820
rect 4598 9818 4622 9820
rect 4678 9818 4684 9820
rect 4438 9766 4440 9818
rect 4620 9766 4622 9818
rect 4376 9764 4382 9766
rect 4438 9764 4462 9766
rect 4518 9764 4542 9766
rect 4598 9764 4622 9766
rect 4678 9764 4684 9766
rect 4376 9755 4684 9764
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 5234 4016 9318
rect 4376 8732 4684 8741
rect 4376 8730 4382 8732
rect 4438 8730 4462 8732
rect 4518 8730 4542 8732
rect 4598 8730 4622 8732
rect 4678 8730 4684 8732
rect 4438 8678 4440 8730
rect 4620 8678 4622 8730
rect 4376 8676 4382 8678
rect 4438 8676 4462 8678
rect 4518 8676 4542 8678
rect 4598 8676 4622 8678
rect 4678 8676 4684 8678
rect 4376 8667 4684 8676
rect 4816 7750 4844 18634
rect 4896 17740 4948 17746
rect 4896 17682 4948 17688
rect 4908 17202 4936 17682
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16794 4936 16934
rect 4896 16788 4948 16794
rect 4896 16730 4948 16736
rect 5000 12442 5028 23802
rect 5184 23118 5212 36654
rect 5446 35592 5502 35601
rect 5446 35527 5502 35536
rect 5460 34678 5488 35527
rect 5448 34672 5500 34678
rect 5448 34614 5500 34620
rect 5736 31754 5764 37606
rect 6090 37564 6398 37573
rect 6090 37562 6096 37564
rect 6152 37562 6176 37564
rect 6232 37562 6256 37564
rect 6312 37562 6336 37564
rect 6392 37562 6398 37564
rect 6152 37510 6154 37562
rect 6334 37510 6336 37562
rect 6090 37508 6096 37510
rect 6152 37508 6176 37510
rect 6232 37508 6256 37510
rect 6312 37508 6336 37510
rect 6392 37508 6398 37510
rect 6090 37499 6398 37508
rect 6564 37194 6592 37606
rect 6552 37188 6604 37194
rect 6552 37130 6604 37136
rect 6090 36476 6398 36485
rect 6090 36474 6096 36476
rect 6152 36474 6176 36476
rect 6232 36474 6256 36476
rect 6312 36474 6336 36476
rect 6392 36474 6398 36476
rect 6152 36422 6154 36474
rect 6334 36422 6336 36474
rect 6090 36420 6096 36422
rect 6152 36420 6176 36422
rect 6232 36420 6256 36422
rect 6312 36420 6336 36422
rect 6392 36420 6398 36422
rect 6090 36411 6398 36420
rect 6090 35388 6398 35397
rect 6090 35386 6096 35388
rect 6152 35386 6176 35388
rect 6232 35386 6256 35388
rect 6312 35386 6336 35388
rect 6392 35386 6398 35388
rect 6152 35334 6154 35386
rect 6334 35334 6336 35386
rect 6090 35332 6096 35334
rect 6152 35332 6176 35334
rect 6232 35332 6256 35334
rect 6312 35332 6336 35334
rect 6392 35332 6398 35334
rect 6090 35323 6398 35332
rect 5908 35148 5960 35154
rect 5908 35090 5960 35096
rect 5816 34604 5868 34610
rect 5816 34546 5868 34552
rect 5644 31726 5764 31754
rect 5448 31340 5500 31346
rect 5448 31282 5500 31288
rect 5356 30932 5408 30938
rect 5356 30874 5408 30880
rect 5264 29028 5316 29034
rect 5264 28970 5316 28976
rect 5172 23112 5224 23118
rect 5172 23054 5224 23060
rect 5080 22636 5132 22642
rect 5080 22578 5132 22584
rect 5092 21690 5120 22578
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5184 19514 5212 23054
rect 5276 20505 5304 28970
rect 5262 20496 5318 20505
rect 5262 20431 5318 20440
rect 5368 19666 5396 30874
rect 5460 26382 5488 31282
rect 5540 29708 5592 29714
rect 5540 29650 5592 29656
rect 5552 28762 5580 29650
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 5460 25294 5488 26318
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5460 22098 5488 23258
rect 5448 22092 5500 22098
rect 5448 22034 5500 22040
rect 5552 21842 5580 27066
rect 5644 22030 5672 31726
rect 5828 29646 5856 34546
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 5736 23118 5764 25230
rect 5828 23118 5856 25230
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5828 22438 5856 23054
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5552 21814 5764 21842
rect 5540 21684 5592 21690
rect 5540 21626 5592 21632
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 21146 5488 21286
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5446 19952 5502 19961
rect 5446 19887 5502 19896
rect 5276 19638 5396 19666
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5276 17354 5304 19638
rect 5460 19530 5488 19887
rect 5184 17326 5304 17354
rect 5368 19502 5488 19530
rect 5184 16590 5212 17326
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 15502 5212 16526
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5276 13433 5304 17138
rect 5262 13424 5318 13433
rect 5262 13359 5318 13368
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5368 10742 5396 19502
rect 5552 19394 5580 21626
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5644 21010 5672 21490
rect 5632 21004 5684 21010
rect 5632 20946 5684 20952
rect 5644 20466 5672 20946
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5644 19718 5672 20402
rect 5736 19854 5764 21814
rect 5920 21400 5948 35090
rect 6460 34536 6512 34542
rect 6460 34478 6512 34484
rect 6090 34300 6398 34309
rect 6090 34298 6096 34300
rect 6152 34298 6176 34300
rect 6232 34298 6256 34300
rect 6312 34298 6336 34300
rect 6392 34298 6398 34300
rect 6152 34246 6154 34298
rect 6334 34246 6336 34298
rect 6090 34244 6096 34246
rect 6152 34244 6176 34246
rect 6232 34244 6256 34246
rect 6312 34244 6336 34246
rect 6392 34244 6398 34246
rect 6090 34235 6398 34244
rect 6472 33658 6500 34478
rect 6460 33652 6512 33658
rect 6460 33594 6512 33600
rect 6460 33448 6512 33454
rect 6460 33390 6512 33396
rect 6090 33212 6398 33221
rect 6090 33210 6096 33212
rect 6152 33210 6176 33212
rect 6232 33210 6256 33212
rect 6312 33210 6336 33212
rect 6392 33210 6398 33212
rect 6152 33158 6154 33210
rect 6334 33158 6336 33210
rect 6090 33156 6096 33158
rect 6152 33156 6176 33158
rect 6232 33156 6256 33158
rect 6312 33156 6336 33158
rect 6392 33156 6398 33158
rect 6090 33147 6398 33156
rect 6090 32124 6398 32133
rect 6090 32122 6096 32124
rect 6152 32122 6176 32124
rect 6232 32122 6256 32124
rect 6312 32122 6336 32124
rect 6392 32122 6398 32124
rect 6152 32070 6154 32122
rect 6334 32070 6336 32122
rect 6090 32068 6096 32070
rect 6152 32068 6176 32070
rect 6232 32068 6256 32070
rect 6312 32068 6336 32070
rect 6392 32068 6398 32070
rect 6090 32059 6398 32068
rect 6090 31036 6398 31045
rect 6090 31034 6096 31036
rect 6152 31034 6176 31036
rect 6232 31034 6256 31036
rect 6312 31034 6336 31036
rect 6392 31034 6398 31036
rect 6152 30982 6154 31034
rect 6334 30982 6336 31034
rect 6090 30980 6096 30982
rect 6152 30980 6176 30982
rect 6232 30980 6256 30982
rect 6312 30980 6336 30982
rect 6392 30980 6398 30982
rect 6090 30971 6398 30980
rect 6090 29948 6398 29957
rect 6090 29946 6096 29948
rect 6152 29946 6176 29948
rect 6232 29946 6256 29948
rect 6312 29946 6336 29948
rect 6392 29946 6398 29948
rect 6152 29894 6154 29946
rect 6334 29894 6336 29946
rect 6090 29892 6096 29894
rect 6152 29892 6176 29894
rect 6232 29892 6256 29894
rect 6312 29892 6336 29894
rect 6392 29892 6398 29894
rect 6090 29883 6398 29892
rect 6090 28860 6398 28869
rect 6090 28858 6096 28860
rect 6152 28858 6176 28860
rect 6232 28858 6256 28860
rect 6312 28858 6336 28860
rect 6392 28858 6398 28860
rect 6152 28806 6154 28858
rect 6334 28806 6336 28858
rect 6090 28804 6096 28806
rect 6152 28804 6176 28806
rect 6232 28804 6256 28806
rect 6312 28804 6336 28806
rect 6392 28804 6398 28806
rect 6090 28795 6398 28804
rect 6000 28756 6052 28762
rect 6000 28698 6052 28704
rect 6012 27470 6040 28698
rect 6090 27772 6398 27781
rect 6090 27770 6096 27772
rect 6152 27770 6176 27772
rect 6232 27770 6256 27772
rect 6312 27770 6336 27772
rect 6392 27770 6398 27772
rect 6152 27718 6154 27770
rect 6334 27718 6336 27770
rect 6090 27716 6096 27718
rect 6152 27716 6176 27718
rect 6232 27716 6256 27718
rect 6312 27716 6336 27718
rect 6392 27716 6398 27718
rect 6090 27707 6398 27716
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6012 26382 6040 27406
rect 6472 27334 6500 33390
rect 6932 31890 6960 41550
rect 7286 41511 7342 41520
rect 12438 41576 12494 41585
rect 12438 41511 12494 41520
rect 7803 41372 8111 41381
rect 7803 41370 7809 41372
rect 7865 41370 7889 41372
rect 7945 41370 7969 41372
rect 8025 41370 8049 41372
rect 8105 41370 8111 41372
rect 7865 41318 7867 41370
rect 8047 41318 8049 41370
rect 7803 41316 7809 41318
rect 7865 41316 7889 41318
rect 7945 41316 7969 41318
rect 8025 41316 8049 41318
rect 8105 41316 8111 41318
rect 7803 41307 8111 41316
rect 11230 41372 11538 41381
rect 11230 41370 11236 41372
rect 11292 41370 11316 41372
rect 11372 41370 11396 41372
rect 11452 41370 11476 41372
rect 11532 41370 11538 41372
rect 11292 41318 11294 41370
rect 11474 41318 11476 41370
rect 11230 41316 11236 41318
rect 11292 41316 11316 41318
rect 11372 41316 11396 41318
rect 11452 41316 11476 41318
rect 11532 41316 11538 41318
rect 11230 41307 11538 41316
rect 14657 41372 14965 41381
rect 14657 41370 14663 41372
rect 14719 41370 14743 41372
rect 14799 41370 14823 41372
rect 14879 41370 14903 41372
rect 14959 41370 14965 41372
rect 14719 41318 14721 41370
rect 14901 41318 14903 41370
rect 14657 41316 14663 41318
rect 14719 41316 14743 41318
rect 14799 41316 14823 41318
rect 14879 41316 14903 41318
rect 14959 41316 14965 41318
rect 14657 41307 14965 41316
rect 8208 40928 8260 40934
rect 8208 40870 8260 40876
rect 7803 40284 8111 40293
rect 7803 40282 7809 40284
rect 7865 40282 7889 40284
rect 7945 40282 7969 40284
rect 8025 40282 8049 40284
rect 8105 40282 8111 40284
rect 7865 40230 7867 40282
rect 8047 40230 8049 40282
rect 7803 40228 7809 40230
rect 7865 40228 7889 40230
rect 7945 40228 7969 40230
rect 8025 40228 8049 40230
rect 8105 40228 8111 40230
rect 7803 40219 8111 40228
rect 7380 39840 7432 39846
rect 7380 39782 7432 39788
rect 7392 39370 7420 39782
rect 8220 39420 8248 40870
rect 9517 40828 9825 40837
rect 9517 40826 9523 40828
rect 9579 40826 9603 40828
rect 9659 40826 9683 40828
rect 9739 40826 9763 40828
rect 9819 40826 9825 40828
rect 9579 40774 9581 40826
rect 9761 40774 9763 40826
rect 9517 40772 9523 40774
rect 9579 40772 9603 40774
rect 9659 40772 9683 40774
rect 9739 40772 9763 40774
rect 9819 40772 9825 40774
rect 9517 40763 9825 40772
rect 12944 40828 13252 40837
rect 12944 40826 12950 40828
rect 13006 40826 13030 40828
rect 13086 40826 13110 40828
rect 13166 40826 13190 40828
rect 13246 40826 13252 40828
rect 13006 40774 13008 40826
rect 13188 40774 13190 40826
rect 12944 40772 12950 40774
rect 13006 40772 13030 40774
rect 13086 40772 13110 40774
rect 13166 40772 13190 40774
rect 13246 40772 13252 40774
rect 12944 40763 13252 40772
rect 11230 40284 11538 40293
rect 11230 40282 11236 40284
rect 11292 40282 11316 40284
rect 11372 40282 11396 40284
rect 11452 40282 11476 40284
rect 11532 40282 11538 40284
rect 11292 40230 11294 40282
rect 11474 40230 11476 40282
rect 11230 40228 11236 40230
rect 11292 40228 11316 40230
rect 11372 40228 11396 40230
rect 11452 40228 11476 40230
rect 11532 40228 11538 40230
rect 11230 40219 11538 40228
rect 14657 40284 14965 40293
rect 14657 40282 14663 40284
rect 14719 40282 14743 40284
rect 14799 40282 14823 40284
rect 14879 40282 14903 40284
rect 14959 40282 14965 40284
rect 14719 40230 14721 40282
rect 14901 40230 14903 40282
rect 14657 40228 14663 40230
rect 14719 40228 14743 40230
rect 14799 40228 14823 40230
rect 14879 40228 14903 40230
rect 14959 40228 14965 40230
rect 14657 40219 14965 40228
rect 13360 40044 13412 40050
rect 13360 39986 13412 39992
rect 10968 39976 11020 39982
rect 10968 39918 11020 39924
rect 9517 39740 9825 39749
rect 9517 39738 9523 39740
rect 9579 39738 9603 39740
rect 9659 39738 9683 39740
rect 9739 39738 9763 39740
rect 9819 39738 9825 39740
rect 9579 39686 9581 39738
rect 9761 39686 9763 39738
rect 9517 39684 9523 39686
rect 9579 39684 9603 39686
rect 9659 39684 9683 39686
rect 9739 39684 9763 39686
rect 9819 39684 9825 39686
rect 9517 39675 9825 39684
rect 10980 39642 11008 39918
rect 12944 39740 13252 39749
rect 12944 39738 12950 39740
rect 13006 39738 13030 39740
rect 13086 39738 13110 39740
rect 13166 39738 13190 39740
rect 13246 39738 13252 39740
rect 13006 39686 13008 39738
rect 13188 39686 13190 39738
rect 12944 39684 12950 39686
rect 13006 39684 13030 39686
rect 13086 39684 13110 39686
rect 13166 39684 13190 39686
rect 13246 39684 13252 39686
rect 12944 39675 13252 39684
rect 13372 39642 13400 39986
rect 14004 39840 14056 39846
rect 14004 39782 14056 39788
rect 14188 39840 14240 39846
rect 14188 39782 14240 39788
rect 10968 39636 11020 39642
rect 10968 39578 11020 39584
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 14016 39545 14044 39782
rect 14200 39545 14228 39782
rect 14002 39536 14058 39545
rect 14002 39471 14058 39480
rect 14186 39536 14242 39545
rect 14186 39471 14242 39480
rect 8392 39432 8444 39438
rect 8220 39392 8392 39420
rect 7380 39364 7432 39370
rect 7380 39306 7432 39312
rect 7286 37224 7342 37233
rect 7286 37159 7342 37168
rect 7300 36378 7328 37159
rect 7288 36372 7340 36378
rect 7288 36314 7340 36320
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 7012 33380 7064 33386
rect 7012 33322 7064 33328
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6932 30546 6960 31826
rect 6840 30518 6960 30546
rect 6840 30326 6868 30518
rect 7024 30410 7052 33322
rect 7116 32434 7144 33934
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 6932 30382 7052 30410
rect 7104 30388 7156 30394
rect 6828 30320 6880 30326
rect 6828 30262 6880 30268
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 6736 29504 6788 29510
rect 6736 29446 6788 29452
rect 6564 29306 6592 29446
rect 6552 29300 6604 29306
rect 6552 29242 6604 29248
rect 6748 29102 6776 29446
rect 6840 29102 6868 29582
rect 6736 29096 6788 29102
rect 6736 29038 6788 29044
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6644 27872 6696 27878
rect 6644 27814 6696 27820
rect 6460 27328 6512 27334
rect 6460 27270 6512 27276
rect 6090 26684 6398 26693
rect 6090 26682 6096 26684
rect 6152 26682 6176 26684
rect 6232 26682 6256 26684
rect 6312 26682 6336 26684
rect 6392 26682 6398 26684
rect 6152 26630 6154 26682
rect 6334 26630 6336 26682
rect 6090 26628 6096 26630
rect 6152 26628 6176 26630
rect 6232 26628 6256 26630
rect 6312 26628 6336 26630
rect 6392 26628 6398 26630
rect 6090 26619 6398 26628
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6380 25838 6408 26318
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6090 25596 6398 25605
rect 6090 25594 6096 25596
rect 6152 25594 6176 25596
rect 6232 25594 6256 25596
rect 6312 25594 6336 25596
rect 6392 25594 6398 25596
rect 6152 25542 6154 25594
rect 6334 25542 6336 25594
rect 6090 25540 6096 25542
rect 6152 25540 6176 25542
rect 6232 25540 6256 25542
rect 6312 25540 6336 25542
rect 6392 25540 6398 25542
rect 6090 25531 6398 25540
rect 6368 25492 6420 25498
rect 6472 25480 6500 27270
rect 6656 26042 6684 27814
rect 6748 26994 6776 29038
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6840 26790 6868 29038
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6736 26376 6788 26382
rect 6932 26364 6960 30382
rect 7104 30330 7156 30336
rect 7012 30252 7064 30258
rect 7012 30194 7064 30200
rect 6788 26336 6960 26364
rect 6736 26318 6788 26324
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6420 25452 6500 25480
rect 6368 25434 6420 25440
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 24410 6040 24686
rect 6090 24508 6398 24517
rect 6090 24506 6096 24508
rect 6152 24506 6176 24508
rect 6232 24506 6256 24508
rect 6312 24506 6336 24508
rect 6392 24506 6398 24508
rect 6152 24454 6154 24506
rect 6334 24454 6336 24506
rect 6090 24452 6096 24454
rect 6152 24452 6176 24454
rect 6232 24452 6256 24454
rect 6312 24452 6336 24454
rect 6392 24452 6398 24454
rect 6090 24443 6398 24452
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 6012 22642 6040 24346
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6380 23508 6408 24210
rect 6472 23730 6500 25452
rect 6552 25288 6604 25294
rect 6552 25230 6604 25236
rect 6460 23724 6512 23730
rect 6460 23666 6512 23672
rect 6380 23480 6500 23508
rect 6090 23420 6398 23429
rect 6090 23418 6096 23420
rect 6152 23418 6176 23420
rect 6232 23418 6256 23420
rect 6312 23418 6336 23420
rect 6392 23418 6398 23420
rect 6152 23366 6154 23418
rect 6334 23366 6336 23418
rect 6090 23364 6096 23366
rect 6152 23364 6176 23366
rect 6232 23364 6256 23366
rect 6312 23364 6336 23366
rect 6392 23364 6398 23366
rect 6090 23355 6398 23364
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 6090 22332 6398 22341
rect 6090 22330 6096 22332
rect 6152 22330 6176 22332
rect 6232 22330 6256 22332
rect 6312 22330 6336 22332
rect 6392 22330 6398 22332
rect 6152 22278 6154 22330
rect 6334 22278 6336 22330
rect 6090 22276 6096 22278
rect 6152 22276 6176 22278
rect 6232 22276 6256 22278
rect 6312 22276 6336 22278
rect 6392 22276 6398 22278
rect 6090 22267 6398 22276
rect 6472 22030 6500 23480
rect 6564 23186 6592 25230
rect 6656 25158 6684 25638
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6748 25158 6776 25230
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6656 24274 6684 25094
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6552 23180 6604 23186
rect 6552 23122 6604 23128
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 6288 21486 6316 21966
rect 6564 21690 6592 23122
rect 6656 23066 6684 24006
rect 6748 23186 6776 25094
rect 6840 24206 6868 26336
rect 6920 24268 6972 24274
rect 6920 24210 6972 24216
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6932 23662 6960 24210
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 23322 6960 23598
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6828 23112 6880 23118
rect 6656 23038 6776 23066
rect 6828 23054 6880 23060
rect 6644 22500 6696 22506
rect 6644 22442 6696 22448
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6276 21480 6328 21486
rect 6276 21422 6328 21428
rect 5828 21372 5948 21400
rect 5828 20942 5856 21372
rect 6656 21332 6684 22442
rect 5920 21304 6684 21332
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5460 19366 5580 19394
rect 5736 19378 5764 19790
rect 5632 19372 5684 19378
rect 5460 17746 5488 19366
rect 5632 19314 5684 19320
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5552 18426 5580 19246
rect 5644 18902 5672 19314
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18970 5764 19110
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5632 18896 5684 18902
rect 5828 18850 5856 20878
rect 5632 18838 5684 18844
rect 5736 18822 5856 18850
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 16658 5488 17682
rect 5644 17134 5672 18566
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5448 16652 5500 16658
rect 5500 16612 5580 16640
rect 5448 16594 5500 16600
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 13938 5488 15438
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5460 13530 5488 13874
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 11898 5580 16612
rect 5644 16522 5672 17070
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5644 15706 5672 16458
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5552 10538 5580 11834
rect 5644 11694 5672 13262
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11218 5672 11630
rect 5736 11354 5764 18822
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5828 18426 5856 18702
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5920 17728 5948 21304
rect 6090 21244 6398 21253
rect 6090 21242 6096 21244
rect 6152 21242 6176 21244
rect 6232 21242 6256 21244
rect 6312 21242 6336 21244
rect 6392 21242 6398 21244
rect 6152 21190 6154 21242
rect 6334 21190 6336 21242
rect 6090 21188 6096 21190
rect 6152 21188 6176 21190
rect 6232 21188 6256 21190
rect 6312 21188 6336 21190
rect 6392 21188 6398 21190
rect 6090 21179 6398 21188
rect 6748 21162 6776 23038
rect 6840 22234 6868 23054
rect 6920 22976 6972 22982
rect 6920 22918 6972 22924
rect 6932 22234 6960 22918
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 7024 22030 7052 30194
rect 7116 28422 7144 30330
rect 7196 30320 7248 30326
rect 7196 30262 7248 30268
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7208 27418 7236 30262
rect 7116 27390 7236 27418
rect 7116 24274 7144 27390
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7208 26926 7236 27270
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 7196 25900 7248 25906
rect 7196 25842 7248 25848
rect 7208 24410 7236 25842
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7104 24268 7156 24274
rect 7104 24210 7156 24216
rect 7208 23526 7236 24346
rect 7196 23520 7248 23526
rect 7196 23462 7248 23468
rect 7196 22636 7248 22642
rect 7196 22578 7248 22584
rect 6828 22024 6880 22030
rect 7012 22024 7064 22030
rect 6880 21984 6960 22012
rect 6828 21966 6880 21972
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6564 21134 6776 21162
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6000 20460 6052 20466
rect 6000 20402 6052 20408
rect 6012 20058 6040 20402
rect 6090 20156 6398 20165
rect 6090 20154 6096 20156
rect 6152 20154 6176 20156
rect 6232 20154 6256 20156
rect 6312 20154 6336 20156
rect 6392 20154 6398 20156
rect 6152 20102 6154 20154
rect 6334 20102 6336 20154
rect 6090 20100 6096 20102
rect 6152 20100 6176 20102
rect 6232 20100 6256 20102
rect 6312 20100 6336 20102
rect 6392 20100 6398 20102
rect 6090 20091 6398 20100
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6380 19854 6408 19994
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6012 18850 6040 19654
rect 6104 19378 6132 19790
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6090 19068 6398 19077
rect 6090 19066 6096 19068
rect 6152 19066 6176 19068
rect 6232 19066 6256 19068
rect 6312 19066 6336 19068
rect 6392 19066 6398 19068
rect 6152 19014 6154 19066
rect 6334 19014 6336 19066
rect 6090 19012 6096 19014
rect 6152 19012 6176 19014
rect 6232 19012 6256 19014
rect 6312 19012 6336 19014
rect 6392 19012 6398 19014
rect 6090 19003 6398 19012
rect 6012 18822 6224 18850
rect 6090 18728 6146 18737
rect 6196 18698 6224 18822
rect 6090 18663 6146 18672
rect 6184 18692 6236 18698
rect 6104 18630 6132 18663
rect 6184 18634 6236 18640
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6012 18426 6040 18566
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6104 18306 6132 18566
rect 6012 18278 6132 18306
rect 6012 17864 6040 18278
rect 6090 17980 6398 17989
rect 6090 17978 6096 17980
rect 6152 17978 6176 17980
rect 6232 17978 6256 17980
rect 6312 17978 6336 17980
rect 6392 17978 6398 17980
rect 6152 17926 6154 17978
rect 6334 17926 6336 17978
rect 6090 17924 6096 17926
rect 6152 17924 6176 17926
rect 6232 17924 6256 17926
rect 6312 17924 6336 17926
rect 6392 17924 6398 17926
rect 6090 17915 6398 17924
rect 6012 17836 6132 17864
rect 5828 17700 5948 17728
rect 5828 15194 5856 17700
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5920 17338 5948 17546
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 6104 17116 6132 17836
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6196 17134 6224 17682
rect 6012 17088 6132 17116
rect 6184 17128 6236 17134
rect 5828 15166 5948 15194
rect 5920 12209 5948 15166
rect 5906 12200 5962 12209
rect 5906 12135 5962 12144
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5276 10198 5304 10406
rect 5460 10198 5488 10406
rect 5264 10192 5316 10198
rect 5264 10134 5316 10140
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5552 10130 5580 10474
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5540 10124 5592 10130
rect 5592 10084 5764 10112
rect 5540 10066 5592 10072
rect 4986 9752 5042 9761
rect 5092 9722 5120 10066
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 4986 9687 5042 9696
rect 5080 9716 5132 9722
rect 5000 8566 5028 9687
rect 5080 9658 5132 9664
rect 5276 9518 5304 9862
rect 5368 9654 5396 9862
rect 5644 9722 5672 9930
rect 5736 9761 5764 10084
rect 5722 9752 5778 9761
rect 5632 9716 5684 9722
rect 5722 9687 5778 9696
rect 5632 9658 5684 9664
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4376 7644 4684 7653
rect 4376 7642 4382 7644
rect 4438 7642 4462 7644
rect 4518 7642 4542 7644
rect 4598 7642 4622 7644
rect 4678 7642 4684 7644
rect 4438 7590 4440 7642
rect 4620 7590 4622 7642
rect 4376 7588 4382 7590
rect 4438 7588 4462 7590
rect 4518 7588 4542 7590
rect 4598 7588 4622 7590
rect 4678 7588 4684 7590
rect 4376 7579 4684 7588
rect 5736 7410 5764 9687
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 4376 6556 4684 6565
rect 4376 6554 4382 6556
rect 4438 6554 4462 6556
rect 4518 6554 4542 6556
rect 4598 6554 4622 6556
rect 4678 6554 4684 6556
rect 4438 6502 4440 6554
rect 4620 6502 4622 6554
rect 4376 6500 4382 6502
rect 4438 6500 4462 6502
rect 4518 6500 4542 6502
rect 4598 6500 4622 6502
rect 4678 6500 4684 6502
rect 4376 6491 4684 6500
rect 5828 5574 5856 11086
rect 5920 9994 5948 12135
rect 6012 10248 6040 17088
rect 6184 17070 6236 17076
rect 6090 16892 6398 16901
rect 6090 16890 6096 16892
rect 6152 16890 6176 16892
rect 6232 16890 6256 16892
rect 6312 16890 6336 16892
rect 6392 16890 6398 16892
rect 6152 16838 6154 16890
rect 6334 16838 6336 16890
rect 6090 16836 6096 16838
rect 6152 16836 6176 16838
rect 6232 16836 6256 16838
rect 6312 16836 6336 16838
rect 6392 16836 6398 16838
rect 6090 16827 6398 16836
rect 6090 15804 6398 15813
rect 6090 15802 6096 15804
rect 6152 15802 6176 15804
rect 6232 15802 6256 15804
rect 6312 15802 6336 15804
rect 6392 15802 6398 15804
rect 6152 15750 6154 15802
rect 6334 15750 6336 15802
rect 6090 15748 6096 15750
rect 6152 15748 6176 15750
rect 6232 15748 6256 15750
rect 6312 15748 6336 15750
rect 6392 15748 6398 15750
rect 6090 15739 6398 15748
rect 6090 14716 6398 14725
rect 6090 14714 6096 14716
rect 6152 14714 6176 14716
rect 6232 14714 6256 14716
rect 6312 14714 6336 14716
rect 6392 14714 6398 14716
rect 6152 14662 6154 14714
rect 6334 14662 6336 14714
rect 6090 14660 6096 14662
rect 6152 14660 6176 14662
rect 6232 14660 6256 14662
rect 6312 14660 6336 14662
rect 6392 14660 6398 14662
rect 6090 14651 6398 14660
rect 6368 14408 6420 14414
rect 6368 14350 6420 14356
rect 6380 13938 6408 14350
rect 6472 14006 6500 20810
rect 6564 20602 6592 21134
rect 6644 20868 6696 20874
rect 6644 20810 6696 20816
rect 6552 20596 6604 20602
rect 6552 20538 6604 20544
rect 6564 19854 6592 20538
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6656 19310 6684 20810
rect 6736 20800 6788 20806
rect 6736 20742 6788 20748
rect 6748 20534 6776 20742
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6840 20482 6868 21422
rect 6932 21010 6960 21984
rect 7012 21966 7064 21972
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7024 20942 7052 21966
rect 7208 21706 7236 22578
rect 7300 21729 7328 36314
rect 7392 30258 7420 39306
rect 7564 39296 7616 39302
rect 7564 39238 7616 39244
rect 7576 39030 7604 39238
rect 7803 39196 8111 39205
rect 7803 39194 7809 39196
rect 7865 39194 7889 39196
rect 7945 39194 7969 39196
rect 8025 39194 8049 39196
rect 8105 39194 8111 39196
rect 7865 39142 7867 39194
rect 8047 39142 8049 39194
rect 7803 39140 7809 39142
rect 7865 39140 7889 39142
rect 7945 39140 7969 39142
rect 8025 39140 8049 39142
rect 8105 39140 8111 39142
rect 7803 39131 8111 39140
rect 7564 39024 7616 39030
rect 7564 38966 7616 38972
rect 7803 38108 8111 38117
rect 7803 38106 7809 38108
rect 7865 38106 7889 38108
rect 7945 38106 7969 38108
rect 8025 38106 8049 38108
rect 8105 38106 8111 38108
rect 7865 38054 7867 38106
rect 8047 38054 8049 38106
rect 7803 38052 7809 38054
rect 7865 38052 7889 38054
rect 7945 38052 7969 38054
rect 8025 38052 8049 38054
rect 8105 38052 8111 38054
rect 7803 38043 8111 38052
rect 7803 37020 8111 37029
rect 7803 37018 7809 37020
rect 7865 37018 7889 37020
rect 7945 37018 7969 37020
rect 8025 37018 8049 37020
rect 8105 37018 8111 37020
rect 7865 36966 7867 37018
rect 8047 36966 8049 37018
rect 7803 36964 7809 36966
rect 7865 36964 7889 36966
rect 7945 36964 7969 36966
rect 8025 36964 8049 36966
rect 8105 36964 8111 36966
rect 7803 36955 8111 36964
rect 7803 35932 8111 35941
rect 7803 35930 7809 35932
rect 7865 35930 7889 35932
rect 7945 35930 7969 35932
rect 8025 35930 8049 35932
rect 8105 35930 8111 35932
rect 7865 35878 7867 35930
rect 8047 35878 8049 35930
rect 7803 35876 7809 35878
rect 7865 35876 7889 35878
rect 7945 35876 7969 35878
rect 8025 35876 8049 35878
rect 8105 35876 8111 35878
rect 7803 35867 8111 35876
rect 7803 34844 8111 34853
rect 7803 34842 7809 34844
rect 7865 34842 7889 34844
rect 7945 34842 7969 34844
rect 8025 34842 8049 34844
rect 8105 34842 8111 34844
rect 7865 34790 7867 34842
rect 8047 34790 8049 34842
rect 7803 34788 7809 34790
rect 7865 34788 7889 34790
rect 7945 34788 7969 34790
rect 8025 34788 8049 34790
rect 8105 34788 8111 34790
rect 7803 34779 8111 34788
rect 7803 33756 8111 33765
rect 7803 33754 7809 33756
rect 7865 33754 7889 33756
rect 7945 33754 7969 33756
rect 8025 33754 8049 33756
rect 8105 33754 8111 33756
rect 7865 33702 7867 33754
rect 8047 33702 8049 33754
rect 7803 33700 7809 33702
rect 7865 33700 7889 33702
rect 7945 33700 7969 33702
rect 8025 33700 8049 33702
rect 8105 33700 8111 33702
rect 7803 33691 8111 33700
rect 7803 32668 8111 32677
rect 7803 32666 7809 32668
rect 7865 32666 7889 32668
rect 7945 32666 7969 32668
rect 8025 32666 8049 32668
rect 8105 32666 8111 32668
rect 7865 32614 7867 32666
rect 8047 32614 8049 32666
rect 7803 32612 7809 32614
rect 7865 32612 7889 32614
rect 7945 32612 7969 32614
rect 8025 32612 8049 32614
rect 8105 32612 8111 32614
rect 7803 32603 8111 32612
rect 7656 32428 7708 32434
rect 7656 32370 7708 32376
rect 7668 31754 7696 32370
rect 8220 32042 8248 39392
rect 8392 39374 8444 39380
rect 12716 39432 12768 39438
rect 12716 39374 12768 39380
rect 13360 39432 13412 39438
rect 13360 39374 13412 39380
rect 11230 39196 11538 39205
rect 11230 39194 11236 39196
rect 11292 39194 11316 39196
rect 11372 39194 11396 39196
rect 11452 39194 11476 39196
rect 11532 39194 11538 39196
rect 11292 39142 11294 39194
rect 11474 39142 11476 39194
rect 11230 39140 11236 39142
rect 11292 39140 11316 39142
rect 11372 39140 11396 39142
rect 11452 39140 11476 39142
rect 11532 39140 11538 39142
rect 11230 39131 11538 39140
rect 12728 39098 12756 39374
rect 12716 39092 12768 39098
rect 12716 39034 12768 39040
rect 12728 38962 12848 38978
rect 12624 38956 12676 38962
rect 12624 38898 12676 38904
rect 12728 38956 12860 38962
rect 12728 38950 12808 38956
rect 9517 38652 9825 38661
rect 9517 38650 9523 38652
rect 9579 38650 9603 38652
rect 9659 38650 9683 38652
rect 9739 38650 9763 38652
rect 9819 38650 9825 38652
rect 9579 38598 9581 38650
rect 9761 38598 9763 38650
rect 9517 38596 9523 38598
rect 9579 38596 9603 38598
rect 9659 38596 9683 38598
rect 9739 38596 9763 38598
rect 9819 38596 9825 38598
rect 9517 38587 9825 38596
rect 12440 38480 12492 38486
rect 12440 38422 12492 38428
rect 11612 38344 11664 38350
rect 11612 38286 11664 38292
rect 9404 38276 9456 38282
rect 9404 38218 9456 38224
rect 8300 36644 8352 36650
rect 8300 36586 8352 36592
rect 8312 34542 8340 36586
rect 9036 35012 9088 35018
rect 9036 34954 9088 34960
rect 9048 34678 9076 34954
rect 9036 34672 9088 34678
rect 9036 34614 9088 34620
rect 9220 34604 9272 34610
rect 9220 34546 9272 34552
rect 9312 34604 9364 34610
rect 9312 34546 9364 34552
rect 8300 34536 8352 34542
rect 8300 34478 8352 34484
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8128 32014 8248 32042
rect 8128 31822 8156 32014
rect 8208 31952 8260 31958
rect 8208 31894 8260 31900
rect 8116 31816 8168 31822
rect 8116 31758 8168 31764
rect 7472 31748 7524 31754
rect 7472 31690 7524 31696
rect 7576 31726 7696 31754
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7380 30048 7432 30054
rect 7380 29990 7432 29996
rect 7392 29850 7420 29990
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 7380 25696 7432 25702
rect 7380 25638 7432 25644
rect 7392 25498 7420 25638
rect 7380 25492 7432 25498
rect 7380 25434 7432 25440
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 7392 24818 7420 25162
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 7116 21678 7236 21706
rect 7286 21720 7342 21729
rect 7012 20936 7064 20942
rect 7012 20878 7064 20884
rect 7116 20602 7144 21678
rect 7286 21655 7342 21664
rect 7392 21622 7420 24754
rect 7196 21616 7248 21622
rect 7380 21616 7432 21622
rect 7196 21558 7248 21564
rect 7286 21584 7342 21593
rect 7104 20596 7156 20602
rect 7104 20538 7156 20544
rect 6748 19854 6776 20470
rect 6840 20454 6960 20482
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6840 20058 6868 20334
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6932 19700 6960 20454
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 7024 20058 7052 20266
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 7102 19952 7158 19961
rect 7102 19887 7158 19896
rect 7116 19854 7144 19887
rect 7104 19848 7156 19854
rect 7010 19816 7066 19825
rect 7104 19790 7156 19796
rect 7010 19751 7066 19760
rect 6748 19672 6960 19700
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6748 18358 6776 19672
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18766 6868 19246
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6736 18352 6788 18358
rect 6736 18294 6788 18300
rect 6840 17610 6868 18362
rect 6552 17604 6604 17610
rect 6552 17546 6604 17552
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6564 16794 6592 17546
rect 6552 16788 6604 16794
rect 6552 16730 6604 16736
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6368 13932 6420 13938
rect 6368 13874 6420 13880
rect 6090 13628 6398 13637
rect 6090 13626 6096 13628
rect 6152 13626 6176 13628
rect 6232 13626 6256 13628
rect 6312 13626 6336 13628
rect 6392 13626 6398 13628
rect 6152 13574 6154 13626
rect 6334 13574 6336 13626
rect 6090 13572 6096 13574
rect 6152 13572 6176 13574
rect 6232 13572 6256 13574
rect 6312 13572 6336 13574
rect 6392 13572 6398 13574
rect 6090 13563 6398 13572
rect 6092 13320 6144 13326
rect 6460 13320 6512 13326
rect 6144 13280 6460 13308
rect 6092 13262 6144 13268
rect 6460 13262 6512 13268
rect 6090 12540 6398 12549
rect 6090 12538 6096 12540
rect 6152 12538 6176 12540
rect 6232 12538 6256 12540
rect 6312 12538 6336 12540
rect 6392 12538 6398 12540
rect 6152 12486 6154 12538
rect 6334 12486 6336 12538
rect 6090 12484 6096 12486
rect 6152 12484 6176 12486
rect 6232 12484 6256 12486
rect 6312 12484 6336 12486
rect 6392 12484 6398 12486
rect 6090 12475 6398 12484
rect 6090 11452 6398 11461
rect 6090 11450 6096 11452
rect 6152 11450 6176 11452
rect 6232 11450 6256 11452
rect 6312 11450 6336 11452
rect 6392 11450 6398 11452
rect 6152 11398 6154 11450
rect 6334 11398 6336 11450
rect 6090 11396 6096 11398
rect 6152 11396 6176 11398
rect 6232 11396 6256 11398
rect 6312 11396 6336 11398
rect 6392 11396 6398 11398
rect 6090 11387 6398 11396
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 10470 6408 10542
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6090 10364 6398 10373
rect 6090 10362 6096 10364
rect 6152 10362 6176 10364
rect 6232 10362 6256 10364
rect 6312 10362 6336 10364
rect 6392 10362 6398 10364
rect 6152 10310 6154 10362
rect 6334 10310 6336 10362
rect 6090 10308 6096 10310
rect 6152 10308 6176 10310
rect 6232 10308 6256 10310
rect 6312 10308 6336 10310
rect 6392 10308 6398 10310
rect 6090 10299 6398 10308
rect 6012 10220 6132 10248
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 6104 9466 6132 10220
rect 6012 9438 6132 9466
rect 6012 7546 6040 9438
rect 6090 9276 6398 9285
rect 6090 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6336 9276
rect 6392 9274 6398 9276
rect 6152 9222 6154 9274
rect 6334 9222 6336 9274
rect 6090 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6336 9222
rect 6392 9220 6398 9222
rect 6090 9211 6398 9220
rect 6472 8634 6500 11154
rect 6564 10062 6592 16526
rect 6656 15008 6684 17546
rect 6932 15502 6960 19450
rect 7024 18272 7052 19751
rect 7116 19718 7144 19790
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7024 18244 7144 18272
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7024 17542 7052 18090
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6656 14980 6868 15008
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 10656 6684 13874
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12986 6776 13194
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6840 12434 6868 14980
rect 7024 12832 7052 17478
rect 7116 16580 7144 18244
rect 7104 16574 7156 16580
rect 7104 16516 7156 16522
rect 7104 16448 7156 16454
rect 7208 16436 7236 21558
rect 7380 21558 7432 21564
rect 7286 21519 7342 21528
rect 7298 21508 7328 21519
rect 7300 20466 7328 21508
rect 7484 21434 7512 31690
rect 7576 31142 7604 31726
rect 7803 31580 8111 31589
rect 7803 31578 7809 31580
rect 7865 31578 7889 31580
rect 7945 31578 7969 31580
rect 8025 31578 8049 31580
rect 8105 31578 8111 31580
rect 7865 31526 7867 31578
rect 8047 31526 8049 31578
rect 7803 31524 7809 31526
rect 7865 31524 7889 31526
rect 7945 31524 7969 31526
rect 8025 31524 8049 31526
rect 8105 31524 8111 31526
rect 7803 31515 8111 31524
rect 7564 31136 7616 31142
rect 7564 31078 7616 31084
rect 7576 28082 7604 31078
rect 7803 30492 8111 30501
rect 7803 30490 7809 30492
rect 7865 30490 7889 30492
rect 7945 30490 7969 30492
rect 8025 30490 8049 30492
rect 8105 30490 8111 30492
rect 7865 30438 7867 30490
rect 8047 30438 8049 30490
rect 7803 30436 7809 30438
rect 7865 30436 7889 30438
rect 7945 30436 7969 30438
rect 8025 30436 8049 30438
rect 8105 30436 8111 30438
rect 7803 30427 8111 30436
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7668 28994 7696 29650
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 8116 29640 8168 29646
rect 8220 29628 8248 31894
rect 8312 31346 8340 33458
rect 9140 32502 9168 33934
rect 8392 32496 8444 32502
rect 8392 32438 8444 32444
rect 9128 32496 9180 32502
rect 9128 32438 9180 32444
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8300 31136 8352 31142
rect 8300 31078 8352 31084
rect 8312 29850 8340 31078
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 8168 29600 8248 29628
rect 8116 29582 8168 29588
rect 7852 29492 7880 29582
rect 7852 29464 8248 29492
rect 7803 29404 8111 29413
rect 7803 29402 7809 29404
rect 7865 29402 7889 29404
rect 7945 29402 7969 29404
rect 8025 29402 8049 29404
rect 8105 29402 8111 29404
rect 7865 29350 7867 29402
rect 8047 29350 8049 29402
rect 7803 29348 7809 29350
rect 7865 29348 7889 29350
rect 7945 29348 7969 29350
rect 8025 29348 8049 29350
rect 8105 29348 8111 29350
rect 7803 29339 8111 29348
rect 8220 29288 8248 29464
rect 8300 29300 8352 29306
rect 8220 29260 8300 29288
rect 8300 29242 8352 29248
rect 7840 29164 7892 29170
rect 7840 29106 7892 29112
rect 8024 29164 8076 29170
rect 8024 29106 8076 29112
rect 7852 28994 7880 29106
rect 7668 28966 7880 28994
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7668 27112 7696 28966
rect 8036 28762 8064 29106
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 7803 28316 8111 28325
rect 7803 28314 7809 28316
rect 7865 28314 7889 28316
rect 7945 28314 7969 28316
rect 8025 28314 8049 28316
rect 8105 28314 8111 28316
rect 7865 28262 7867 28314
rect 8047 28262 8049 28314
rect 7803 28260 7809 28262
rect 7865 28260 7889 28262
rect 7945 28260 7969 28262
rect 8025 28260 8049 28262
rect 8105 28260 8111 28262
rect 7803 28251 8111 28260
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8220 27470 8248 28018
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 7803 27228 8111 27237
rect 7803 27226 7809 27228
rect 7865 27226 7889 27228
rect 7945 27226 7969 27228
rect 8025 27226 8049 27228
rect 8105 27226 8111 27228
rect 7865 27174 7867 27226
rect 8047 27174 8049 27226
rect 7803 27172 7809 27174
rect 7865 27172 7889 27174
rect 7945 27172 7969 27174
rect 8025 27172 8049 27174
rect 8105 27172 8111 27174
rect 7803 27163 8111 27172
rect 7668 27084 7788 27112
rect 7760 26926 7788 27084
rect 7564 26920 7616 26926
rect 7564 26862 7616 26868
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 7576 26518 7604 26862
rect 7760 26790 7788 26862
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7748 26784 7800 26790
rect 7748 26726 7800 26732
rect 7564 26512 7616 26518
rect 7564 26454 7616 26460
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7576 24886 7604 26250
rect 7564 24880 7616 24886
rect 7564 24822 7616 24828
rect 7564 24744 7616 24750
rect 7564 24686 7616 24692
rect 7576 22642 7604 24686
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7392 21418 7512 21434
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7380 21412 7512 21418
rect 7432 21406 7512 21412
rect 7380 21354 7432 21360
rect 7392 20942 7420 21354
rect 7576 21298 7604 21422
rect 7484 21270 7604 21298
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7484 20806 7512 21270
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 20369 7328 20402
rect 7286 20360 7342 20369
rect 7286 20295 7342 20304
rect 7392 19258 7420 20538
rect 7156 16408 7236 16436
rect 7300 19230 7420 19258
rect 7104 16390 7156 16396
rect 7116 16182 7144 16390
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 7194 16144 7250 16153
rect 7300 16114 7328 19230
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7392 18630 7420 18702
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7380 18216 7432 18222
rect 7380 18158 7432 18164
rect 7194 16079 7250 16088
rect 7288 16108 7340 16114
rect 7208 16028 7236 16079
rect 7288 16050 7340 16056
rect 7116 16000 7236 16028
rect 7116 13938 7144 16000
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 14958 7236 15302
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7116 12986 7144 13126
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7022 12804 7052 12832
rect 7102 12880 7158 12889
rect 7102 12815 7158 12824
rect 7022 12764 7050 12804
rect 7022 12736 7052 12764
rect 7024 12646 7052 12736
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 6748 12406 6868 12434
rect 6748 12238 6776 12406
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6748 11626 6776 12174
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6828 10668 6880 10674
rect 6656 10628 6828 10656
rect 6828 10610 6880 10616
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6564 8634 6592 9386
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6090 8188 6398 8197
rect 6090 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6336 8188
rect 6392 8186 6398 8188
rect 6152 8134 6154 8186
rect 6334 8134 6336 8186
rect 6090 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6336 8134
rect 6392 8132 6398 8134
rect 6090 8123 6398 8132
rect 6748 8090 6776 8434
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6550 7783 6606 7792
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6090 7100 6398 7109
rect 6090 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6336 7100
rect 6392 7098 6398 7100
rect 6152 7046 6154 7098
rect 6334 7046 6336 7098
rect 6090 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6336 7046
rect 6392 7044 6398 7046
rect 6090 7035 6398 7044
rect 6090 6012 6398 6021
rect 6090 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6336 6012
rect 6392 6010 6398 6012
rect 6152 5958 6154 6010
rect 6334 5958 6336 6010
rect 6090 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6336 5958
rect 6392 5956 6398 5958
rect 6090 5947 6398 5956
rect 6748 5710 6776 7686
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6840 7410 6868 7482
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 7002 6868 7346
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6932 6798 6960 11698
rect 7024 7993 7052 12174
rect 7010 7984 7066 7993
rect 7010 7919 7012 7928
rect 7064 7919 7066 7928
rect 7012 7890 7064 7896
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6322 6960 6734
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 4376 5468 4684 5477
rect 4376 5466 4382 5468
rect 4438 5466 4462 5468
rect 4518 5466 4542 5468
rect 4598 5466 4622 5468
rect 4678 5466 4684 5468
rect 4438 5414 4440 5466
rect 4620 5414 4622 5466
rect 4376 5412 4382 5414
rect 4438 5412 4462 5414
rect 4518 5412 4542 5414
rect 4598 5412 4622 5414
rect 4678 5412 4684 5414
rect 4376 5403 4684 5412
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 6090 4924 6398 4933
rect 6090 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6336 4924
rect 6392 4922 6398 4924
rect 6152 4870 6154 4922
rect 6334 4870 6336 4922
rect 6090 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6336 4870
rect 6392 4868 6398 4870
rect 6090 4859 6398 4868
rect 4376 4380 4684 4389
rect 4376 4378 4382 4380
rect 4438 4378 4462 4380
rect 4518 4378 4542 4380
rect 4598 4378 4622 4380
rect 4678 4378 4684 4380
rect 4438 4326 4440 4378
rect 4620 4326 4622 4378
rect 4376 4324 4382 4326
rect 4438 4324 4462 4326
rect 4518 4324 4542 4326
rect 4598 4324 4622 4326
rect 4678 4324 4684 4326
rect 4376 4315 4684 4324
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 6090 3836 6398 3845
rect 6090 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6336 3836
rect 6392 3834 6398 3836
rect 6152 3782 6154 3834
rect 6334 3782 6336 3834
rect 6090 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6336 3782
rect 6392 3780 6398 3782
rect 6090 3771 6398 3780
rect 4376 3292 4684 3301
rect 4376 3290 4382 3292
rect 4438 3290 4462 3292
rect 4518 3290 4542 3292
rect 4598 3290 4622 3292
rect 4678 3290 4684 3292
rect 4438 3238 4440 3290
rect 4620 3238 4622 3290
rect 4376 3236 4382 3238
rect 4438 3236 4462 3238
rect 4518 3236 4542 3238
rect 4598 3236 4622 3238
rect 4678 3236 4684 3238
rect 4376 3227 4684 3236
rect 7116 2774 7144 12815
rect 7208 8616 7236 14282
rect 7300 11830 7328 15438
rect 7392 12374 7420 18158
rect 7484 14906 7512 20742
rect 7564 20256 7616 20262
rect 7564 20198 7616 20204
rect 7576 18970 7604 20198
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7668 18850 7696 26726
rect 7852 26586 7880 26862
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 7803 26140 8111 26149
rect 7803 26138 7809 26140
rect 7865 26138 7889 26140
rect 7945 26138 7969 26140
rect 8025 26138 8049 26140
rect 8105 26138 8111 26140
rect 7865 26086 7867 26138
rect 8047 26086 8049 26138
rect 7803 26084 7809 26086
rect 7865 26084 7889 26086
rect 7945 26084 7969 26086
rect 8025 26084 8049 26086
rect 8105 26084 8111 26086
rect 7803 26075 8111 26084
rect 8220 26042 8248 27406
rect 8312 27130 8340 29242
rect 8404 27878 8432 32438
rect 9036 32224 9088 32230
rect 8956 32184 9036 32212
rect 8758 31240 8814 31249
rect 8758 31175 8814 31184
rect 8484 30320 8536 30326
rect 8484 30262 8536 30268
rect 8392 27872 8444 27878
rect 8392 27814 8444 27820
rect 8300 27124 8352 27130
rect 8300 27066 8352 27072
rect 8496 26246 8524 30262
rect 8772 29782 8800 31175
rect 8956 29782 8984 32184
rect 9232 32212 9260 34546
rect 9324 34202 9352 34546
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9416 34082 9444 38218
rect 11230 38108 11538 38117
rect 11230 38106 11236 38108
rect 11292 38106 11316 38108
rect 11372 38106 11396 38108
rect 11452 38106 11476 38108
rect 11532 38106 11538 38108
rect 11292 38054 11294 38106
rect 11474 38054 11476 38106
rect 11230 38052 11236 38054
rect 11292 38052 11316 38054
rect 11372 38052 11396 38054
rect 11452 38052 11476 38054
rect 11532 38052 11538 38054
rect 11230 38043 11538 38052
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 9517 37564 9825 37573
rect 9517 37562 9523 37564
rect 9579 37562 9603 37564
rect 9659 37562 9683 37564
rect 9739 37562 9763 37564
rect 9819 37562 9825 37564
rect 9579 37510 9581 37562
rect 9761 37510 9763 37562
rect 9517 37508 9523 37510
rect 9579 37508 9603 37510
rect 9659 37508 9683 37510
rect 9739 37508 9763 37510
rect 9819 37508 9825 37510
rect 9517 37499 9825 37508
rect 10796 37466 10824 37810
rect 10784 37460 10836 37466
rect 10784 37402 10836 37408
rect 10968 37256 11020 37262
rect 10968 37198 11020 37204
rect 10980 36922 11008 37198
rect 11230 37020 11538 37029
rect 11230 37018 11236 37020
rect 11292 37018 11316 37020
rect 11372 37018 11396 37020
rect 11452 37018 11476 37020
rect 11532 37018 11538 37020
rect 11292 36966 11294 37018
rect 11474 36966 11476 37018
rect 11230 36964 11236 36966
rect 11292 36964 11316 36966
rect 11372 36964 11396 36966
rect 11452 36964 11476 36966
rect 11532 36964 11538 36966
rect 11230 36955 11538 36964
rect 11624 36922 11652 38286
rect 11794 38176 11850 38185
rect 11794 38111 11850 38120
rect 11808 38010 11836 38111
rect 11796 38004 11848 38010
rect 11796 37946 11848 37952
rect 12452 37942 12480 38422
rect 12636 38298 12664 38898
rect 12728 38486 12756 38950
rect 12808 38898 12860 38904
rect 13268 38752 13320 38758
rect 13268 38694 13320 38700
rect 12944 38652 13252 38661
rect 12944 38650 12950 38652
rect 13006 38650 13030 38652
rect 13086 38650 13110 38652
rect 13166 38650 13190 38652
rect 13246 38650 13252 38652
rect 13006 38598 13008 38650
rect 13188 38598 13190 38650
rect 12944 38596 12950 38598
rect 13006 38596 13030 38598
rect 13086 38596 13110 38598
rect 13166 38596 13190 38598
rect 13246 38596 13252 38598
rect 12944 38587 13252 38596
rect 12716 38480 12768 38486
rect 12716 38422 12768 38428
rect 13280 38350 13308 38694
rect 13372 38554 13400 39374
rect 13912 39364 13964 39370
rect 13912 39306 13964 39312
rect 13924 39001 13952 39306
rect 14372 39296 14424 39302
rect 14372 39238 14424 39244
rect 13910 38992 13966 39001
rect 13452 38956 13504 38962
rect 13910 38927 13966 38936
rect 13452 38898 13504 38904
rect 13360 38548 13412 38554
rect 13360 38490 13412 38496
rect 12544 38270 12664 38298
rect 13176 38344 13228 38350
rect 13176 38286 13228 38292
rect 13268 38344 13320 38350
rect 13268 38286 13320 38292
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 12544 38010 12572 38270
rect 12624 38208 12676 38214
rect 12624 38150 12676 38156
rect 12532 38004 12584 38010
rect 12532 37946 12584 37952
rect 12440 37936 12492 37942
rect 12440 37878 12492 37884
rect 12072 37868 12124 37874
rect 12072 37810 12124 37816
rect 12532 37868 12584 37874
rect 12532 37810 12584 37816
rect 12084 37466 12112 37810
rect 12348 37732 12400 37738
rect 12348 37674 12400 37680
rect 12360 37466 12388 37674
rect 12072 37460 12124 37466
rect 12072 37402 12124 37408
rect 12348 37460 12400 37466
rect 12348 37402 12400 37408
rect 12544 37312 12572 37810
rect 12636 37670 12664 38150
rect 13188 38010 13216 38286
rect 13268 38208 13320 38214
rect 13268 38150 13320 38156
rect 13176 38004 13228 38010
rect 13176 37946 13228 37952
rect 13280 37874 13308 38150
rect 13084 37868 13136 37874
rect 12728 37828 13084 37856
rect 12624 37664 12676 37670
rect 12624 37606 12676 37612
rect 12624 37324 12676 37330
rect 12544 37284 12624 37312
rect 12624 37266 12676 37272
rect 11888 37256 11940 37262
rect 12728 37210 12756 37828
rect 13084 37810 13136 37816
rect 13268 37868 13320 37874
rect 13268 37810 13320 37816
rect 12944 37564 13252 37573
rect 12944 37562 12950 37564
rect 13006 37562 13030 37564
rect 13086 37562 13110 37564
rect 13166 37562 13190 37564
rect 13246 37562 13252 37564
rect 13006 37510 13008 37562
rect 13188 37510 13190 37562
rect 12944 37508 12950 37510
rect 13006 37508 13030 37510
rect 13086 37508 13110 37510
rect 13166 37508 13190 37510
rect 13246 37508 13252 37510
rect 12944 37499 13252 37508
rect 12808 37256 12860 37262
rect 11888 37198 11940 37204
rect 11900 36922 11928 37198
rect 12164 37188 12216 37194
rect 12164 37130 12216 37136
rect 12360 37182 12756 37210
rect 12806 37224 12808 37233
rect 12900 37256 12952 37262
rect 12860 37224 12862 37233
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 11612 36916 11664 36922
rect 11612 36858 11664 36864
rect 11888 36916 11940 36922
rect 11888 36858 11940 36864
rect 11888 36712 11940 36718
rect 11334 36680 11390 36689
rect 11334 36615 11336 36624
rect 11388 36615 11390 36624
rect 11808 36672 11888 36700
rect 11336 36586 11388 36592
rect 9517 36476 9825 36485
rect 9517 36474 9523 36476
rect 9579 36474 9603 36476
rect 9659 36474 9683 36476
rect 9739 36474 9763 36476
rect 9819 36474 9825 36476
rect 9579 36422 9581 36474
rect 9761 36422 9763 36474
rect 9517 36420 9523 36422
rect 9579 36420 9603 36422
rect 9659 36420 9683 36422
rect 9739 36420 9763 36422
rect 9819 36420 9825 36422
rect 9517 36411 9825 36420
rect 10968 36100 11020 36106
rect 10968 36042 11020 36048
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10692 35692 10744 35698
rect 10692 35634 10744 35640
rect 9517 35388 9825 35397
rect 9517 35386 9523 35388
rect 9579 35386 9603 35388
rect 9659 35386 9683 35388
rect 9739 35386 9763 35388
rect 9819 35386 9825 35388
rect 9579 35334 9581 35386
rect 9761 35334 9763 35386
rect 9517 35332 9523 35334
rect 9579 35332 9603 35334
rect 9659 35332 9683 35334
rect 9739 35332 9763 35334
rect 9819 35332 9825 35334
rect 9517 35323 9825 35332
rect 10428 35290 10456 35634
rect 10704 35290 10732 35634
rect 10980 35562 11008 36042
rect 11230 35932 11538 35941
rect 11230 35930 11236 35932
rect 11292 35930 11316 35932
rect 11372 35930 11396 35932
rect 11452 35930 11476 35932
rect 11532 35930 11538 35932
rect 11292 35878 11294 35930
rect 11474 35878 11476 35930
rect 11230 35876 11236 35878
rect 11292 35876 11316 35878
rect 11372 35876 11396 35878
rect 11452 35876 11476 35878
rect 11532 35876 11538 35878
rect 11230 35867 11538 35876
rect 11520 35624 11572 35630
rect 11572 35584 11652 35612
rect 11520 35566 11572 35572
rect 10968 35556 11020 35562
rect 10968 35498 11020 35504
rect 11152 35488 11204 35494
rect 11152 35430 11204 35436
rect 10416 35284 10468 35290
rect 10416 35226 10468 35232
rect 10692 35284 10744 35290
rect 10692 35226 10744 35232
rect 9680 35080 9732 35086
rect 11060 35080 11112 35086
rect 9680 35022 9732 35028
rect 10966 35048 11022 35057
rect 9692 34746 9720 35022
rect 11060 35022 11112 35028
rect 10966 34983 11022 34992
rect 10980 34746 11008 34983
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 9517 34300 9825 34309
rect 9517 34298 9523 34300
rect 9579 34298 9603 34300
rect 9659 34298 9683 34300
rect 9739 34298 9763 34300
rect 9819 34298 9825 34300
rect 9579 34246 9581 34298
rect 9761 34246 9763 34298
rect 9517 34244 9523 34246
rect 9579 34244 9603 34246
rect 9659 34244 9683 34246
rect 9739 34244 9763 34246
rect 9819 34244 9825 34246
rect 9517 34235 9825 34244
rect 9968 34202 9996 34546
rect 10140 34468 10192 34474
rect 10140 34410 10192 34416
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9036 32166 9088 32172
rect 9140 32184 9260 32212
rect 9324 34054 9444 34082
rect 9140 30394 9168 32184
rect 9220 31816 9272 31822
rect 9220 31758 9272 31764
rect 9232 31414 9260 31758
rect 9324 31754 9352 34054
rect 9404 33992 9456 33998
rect 9404 33934 9456 33940
rect 9588 33992 9640 33998
rect 9588 33934 9640 33940
rect 9416 33658 9444 33934
rect 9600 33658 9628 33934
rect 9864 33924 9916 33930
rect 9864 33866 9916 33872
rect 9876 33658 9904 33866
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 9588 33652 9640 33658
rect 9588 33594 9640 33600
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9517 33212 9825 33221
rect 9517 33210 9523 33212
rect 9579 33210 9603 33212
rect 9659 33210 9683 33212
rect 9739 33210 9763 33212
rect 9819 33210 9825 33212
rect 9579 33158 9581 33210
rect 9761 33158 9763 33210
rect 9517 33156 9523 33158
rect 9579 33156 9603 33158
rect 9659 33156 9683 33158
rect 9739 33156 9763 33158
rect 9819 33156 9825 33158
rect 9517 33147 9825 33156
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9517 32124 9825 32133
rect 9517 32122 9523 32124
rect 9579 32122 9603 32124
rect 9659 32122 9683 32124
rect 9739 32122 9763 32124
rect 9819 32122 9825 32124
rect 9579 32070 9581 32122
rect 9761 32070 9763 32122
rect 9517 32068 9523 32070
rect 9579 32068 9603 32070
rect 9659 32068 9683 32070
rect 9739 32068 9763 32070
rect 9819 32068 9825 32070
rect 9517 32059 9825 32068
rect 9324 31726 9444 31754
rect 9220 31408 9272 31414
rect 9220 31350 9272 31356
rect 9128 30388 9180 30394
rect 9128 30330 9180 30336
rect 9232 30240 9260 31350
rect 9140 30212 9260 30240
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 8760 29776 8812 29782
rect 8760 29718 8812 29724
rect 8944 29776 8996 29782
rect 8944 29718 8996 29724
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8760 29096 8812 29102
rect 8956 29073 8984 29582
rect 9048 29170 9076 30126
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 8760 29038 8812 29044
rect 8942 29064 8998 29073
rect 8668 29028 8720 29034
rect 8668 28970 8720 28976
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8588 26314 8616 27270
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 7803 25052 8111 25061
rect 7803 25050 7809 25052
rect 7865 25050 7889 25052
rect 7945 25050 7969 25052
rect 8025 25050 8049 25052
rect 8105 25050 8111 25052
rect 7865 24998 7867 25050
rect 8047 24998 8049 25050
rect 7803 24996 7809 24998
rect 7865 24996 7889 24998
rect 7945 24996 7969 24998
rect 8025 24996 8049 24998
rect 8105 24996 8111 24998
rect 7803 24987 8111 24996
rect 7803 23964 8111 23973
rect 7803 23962 7809 23964
rect 7865 23962 7889 23964
rect 7945 23962 7969 23964
rect 8025 23962 8049 23964
rect 8105 23962 8111 23964
rect 7865 23910 7867 23962
rect 8047 23910 8049 23962
rect 7803 23908 7809 23910
rect 7865 23908 7889 23910
rect 7945 23908 7969 23910
rect 8025 23908 8049 23910
rect 8105 23908 8111 23910
rect 7803 23899 8111 23908
rect 8116 23792 8168 23798
rect 8116 23734 8168 23740
rect 8128 22982 8156 23734
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8116 22976 8168 22982
rect 8116 22918 8168 22924
rect 7803 22876 8111 22885
rect 7803 22874 7809 22876
rect 7865 22874 7889 22876
rect 7945 22874 7969 22876
rect 8025 22874 8049 22876
rect 8105 22874 8111 22876
rect 7865 22822 7867 22874
rect 8047 22822 8049 22874
rect 7803 22820 7809 22822
rect 7865 22820 7889 22822
rect 7945 22820 7969 22822
rect 8025 22820 8049 22822
rect 8105 22820 8111 22822
rect 7803 22811 8111 22820
rect 8220 22574 8248 23462
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 7803 21788 8111 21797
rect 7803 21786 7809 21788
rect 7865 21786 7889 21788
rect 7945 21786 7969 21788
rect 8025 21786 8049 21788
rect 8105 21786 8111 21788
rect 7865 21734 7867 21786
rect 8047 21734 8049 21786
rect 7803 21732 7809 21734
rect 7865 21732 7889 21734
rect 7945 21732 7969 21734
rect 8025 21732 8049 21734
rect 8105 21732 8111 21734
rect 7803 21723 8111 21732
rect 8220 21672 8248 21830
rect 8128 21644 8248 21672
rect 8128 21486 8156 21644
rect 8116 21480 8168 21486
rect 8116 21422 8168 21428
rect 7803 20700 8111 20709
rect 7803 20698 7809 20700
rect 7865 20698 7889 20700
rect 7945 20698 7969 20700
rect 8025 20698 8049 20700
rect 8105 20698 8111 20700
rect 7865 20646 7867 20698
rect 8047 20646 8049 20698
rect 7803 20644 7809 20646
rect 7865 20644 7889 20646
rect 7945 20644 7969 20646
rect 8025 20644 8049 20646
rect 8105 20644 8111 20646
rect 7803 20635 8111 20644
rect 8206 20632 8262 20641
rect 8206 20567 8262 20576
rect 8220 19825 8248 20567
rect 8206 19816 8262 19825
rect 8206 19751 8262 19760
rect 7803 19612 8111 19621
rect 7803 19610 7809 19612
rect 7865 19610 7889 19612
rect 7945 19610 7969 19612
rect 8025 19610 8049 19612
rect 8105 19610 8111 19612
rect 7865 19558 7867 19610
rect 8047 19558 8049 19610
rect 7803 19556 7809 19558
rect 7865 19556 7889 19558
rect 7945 19556 7969 19558
rect 8025 19556 8049 19558
rect 8105 19556 8111 19558
rect 7803 19547 8111 19556
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7576 18822 7696 18850
rect 7576 17338 7604 18822
rect 7656 18760 7708 18766
rect 7656 18702 7708 18708
rect 7668 18358 7696 18702
rect 7760 18630 7788 19246
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7803 18524 8111 18533
rect 7803 18522 7809 18524
rect 7865 18522 7889 18524
rect 7945 18522 7969 18524
rect 8025 18522 8049 18524
rect 8105 18522 8111 18524
rect 7865 18470 7867 18522
rect 8047 18470 8049 18522
rect 7803 18468 7809 18470
rect 7865 18468 7889 18470
rect 7945 18468 7969 18470
rect 8025 18468 8049 18470
rect 8105 18468 8111 18470
rect 7803 18459 8111 18468
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16046 7604 16934
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7484 14890 7604 14906
rect 7472 14884 7604 14890
rect 7524 14878 7604 14884
rect 7472 14826 7524 14832
rect 7472 14068 7524 14074
rect 7472 14010 7524 14016
rect 7484 13530 7512 14010
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 12986 7604 14878
rect 7668 14346 7696 18294
rect 8220 18222 8248 19110
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 7803 17436 8111 17445
rect 7803 17434 7809 17436
rect 7865 17434 7889 17436
rect 7945 17434 7969 17436
rect 8025 17434 8049 17436
rect 8105 17434 8111 17436
rect 7865 17382 7867 17434
rect 8047 17382 8049 17434
rect 7803 17380 7809 17382
rect 7865 17380 7889 17382
rect 7945 17380 7969 17382
rect 8025 17380 8049 17382
rect 8105 17380 8111 17382
rect 7803 17371 8111 17380
rect 8220 17377 8248 18022
rect 8206 17368 8262 17377
rect 7748 17332 7800 17338
rect 8206 17303 8262 17312
rect 7748 17274 7800 17280
rect 7760 16522 7788 17274
rect 8312 17066 8340 25842
rect 8680 25226 8708 28970
rect 8772 28694 8800 29038
rect 8942 28999 8998 29008
rect 8760 28688 8812 28694
rect 8760 28630 8812 28636
rect 8852 28552 8904 28558
rect 8852 28494 8904 28500
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8772 26353 8800 26862
rect 8864 26518 8892 28494
rect 9140 28370 9168 30212
rect 9312 30184 9364 30190
rect 9232 30132 9312 30138
rect 9232 30126 9364 30132
rect 9232 30110 9352 30126
rect 9232 29714 9260 30110
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 9232 29073 9260 29650
rect 9218 29064 9274 29073
rect 9218 28999 9274 29008
rect 9140 28342 9352 28370
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 9140 27010 9168 27814
rect 9140 26982 9260 27010
rect 9232 26926 9260 26982
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9036 26852 9088 26858
rect 9036 26794 9088 26800
rect 8944 26784 8996 26790
rect 8944 26726 8996 26732
rect 8852 26512 8904 26518
rect 8852 26454 8904 26460
rect 8758 26344 8814 26353
rect 8758 26279 8814 26288
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8496 23780 8524 24550
rect 8588 24018 8616 24686
rect 8760 24676 8812 24682
rect 8760 24618 8812 24624
rect 8772 24342 8800 24618
rect 8760 24336 8812 24342
rect 8680 24284 8760 24290
rect 8680 24278 8812 24284
rect 8680 24262 8800 24278
rect 8680 24138 8708 24262
rect 8864 24154 8892 26454
rect 8668 24132 8720 24138
rect 8668 24074 8720 24080
rect 8772 24126 8892 24154
rect 8588 23990 8708 24018
rect 8576 23792 8628 23798
rect 8496 23752 8576 23780
rect 8576 23734 8628 23740
rect 8484 23248 8536 23254
rect 8482 23216 8484 23225
rect 8536 23216 8538 23225
rect 8482 23151 8538 23160
rect 8482 23080 8538 23089
rect 8482 23015 8484 23024
rect 8536 23015 8538 23024
rect 8484 22986 8536 22992
rect 8588 22574 8616 23734
rect 8680 22574 8708 23990
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8668 22568 8720 22574
rect 8668 22510 8720 22516
rect 8772 22522 8800 24126
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 22642 8892 24006
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 8482 21856 8538 21865
rect 8482 21791 8538 21800
rect 8496 21690 8524 21791
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8484 21684 8536 21690
rect 8484 21626 8536 21632
rect 8404 21554 8432 21626
rect 8496 21554 8524 21626
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8484 21548 8536 21554
rect 8484 21490 8536 21496
rect 8404 19446 8432 21490
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8588 17898 8616 22510
rect 8680 22420 8708 22510
rect 8772 22494 8892 22522
rect 8680 22392 8800 22420
rect 8772 21706 8800 22392
rect 8864 21865 8892 22494
rect 8850 21856 8906 21865
rect 8850 21791 8906 21800
rect 8772 21678 8892 21706
rect 8668 21548 8720 21554
rect 8668 21490 8720 21496
rect 8680 21146 8708 21490
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8680 20602 8708 20810
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8404 17870 8616 17898
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16794 8340 17002
rect 8300 16788 8352 16794
rect 8300 16730 8352 16736
rect 7748 16516 7800 16522
rect 7748 16458 7800 16464
rect 7803 16348 8111 16357
rect 7803 16346 7809 16348
rect 7865 16346 7889 16348
rect 7945 16346 7969 16348
rect 8025 16346 8049 16348
rect 8105 16346 8111 16348
rect 7865 16294 7867 16346
rect 8047 16294 8049 16346
rect 7803 16292 7809 16294
rect 7865 16292 7889 16294
rect 7945 16292 7969 16294
rect 8025 16292 8049 16294
rect 8105 16292 8111 16294
rect 7803 16283 8111 16292
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7852 16130 7880 16186
rect 7760 16102 7880 16130
rect 8404 16114 8432 17870
rect 8680 17626 8708 19654
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8772 18426 8800 19382
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8772 18290 8800 18362
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8496 17598 8708 17626
rect 8392 16108 8444 16114
rect 7760 16046 7788 16102
rect 8392 16050 8444 16056
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7803 15260 8111 15269
rect 7803 15258 7809 15260
rect 7865 15258 7889 15260
rect 7945 15258 7969 15260
rect 8025 15258 8049 15260
rect 8105 15258 8111 15260
rect 7865 15206 7867 15258
rect 8047 15206 8049 15258
rect 7803 15204 7809 15206
rect 7865 15204 7889 15206
rect 7945 15204 7969 15206
rect 8025 15204 8049 15206
rect 8105 15204 8111 15206
rect 7803 15195 8111 15204
rect 7840 15020 7892 15026
rect 7840 14962 7892 14968
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 7852 14482 7880 14962
rect 8128 14618 8156 14962
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 8220 14385 8248 15982
rect 8404 15706 8432 16050
rect 8392 15700 8444 15706
rect 8392 15642 8444 15648
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8206 14376 8262 14385
rect 7656 14340 7708 14346
rect 8206 14311 8262 14320
rect 7656 14282 7708 14288
rect 7803 14172 8111 14181
rect 7803 14170 7809 14172
rect 7865 14170 7889 14172
rect 7945 14170 7969 14172
rect 8025 14170 8049 14172
rect 8105 14170 8111 14172
rect 7865 14118 7867 14170
rect 8047 14118 8049 14170
rect 7803 14116 7809 14118
rect 7865 14116 7889 14118
rect 7945 14116 7969 14118
rect 8025 14116 8049 14118
rect 8105 14116 8111 14118
rect 7803 14107 8111 14116
rect 8312 13977 8340 14554
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8298 13968 8354 13977
rect 8298 13903 8354 13912
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 8208 13864 8260 13870
rect 8300 13864 8352 13870
rect 8260 13824 8300 13852
rect 8208 13806 8260 13812
rect 8300 13806 8352 13812
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7668 12782 7696 13806
rect 8298 13696 8354 13705
rect 8298 13631 8354 13640
rect 7803 13084 8111 13093
rect 7803 13082 7809 13084
rect 7865 13082 7889 13084
rect 7945 13082 7969 13084
rect 8025 13082 8049 13084
rect 8105 13082 8111 13084
rect 7865 13030 7867 13082
rect 8047 13030 8049 13082
rect 7803 13028 7809 13030
rect 7865 13028 7889 13030
rect 7945 13028 7969 13030
rect 8025 13028 8049 13030
rect 8105 13028 8111 13030
rect 7803 13019 8111 13028
rect 7656 12776 7708 12782
rect 7654 12744 7656 12753
rect 7708 12744 7710 12753
rect 7472 12708 7524 12714
rect 7654 12679 7710 12688
rect 7472 12650 7524 12656
rect 7380 12368 7432 12374
rect 7380 12310 7432 12316
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 9518 7420 10406
rect 7484 10130 7512 12650
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7564 12300 7616 12306
rect 7564 12242 7616 12248
rect 7576 11354 7604 12242
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7668 10792 7696 12582
rect 7944 12306 7972 12582
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8116 12232 8168 12238
rect 8168 12192 8248 12220
rect 8116 12174 8168 12180
rect 7852 12102 7880 12174
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7803 11996 8111 12005
rect 7803 11994 7809 11996
rect 7865 11994 7889 11996
rect 7945 11994 7969 11996
rect 8025 11994 8049 11996
rect 8105 11994 8111 11996
rect 7865 11942 7867 11994
rect 8047 11942 8049 11994
rect 7803 11940 7809 11942
rect 7865 11940 7889 11942
rect 7945 11940 7969 11942
rect 8025 11940 8049 11942
rect 8105 11940 8111 11942
rect 7803 11931 8111 11940
rect 8220 11898 8248 12192
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7803 10908 8111 10917
rect 7803 10906 7809 10908
rect 7865 10906 7889 10908
rect 7945 10906 7969 10908
rect 8025 10906 8049 10908
rect 8105 10906 8111 10908
rect 7865 10854 7867 10906
rect 8047 10854 8049 10906
rect 7803 10852 7809 10854
rect 7865 10852 7889 10854
rect 7945 10852 7969 10854
rect 8025 10852 8049 10854
rect 8105 10852 8111 10854
rect 7803 10843 8111 10852
rect 7668 10764 7788 10792
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7472 10124 7524 10130
rect 7524 10084 7604 10112
rect 7472 10066 7524 10072
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9722 7512 9862
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9042 7328 9318
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7208 8588 7328 8616
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 8090 7236 8434
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7208 6254 7236 7414
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5778 7236 6190
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7208 5234 7236 5714
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7300 4554 7328 8588
rect 7484 8362 7512 8910
rect 7576 8498 7604 10084
rect 7668 9518 7696 10134
rect 7760 9908 7788 10764
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7852 10130 7880 10542
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7840 10124 7892 10130
rect 7840 10066 7892 10072
rect 8128 10062 8156 10406
rect 8312 10112 8340 13631
rect 8404 13530 8432 14350
rect 8496 14249 8524 17598
rect 8680 17338 8708 17598
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8864 17218 8892 21678
rect 8956 19718 8984 26726
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 9048 19258 9076 26794
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9232 24818 9260 25638
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9128 24744 9180 24750
rect 9128 24686 9180 24692
rect 9140 24614 9168 24686
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9232 24426 9260 24550
rect 9140 24398 9260 24426
rect 9140 23662 9168 24398
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9140 23322 9168 23598
rect 9128 23316 9180 23322
rect 9128 23258 9180 23264
rect 9128 23112 9180 23118
rect 9128 23054 9180 23060
rect 9140 20058 9168 23054
rect 9128 20052 9180 20058
rect 9128 19994 9180 20000
rect 9126 19680 9182 19689
rect 9126 19615 9182 19624
rect 9140 19378 9168 19615
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9048 19230 9168 19258
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9048 18766 9076 19110
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18272 8984 18566
rect 9036 18284 9088 18290
rect 8956 18244 9036 18272
rect 9036 18226 9088 18232
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 8588 17190 8892 17218
rect 9048 17202 9076 17478
rect 9036 17196 9088 17202
rect 8588 16114 8616 17190
rect 9036 17138 9088 17144
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8680 16114 8708 16662
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8588 15434 8616 16050
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8588 14618 8616 15098
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8482 14240 8538 14249
rect 8482 14175 8538 14184
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8496 12850 8524 14175
rect 8588 12850 8616 14282
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11898 8432 12038
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8588 11082 8616 12786
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10266 8524 10406
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8312 10084 8432 10112
rect 8116 10056 8168 10062
rect 8168 10004 8340 10010
rect 8116 9998 8340 10004
rect 8128 9982 8340 9998
rect 7742 9880 7788 9908
rect 7742 9704 7770 9880
rect 7803 9820 8111 9829
rect 7803 9818 7809 9820
rect 7865 9818 7889 9820
rect 7945 9818 7969 9820
rect 8025 9818 8049 9820
rect 8105 9818 8111 9820
rect 7865 9766 7867 9818
rect 8047 9766 8049 9818
rect 7803 9764 7809 9766
rect 7865 9764 7889 9766
rect 7945 9764 7969 9766
rect 8025 9764 8049 9766
rect 8105 9764 8111 9766
rect 7803 9755 8111 9764
rect 7742 9676 7788 9704
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7760 8820 7788 9676
rect 8312 9586 8340 9982
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7840 9444 7892 9450
rect 7840 9386 7892 9392
rect 7852 8906 7880 9386
rect 8036 8974 8064 9454
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 7668 8792 7788 8820
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7484 7954 7512 8298
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7546 7604 7890
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7668 5370 7696 8792
rect 7803 8732 8111 8741
rect 7803 8730 7809 8732
rect 7865 8730 7889 8732
rect 7945 8730 7969 8732
rect 8025 8730 8049 8732
rect 8105 8730 8111 8732
rect 7865 8678 7867 8730
rect 8047 8678 8049 8730
rect 7803 8676 7809 8678
rect 7865 8676 7889 8678
rect 7945 8676 7969 8678
rect 8025 8676 8049 8678
rect 8105 8676 8111 8678
rect 7803 8667 8111 8676
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7954 7972 8230
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7803 7644 8111 7653
rect 7803 7642 7809 7644
rect 7865 7642 7889 7644
rect 7945 7642 7969 7644
rect 8025 7642 8049 7644
rect 8105 7642 8111 7644
rect 7865 7590 7867 7642
rect 8047 7590 8049 7642
rect 7803 7588 7809 7590
rect 7865 7588 7889 7590
rect 7945 7588 7969 7590
rect 8025 7588 8049 7590
rect 8105 7588 8111 7590
rect 7803 7579 8111 7588
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8128 6934 8156 7278
rect 8220 7274 8248 9454
rect 8404 9042 8432 10084
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 8090 8616 8366
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7803 6556 8111 6565
rect 7803 6554 7809 6556
rect 7865 6554 7889 6556
rect 7945 6554 7969 6556
rect 8025 6554 8049 6556
rect 8105 6554 8111 6556
rect 7865 6502 7867 6554
rect 8047 6502 8049 6554
rect 7803 6500 7809 6502
rect 7865 6500 7889 6502
rect 7945 6500 7969 6502
rect 8025 6500 8049 6502
rect 8105 6500 8111 6502
rect 7803 6491 8111 6500
rect 8300 6384 8352 6390
rect 8298 6352 8300 6361
rect 8352 6352 8354 6361
rect 8298 6287 8354 6296
rect 8208 5704 8260 5710
rect 8206 5672 8208 5681
rect 8260 5672 8262 5681
rect 8206 5607 8262 5616
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7803 5468 8111 5477
rect 7803 5466 7809 5468
rect 7865 5466 7889 5468
rect 7945 5466 7969 5468
rect 8025 5466 8049 5468
rect 8105 5466 8111 5468
rect 7865 5414 7867 5466
rect 8047 5414 8049 5466
rect 7803 5412 7809 5414
rect 7865 5412 7889 5414
rect 7945 5412 7969 5414
rect 8025 5412 8049 5414
rect 8105 5412 8111 5414
rect 7803 5403 8111 5412
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 8312 5302 8340 5510
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4690 8340 4966
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7803 4380 8111 4389
rect 7803 4378 7809 4380
rect 7865 4378 7889 4380
rect 7945 4378 7969 4380
rect 8025 4378 8049 4380
rect 8105 4378 8111 4380
rect 7865 4326 7867 4378
rect 8047 4326 8049 4378
rect 7803 4324 7809 4326
rect 7865 4324 7889 4326
rect 7945 4324 7969 4326
rect 8025 4324 8049 4326
rect 8105 4324 8111 4326
rect 7803 4315 8111 4324
rect 8312 4078 8340 4626
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7803 3292 8111 3301
rect 7803 3290 7809 3292
rect 7865 3290 7889 3292
rect 7945 3290 7969 3292
rect 8025 3290 8049 3292
rect 8105 3290 8111 3292
rect 7865 3238 7867 3290
rect 8047 3238 8049 3290
rect 7803 3236 7809 3238
rect 7865 3236 7889 3238
rect 7945 3236 7969 3238
rect 8025 3236 8049 3238
rect 8105 3236 8111 3238
rect 7803 3227 8111 3236
rect 8312 2774 8340 4014
rect 6090 2748 6398 2757
rect 6090 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6336 2748
rect 6392 2746 6398 2748
rect 7116 2746 7236 2774
rect 8312 2746 8432 2774
rect 6152 2694 6154 2746
rect 6334 2694 6336 2746
rect 6090 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6336 2694
rect 6392 2692 6398 2694
rect 5814 2680 5870 2689
rect 6090 2683 6398 2692
rect 5814 2615 5870 2624
rect 6642 2680 6698 2689
rect 6642 2615 6698 2624
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 4080 2106 4108 2314
rect 4376 2204 4684 2213
rect 4376 2202 4382 2204
rect 4438 2202 4462 2204
rect 4518 2202 4542 2204
rect 4598 2202 4622 2204
rect 4678 2202 4684 2204
rect 4438 2150 4440 2202
rect 4620 2150 4622 2202
rect 4376 2148 4382 2150
rect 4438 2148 4462 2150
rect 4518 2148 4542 2150
rect 4598 2148 4622 2150
rect 4678 2148 4684 2150
rect 4376 2139 4684 2148
rect 5828 2106 5856 2615
rect 6656 2106 6684 2615
rect 7208 2106 7236 2746
rect 7654 2680 7710 2689
rect 7654 2615 7710 2624
rect 7668 2106 7696 2615
rect 7803 2204 8111 2213
rect 7803 2202 7809 2204
rect 7865 2202 7889 2204
rect 7945 2202 7969 2204
rect 8025 2202 8049 2204
rect 8105 2202 8111 2204
rect 7865 2150 7867 2202
rect 8047 2150 8049 2202
rect 7803 2148 7809 2150
rect 7865 2148 7889 2150
rect 7945 2148 7969 2150
rect 8025 2148 8049 2150
rect 8105 2148 8111 2150
rect 7803 2139 8111 2148
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 4252 1964 4304 1970
rect 4252 1906 4304 1912
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 3240 1828 3292 1834
rect 3240 1770 3292 1776
rect 2412 1760 2464 1766
rect 2412 1702 2464 1708
rect 2663 1660 2971 1669
rect 2663 1658 2669 1660
rect 2725 1658 2749 1660
rect 2805 1658 2829 1660
rect 2885 1658 2909 1660
rect 2965 1658 2971 1660
rect 2725 1606 2727 1658
rect 2907 1606 2909 1658
rect 2663 1604 2669 1606
rect 2725 1604 2749 1606
rect 2805 1604 2829 1606
rect 2885 1604 2909 1606
rect 2965 1604 2971 1606
rect 2663 1595 2971 1604
rect 4264 1562 4292 1906
rect 5000 1562 5028 1906
rect 5736 1562 5764 1906
rect 6090 1660 6398 1669
rect 6090 1658 6096 1660
rect 6152 1658 6176 1660
rect 6232 1658 6256 1660
rect 6312 1658 6336 1660
rect 6392 1658 6398 1660
rect 6152 1606 6154 1658
rect 6334 1606 6336 1658
rect 6090 1604 6096 1606
rect 6152 1604 6176 1606
rect 6232 1604 6256 1606
rect 6312 1604 6336 1606
rect 6392 1604 6398 1606
rect 6090 1595 6398 1604
rect 6472 1562 6500 1906
rect 7116 1562 7144 1906
rect 7852 1562 7880 1906
rect 4252 1556 4304 1562
rect 4252 1498 4304 1504
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 7104 1556 7156 1562
rect 7104 1498 7156 1504
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 2780 1352 2832 1358
rect 2780 1294 2832 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 2228 1284 2280 1290
rect 2228 1226 2280 1232
rect 2240 1018 2268 1226
rect 2228 1012 2280 1018
rect 2228 954 2280 960
rect 2792 160 2820 1294
rect 2042 54 2176 82
rect 2042 0 2098 54
rect 2778 0 2834 160
rect 3514 82 3570 160
rect 3804 82 3832 1294
rect 4264 160 4292 1294
rect 4376 1116 4684 1125
rect 4376 1114 4382 1116
rect 4438 1114 4462 1116
rect 4518 1114 4542 1116
rect 4598 1114 4622 1116
rect 4678 1114 4684 1116
rect 4438 1062 4440 1114
rect 4620 1062 4622 1114
rect 4376 1060 4382 1062
rect 4438 1060 4462 1062
rect 4518 1060 4542 1062
rect 4598 1060 4622 1062
rect 4678 1060 4684 1062
rect 4376 1051 4684 1060
rect 5000 160 5028 1294
rect 5736 160 5764 1294
rect 6472 160 6500 1294
rect 3514 54 3832 82
rect 3514 0 3570 54
rect 4250 0 4306 160
rect 4986 0 5042 160
rect 5722 0 5778 160
rect 6458 0 6514 160
rect 7194 82 7250 160
rect 7484 82 7512 1294
rect 7803 1116 8111 1125
rect 7803 1114 7809 1116
rect 7865 1114 7889 1116
rect 7945 1114 7969 1116
rect 8025 1114 8049 1116
rect 8105 1114 8111 1116
rect 7865 1062 7867 1114
rect 8047 1062 8049 1114
rect 7803 1060 7809 1062
rect 7865 1060 7889 1062
rect 7945 1060 7969 1062
rect 8025 1060 8049 1062
rect 8105 1060 8111 1062
rect 7803 1051 8111 1060
rect 7194 54 7512 82
rect 7930 82 7986 160
rect 8220 82 8248 1294
rect 8404 1018 8432 2746
rect 8680 2106 8708 14486
rect 8772 13530 8800 14758
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8772 12850 8800 13126
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8864 12434 8892 17070
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8956 14414 8984 15438
rect 9140 15008 9168 19230
rect 9232 17202 9260 24278
rect 9324 19854 9352 28342
rect 9416 24750 9444 31726
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9517 31036 9825 31045
rect 9517 31034 9523 31036
rect 9579 31034 9603 31036
rect 9659 31034 9683 31036
rect 9739 31034 9763 31036
rect 9819 31034 9825 31036
rect 9579 30982 9581 31034
rect 9761 30982 9763 31034
rect 9517 30980 9523 30982
rect 9579 30980 9603 30982
rect 9659 30980 9683 30982
rect 9739 30980 9763 30982
rect 9819 30980 9825 30982
rect 9517 30971 9825 30980
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9692 30122 9720 30670
rect 9876 30190 9904 31078
rect 9968 30682 9996 32846
rect 10048 32496 10100 32502
rect 10048 32438 10100 32444
rect 10060 31754 10088 32438
rect 10152 32026 10180 34410
rect 10796 34202 10824 34546
rect 10784 34196 10836 34202
rect 10784 34138 10836 34144
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10612 33114 10640 33458
rect 11072 33114 11100 35022
rect 11164 34746 11192 35430
rect 11230 34844 11538 34853
rect 11230 34842 11236 34844
rect 11292 34842 11316 34844
rect 11372 34842 11396 34844
rect 11452 34842 11476 34844
rect 11532 34842 11538 34844
rect 11292 34790 11294 34842
rect 11474 34790 11476 34842
rect 11230 34788 11236 34790
rect 11292 34788 11316 34790
rect 11372 34788 11396 34790
rect 11452 34788 11476 34790
rect 11532 34788 11538 34790
rect 11230 34779 11538 34788
rect 11152 34740 11204 34746
rect 11152 34682 11204 34688
rect 11624 34082 11652 35584
rect 11808 35154 11836 36672
rect 11888 36654 11940 36660
rect 12176 36378 12204 37130
rect 12360 36922 12388 37182
rect 12900 37198 12952 37204
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 12806 37159 12862 37168
rect 12716 37120 12768 37126
rect 12452 37080 12716 37108
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12452 36174 12480 37080
rect 12716 37062 12768 37068
rect 12716 36780 12768 36786
rect 12636 36740 12716 36768
rect 12532 36576 12584 36582
rect 12532 36518 12584 36524
rect 12544 36378 12572 36518
rect 12532 36372 12584 36378
rect 12532 36314 12584 36320
rect 12636 36310 12664 36740
rect 12716 36722 12768 36728
rect 12912 36666 12940 37198
rect 13176 37120 13228 37126
rect 13176 37062 13228 37068
rect 13188 36922 13216 37062
rect 13176 36916 13228 36922
rect 13176 36858 13228 36864
rect 12992 36780 13044 36786
rect 12992 36722 13044 36728
rect 13004 36689 13032 36722
rect 12820 36638 12940 36666
rect 12990 36680 13046 36689
rect 12716 36372 12768 36378
rect 12716 36314 12768 36320
rect 12624 36304 12676 36310
rect 12624 36246 12676 36252
rect 12728 36174 12756 36314
rect 12820 36174 12848 36638
rect 12990 36615 13046 36624
rect 12944 36476 13252 36485
rect 12944 36474 12950 36476
rect 13006 36474 13030 36476
rect 13086 36474 13110 36476
rect 13166 36474 13190 36476
rect 13246 36474 13252 36476
rect 13006 36422 13008 36474
rect 13188 36422 13190 36474
rect 12944 36420 12950 36422
rect 13006 36420 13030 36422
rect 13086 36420 13110 36422
rect 13166 36420 13190 36422
rect 13246 36420 13252 36422
rect 12944 36411 13252 36420
rect 12900 36304 12952 36310
rect 12900 36246 12952 36252
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 12624 36168 12676 36174
rect 12624 36110 12676 36116
rect 12716 36168 12768 36174
rect 12716 36110 12768 36116
rect 12808 36168 12860 36174
rect 12808 36110 12860 36116
rect 12636 35894 12664 36110
rect 11992 35866 12664 35894
rect 11992 35766 12020 35866
rect 11980 35760 12032 35766
rect 11980 35702 12032 35708
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11716 34202 11744 34886
rect 11900 34678 11928 35634
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11796 34604 11848 34610
rect 11796 34546 11848 34552
rect 11704 34196 11756 34202
rect 11704 34138 11756 34144
rect 11164 34054 11652 34082
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 11164 32994 11192 34054
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 11230 33756 11538 33765
rect 11230 33754 11236 33756
rect 11292 33754 11316 33756
rect 11372 33754 11396 33756
rect 11452 33754 11476 33756
rect 11532 33754 11538 33756
rect 11292 33702 11294 33754
rect 11474 33702 11476 33754
rect 11230 33700 11236 33702
rect 11292 33700 11316 33702
rect 11372 33700 11396 33702
rect 11452 33700 11476 33702
rect 11532 33700 11538 33702
rect 11230 33691 11538 33700
rect 11624 33538 11652 33934
rect 11704 33856 11756 33862
rect 11704 33798 11756 33804
rect 11532 33510 11652 33538
rect 11532 33454 11560 33510
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11426 33144 11482 33153
rect 11426 33079 11482 33088
rect 11440 33046 11468 33079
rect 11072 32966 11192 32994
rect 11428 33040 11480 33046
rect 11428 32982 11480 32988
rect 11072 32858 11100 32966
rect 10796 32830 11100 32858
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11532 32858 11560 33390
rect 10416 32224 10468 32230
rect 10416 32166 10468 32172
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10060 31726 10272 31754
rect 9968 30654 10180 30682
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9772 30184 9824 30190
rect 9772 30126 9824 30132
rect 9864 30184 9916 30190
rect 9864 30126 9916 30132
rect 9680 30116 9732 30122
rect 9680 30058 9732 30064
rect 9784 30036 9812 30126
rect 9784 30008 9904 30036
rect 9517 29948 9825 29957
rect 9517 29946 9523 29948
rect 9579 29946 9603 29948
rect 9659 29946 9683 29948
rect 9739 29946 9763 29948
rect 9819 29946 9825 29948
rect 9579 29894 9581 29946
rect 9761 29894 9763 29946
rect 9517 29892 9523 29894
rect 9579 29892 9603 29894
rect 9659 29892 9683 29894
rect 9739 29892 9763 29894
rect 9819 29892 9825 29894
rect 9517 29883 9825 29892
rect 9876 29646 9904 30008
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9876 29306 9904 29582
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9517 28860 9825 28869
rect 9517 28858 9523 28860
rect 9579 28858 9603 28860
rect 9659 28858 9683 28860
rect 9739 28858 9763 28860
rect 9819 28858 9825 28860
rect 9579 28806 9581 28858
rect 9761 28806 9763 28858
rect 9517 28804 9523 28806
rect 9579 28804 9603 28806
rect 9659 28804 9683 28806
rect 9739 28804 9763 28806
rect 9819 28804 9825 28806
rect 9517 28795 9825 28804
rect 9680 28620 9732 28626
rect 9732 28580 9812 28608
rect 9680 28562 9732 28568
rect 9784 28150 9812 28580
rect 9772 28144 9824 28150
rect 9772 28086 9824 28092
rect 9864 28076 9916 28082
rect 9968 28064 9996 30534
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10060 29510 10088 29582
rect 10048 29504 10100 29510
rect 10048 29446 10100 29452
rect 10152 29322 10180 30654
rect 9916 28036 9996 28064
rect 10060 29294 10180 29322
rect 9864 28018 9916 28024
rect 9517 27772 9825 27781
rect 9517 27770 9523 27772
rect 9579 27770 9603 27772
rect 9659 27770 9683 27772
rect 9739 27770 9763 27772
rect 9819 27770 9825 27772
rect 9579 27718 9581 27770
rect 9761 27718 9763 27770
rect 9517 27716 9523 27718
rect 9579 27716 9603 27718
rect 9659 27716 9683 27718
rect 9739 27716 9763 27718
rect 9819 27716 9825 27718
rect 9517 27707 9825 27716
rect 9680 27396 9732 27402
rect 9680 27338 9732 27344
rect 9692 27130 9720 27338
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9784 26994 9812 27270
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9600 26790 9628 26862
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9517 26684 9825 26693
rect 9517 26682 9523 26684
rect 9579 26682 9603 26684
rect 9659 26682 9683 26684
rect 9739 26682 9763 26684
rect 9819 26682 9825 26684
rect 9579 26630 9581 26682
rect 9761 26630 9763 26682
rect 9517 26628 9523 26630
rect 9579 26628 9603 26630
rect 9659 26628 9683 26630
rect 9739 26628 9763 26630
rect 9819 26628 9825 26630
rect 9517 26619 9825 26628
rect 9876 25974 9904 28018
rect 10060 27878 10088 29294
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10152 28694 10180 28902
rect 10140 28688 10192 28694
rect 10140 28630 10192 28636
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10048 27872 10100 27878
rect 10048 27814 10100 27820
rect 9956 26580 10008 26586
rect 9956 26522 10008 26528
rect 9968 26042 9996 26522
rect 10060 26382 10088 27814
rect 10048 26376 10100 26382
rect 10048 26318 10100 26324
rect 9956 26036 10008 26042
rect 9956 25978 10008 25984
rect 9864 25968 9916 25974
rect 9864 25910 9916 25916
rect 9954 25936 10010 25945
rect 9954 25871 10010 25880
rect 9517 25596 9825 25605
rect 9517 25594 9523 25596
rect 9579 25594 9603 25596
rect 9659 25594 9683 25596
rect 9739 25594 9763 25596
rect 9819 25594 9825 25596
rect 9579 25542 9581 25594
rect 9761 25542 9763 25594
rect 9517 25540 9523 25542
rect 9579 25540 9603 25542
rect 9659 25540 9683 25542
rect 9739 25540 9763 25542
rect 9819 25540 9825 25542
rect 9517 25531 9825 25540
rect 9968 25498 9996 25871
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9770 24848 9826 24857
rect 9770 24783 9826 24792
rect 9784 24750 9812 24783
rect 9404 24744 9456 24750
rect 9404 24686 9456 24692
rect 9772 24744 9824 24750
rect 9772 24686 9824 24692
rect 9862 24712 9918 24721
rect 9862 24647 9918 24656
rect 9517 24508 9825 24517
rect 9517 24506 9523 24508
rect 9579 24506 9603 24508
rect 9659 24506 9683 24508
rect 9739 24506 9763 24508
rect 9819 24506 9825 24508
rect 9579 24454 9581 24506
rect 9761 24454 9763 24506
rect 9517 24452 9523 24454
rect 9579 24452 9603 24454
rect 9659 24452 9683 24454
rect 9739 24452 9763 24454
rect 9819 24452 9825 24454
rect 9517 24443 9825 24452
rect 9772 24336 9824 24342
rect 9772 24278 9824 24284
rect 9784 24206 9812 24278
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9876 23866 9904 24647
rect 9968 24410 9996 25230
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9968 23662 9996 24346
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9404 23520 9456 23526
rect 9404 23462 9456 23468
rect 9416 21690 9444 23462
rect 9517 23420 9825 23429
rect 9517 23418 9523 23420
rect 9579 23418 9603 23420
rect 9659 23418 9683 23420
rect 9739 23418 9763 23420
rect 9819 23418 9825 23420
rect 9579 23366 9581 23418
rect 9761 23366 9763 23418
rect 9517 23364 9523 23366
rect 9579 23364 9603 23366
rect 9659 23364 9683 23366
rect 9739 23364 9763 23366
rect 9819 23364 9825 23366
rect 9517 23355 9825 23364
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9772 23112 9824 23118
rect 9600 23072 9772 23100
rect 9600 22982 9628 23072
rect 9772 23054 9824 23060
rect 9588 22976 9640 22982
rect 9588 22918 9640 22924
rect 9517 22332 9825 22341
rect 9517 22330 9523 22332
rect 9579 22330 9603 22332
rect 9659 22330 9683 22332
rect 9739 22330 9763 22332
rect 9819 22330 9825 22332
rect 9579 22278 9581 22330
rect 9761 22278 9763 22330
rect 9517 22276 9523 22278
rect 9579 22276 9603 22278
rect 9659 22276 9683 22278
rect 9739 22276 9763 22278
rect 9819 22276 9825 22278
rect 9517 22267 9825 22276
rect 9968 22234 9996 23258
rect 10060 23050 10088 26318
rect 10152 25974 10180 28154
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10152 24410 10180 24890
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 10048 23044 10100 23050
rect 10048 22986 10100 22992
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9496 21956 9548 21962
rect 9496 21898 9548 21904
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 21078 9444 21490
rect 9508 21457 9536 21898
rect 9600 21894 9628 22170
rect 10244 22166 10272 31726
rect 10322 31376 10378 31385
rect 10322 31311 10378 31320
rect 10336 30938 10364 31311
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10428 30258 10456 32166
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10324 30184 10376 30190
rect 10324 30126 10376 30132
rect 10336 28626 10364 30126
rect 10416 29504 10468 29510
rect 10416 29446 10468 29452
rect 10324 28620 10376 28626
rect 10324 28562 10376 28568
rect 10428 24970 10456 29446
rect 10520 28218 10548 31282
rect 10796 28994 10824 32830
rect 10968 32768 11020 32774
rect 11440 32756 11468 32846
rect 11532 32830 11652 32858
rect 10968 32710 11020 32716
rect 11164 32728 11468 32756
rect 10980 32502 11008 32710
rect 11060 32564 11112 32570
rect 11060 32506 11112 32512
rect 10968 32496 11020 32502
rect 11072 32473 11100 32506
rect 10968 32438 11020 32444
rect 11058 32464 11114 32473
rect 11058 32399 11114 32408
rect 11164 32314 11192 32728
rect 11230 32668 11538 32677
rect 11230 32666 11236 32668
rect 11292 32666 11316 32668
rect 11372 32666 11396 32668
rect 11452 32666 11476 32668
rect 11532 32666 11538 32668
rect 11292 32614 11294 32666
rect 11474 32614 11476 32666
rect 11230 32612 11236 32614
rect 11292 32612 11316 32614
rect 11372 32612 11396 32614
rect 11452 32612 11476 32614
rect 11532 32612 11538 32614
rect 11230 32603 11538 32612
rect 11336 32564 11388 32570
rect 11336 32506 11388 32512
rect 11072 32286 11192 32314
rect 10966 31920 11022 31929
rect 10966 31855 11022 31864
rect 10980 31482 11008 31855
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 10876 30728 10928 30734
rect 10876 30670 10928 30676
rect 10888 29850 10916 30670
rect 11072 30138 11100 32286
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11164 32026 11192 32166
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 11348 31958 11376 32506
rect 11624 32230 11652 32830
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11336 31952 11388 31958
rect 11336 31894 11388 31900
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11532 31686 11560 31758
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11230 31580 11538 31589
rect 11230 31578 11236 31580
rect 11292 31578 11316 31580
rect 11372 31578 11396 31580
rect 11452 31578 11476 31580
rect 11532 31578 11538 31580
rect 11292 31526 11294 31578
rect 11474 31526 11476 31578
rect 11230 31524 11236 31526
rect 11292 31524 11316 31526
rect 11372 31524 11396 31526
rect 11452 31524 11476 31526
rect 11532 31524 11538 31526
rect 11230 31515 11538 31524
rect 11624 31362 11652 32166
rect 11716 31958 11744 33798
rect 11808 33640 11836 34546
rect 11992 34474 12020 35702
rect 12440 35624 12492 35630
rect 12912 35578 12940 36246
rect 13176 36168 13228 36174
rect 13176 36110 13228 36116
rect 13188 35630 13216 36110
rect 12440 35566 12492 35572
rect 12348 35148 12400 35154
rect 12348 35090 12400 35096
rect 12072 35012 12124 35018
rect 12072 34954 12124 34960
rect 12084 34746 12112 34954
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 11980 34468 12032 34474
rect 11980 34410 12032 34416
rect 12268 33998 12296 34546
rect 12256 33992 12308 33998
rect 12176 33940 12256 33946
rect 12176 33934 12308 33940
rect 12176 33918 12296 33934
rect 11808 33612 12020 33640
rect 11888 33516 11940 33522
rect 11888 33458 11940 33464
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11808 32434 11836 32710
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11808 32337 11836 32370
rect 11794 32328 11850 32337
rect 11794 32263 11850 32272
rect 11704 31952 11756 31958
rect 11704 31894 11756 31900
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 11796 31680 11848 31686
rect 11796 31622 11848 31628
rect 11152 31340 11204 31346
rect 11152 31282 11204 31288
rect 11532 31334 11652 31362
rect 11164 30938 11192 31282
rect 11532 31278 11560 31334
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11518 31104 11574 31113
rect 11518 31039 11574 31048
rect 11532 30938 11560 31039
rect 11152 30932 11204 30938
rect 11152 30874 11204 30880
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11230 30492 11538 30501
rect 11230 30490 11236 30492
rect 11292 30490 11316 30492
rect 11372 30490 11396 30492
rect 11452 30490 11476 30492
rect 11532 30490 11538 30492
rect 11292 30438 11294 30490
rect 11474 30438 11476 30490
rect 11230 30436 11236 30438
rect 11292 30436 11316 30438
rect 11372 30436 11396 30438
rect 11452 30436 11476 30438
rect 11532 30436 11538 30438
rect 11230 30427 11538 30436
rect 11612 30184 11664 30190
rect 11072 30110 11192 30138
rect 11612 30126 11664 30132
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29850 11100 29990
rect 10876 29844 10928 29850
rect 10876 29786 10928 29792
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 11060 29640 11112 29646
rect 11060 29582 11112 29588
rect 10796 28966 10916 28994
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 28558 10732 28902
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10796 28558 10824 28698
rect 10692 28552 10744 28558
rect 10612 28512 10692 28540
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10520 25294 10548 27814
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10428 24942 10548 24970
rect 10414 24848 10470 24857
rect 10414 24783 10470 24792
rect 10428 24410 10456 24783
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10336 23866 10364 24210
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10428 23746 10456 24210
rect 10336 23718 10456 23746
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9494 21448 9550 21457
rect 9494 21383 9550 21392
rect 9692 21350 9720 22034
rect 9956 22024 10008 22030
rect 9954 21992 9956 22001
rect 10048 22024 10100 22030
rect 10008 21992 10010 22001
rect 10048 21966 10100 21972
rect 9954 21927 10010 21936
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9876 21457 9904 21626
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9517 21244 9825 21253
rect 9517 21242 9523 21244
rect 9579 21242 9603 21244
rect 9659 21242 9683 21244
rect 9739 21242 9763 21244
rect 9819 21242 9825 21244
rect 9579 21190 9581 21242
rect 9761 21190 9763 21242
rect 9517 21188 9523 21190
rect 9579 21188 9603 21190
rect 9659 21188 9683 21190
rect 9739 21188 9763 21190
rect 9819 21188 9825 21190
rect 9517 21179 9825 21188
rect 9876 21146 9904 21286
rect 9772 21140 9824 21146
rect 9692 21100 9772 21128
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9692 20942 9720 21100
rect 9772 21082 9824 21088
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9864 20936 9916 20942
rect 9864 20878 9916 20884
rect 9876 20602 9904 20878
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9968 20244 9996 21490
rect 9416 20216 9996 20244
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19514 9352 19790
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9324 18426 9352 18702
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 15348 9260 17138
rect 9324 16590 9352 17614
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9324 16046 9352 16526
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15502 9352 15982
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9232 15320 9352 15348
rect 9048 14980 9168 15008
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 9048 14346 9076 14980
rect 9126 14920 9182 14929
rect 9324 14890 9352 15320
rect 9126 14855 9182 14864
rect 9312 14884 9364 14890
rect 9036 14340 9088 14346
rect 9036 14282 9088 14288
rect 8942 14240 8998 14249
rect 8942 14175 8998 14184
rect 8956 13870 8984 14175
rect 9048 13938 9076 14282
rect 9036 13932 9088 13938
rect 9140 13920 9168 14855
rect 9312 14826 9364 14832
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9232 14414 9260 14758
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9232 13938 9260 14010
rect 9036 13874 9088 13880
rect 9122 13892 9168 13920
rect 9220 13932 9272 13938
rect 8944 13864 8996 13870
rect 8944 13806 8996 13812
rect 9034 13832 9090 13841
rect 9034 13767 9090 13776
rect 9122 13784 9150 13892
rect 9220 13874 9272 13880
rect 9048 13734 9076 13767
rect 9122 13756 9260 13784
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8864 12406 8984 12434
rect 8758 11792 8814 11801
rect 8758 11727 8814 11736
rect 8852 11756 8904 11762
rect 8772 4146 8800 11727
rect 8852 11698 8904 11704
rect 8864 11354 8892 11698
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8956 9024 8984 12406
rect 9232 10062 9260 13756
rect 9220 10056 9272 10062
rect 9324 10033 9352 14826
rect 9416 12986 9444 20216
rect 9517 20156 9825 20165
rect 9517 20154 9523 20156
rect 9579 20154 9603 20156
rect 9659 20154 9683 20156
rect 9739 20154 9763 20156
rect 9819 20154 9825 20156
rect 9579 20102 9581 20154
rect 9761 20102 9763 20154
rect 9517 20100 9523 20102
rect 9579 20100 9603 20102
rect 9659 20100 9683 20102
rect 9739 20100 9763 20102
rect 9819 20100 9825 20102
rect 9517 20091 9825 20100
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9678 19272 9734 19281
rect 9678 19207 9680 19216
rect 9732 19207 9734 19216
rect 9680 19178 9732 19184
rect 9784 19156 9812 19994
rect 10060 19802 10088 21966
rect 10140 21684 10192 21690
rect 10140 21626 10192 21632
rect 10152 21078 10180 21626
rect 10140 21072 10192 21078
rect 10336 21026 10364 23718
rect 10520 23644 10548 24942
rect 10612 24206 10640 28512
rect 10692 28494 10744 28500
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10704 25158 10732 25842
rect 10692 25152 10744 25158
rect 10692 25094 10744 25100
rect 10704 24274 10732 25094
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10140 21014 10192 21020
rect 10244 20998 10364 21026
rect 10428 23616 10548 23644
rect 10060 19774 10180 19802
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9864 19372 9916 19378
rect 9916 19332 9996 19360
rect 9864 19314 9916 19320
rect 9784 19128 9904 19156
rect 9517 19068 9825 19077
rect 9517 19066 9523 19068
rect 9579 19066 9603 19068
rect 9659 19066 9683 19068
rect 9739 19066 9763 19068
rect 9819 19066 9825 19068
rect 9579 19014 9581 19066
rect 9761 19014 9763 19066
rect 9517 19012 9523 19014
rect 9579 19012 9603 19014
rect 9659 19012 9683 19014
rect 9739 19012 9763 19014
rect 9819 19012 9825 19014
rect 9517 19003 9825 19012
rect 9678 18864 9734 18873
rect 9876 18834 9904 19128
rect 9678 18799 9734 18808
rect 9864 18828 9916 18834
rect 9692 18290 9720 18799
rect 9864 18770 9916 18776
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9517 17980 9825 17989
rect 9517 17978 9523 17980
rect 9579 17978 9603 17980
rect 9659 17978 9683 17980
rect 9739 17978 9763 17980
rect 9819 17978 9825 17980
rect 9579 17926 9581 17978
rect 9761 17926 9763 17978
rect 9517 17924 9523 17926
rect 9579 17924 9603 17926
rect 9659 17924 9683 17926
rect 9739 17924 9763 17926
rect 9819 17924 9825 17926
rect 9517 17915 9825 17924
rect 9876 17762 9904 18770
rect 9784 17746 9904 17762
rect 9772 17740 9904 17746
rect 9824 17734 9904 17740
rect 9772 17682 9824 17688
rect 9864 17672 9916 17678
rect 9864 17614 9916 17620
rect 9517 16892 9825 16901
rect 9517 16890 9523 16892
rect 9579 16890 9603 16892
rect 9659 16890 9683 16892
rect 9739 16890 9763 16892
rect 9819 16890 9825 16892
rect 9579 16838 9581 16890
rect 9761 16838 9763 16890
rect 9517 16836 9523 16838
rect 9579 16836 9603 16838
rect 9659 16836 9683 16838
rect 9739 16836 9763 16838
rect 9819 16836 9825 16838
rect 9517 16827 9825 16836
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9692 16590 9720 16730
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9600 16114 9628 16390
rect 9876 16182 9904 17614
rect 9864 16176 9916 16182
rect 9864 16118 9916 16124
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9517 15804 9825 15813
rect 9517 15802 9523 15804
rect 9579 15802 9603 15804
rect 9659 15802 9683 15804
rect 9739 15802 9763 15804
rect 9819 15802 9825 15804
rect 9579 15750 9581 15802
rect 9761 15750 9763 15802
rect 9517 15748 9523 15750
rect 9579 15748 9603 15750
rect 9659 15748 9683 15750
rect 9739 15748 9763 15750
rect 9819 15748 9825 15750
rect 9517 15739 9825 15748
rect 9876 15502 9904 15846
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 14804 9720 14894
rect 9692 14776 9904 14804
rect 9517 14716 9825 14725
rect 9517 14714 9523 14716
rect 9579 14714 9603 14716
rect 9659 14714 9683 14716
rect 9739 14714 9763 14716
rect 9819 14714 9825 14716
rect 9579 14662 9581 14714
rect 9761 14662 9763 14714
rect 9517 14660 9523 14662
rect 9579 14660 9603 14662
rect 9659 14660 9683 14662
rect 9739 14660 9763 14662
rect 9819 14660 9825 14662
rect 9517 14651 9825 14660
rect 9517 13628 9825 13637
rect 9517 13626 9523 13628
rect 9579 13626 9603 13628
rect 9659 13626 9683 13628
rect 9739 13626 9763 13628
rect 9819 13626 9825 13628
rect 9579 13574 9581 13626
rect 9761 13574 9763 13626
rect 9517 13572 9523 13574
rect 9579 13572 9603 13574
rect 9659 13572 9683 13574
rect 9739 13572 9763 13574
rect 9819 13572 9825 13574
rect 9517 13563 9825 13572
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9404 12776 9456 12782
rect 9508 12764 9536 13262
rect 9770 12880 9826 12889
rect 9770 12815 9772 12824
rect 9824 12815 9826 12824
rect 9772 12786 9824 12792
rect 9456 12736 9536 12764
rect 9404 12718 9456 12724
rect 9416 10266 9444 12718
rect 9517 12540 9825 12549
rect 9517 12538 9523 12540
rect 9579 12538 9603 12540
rect 9659 12538 9683 12540
rect 9739 12538 9763 12540
rect 9819 12538 9825 12540
rect 9579 12486 9581 12538
rect 9761 12486 9763 12538
rect 9517 12484 9523 12486
rect 9579 12484 9603 12486
rect 9659 12484 9683 12486
rect 9739 12484 9763 12486
rect 9819 12484 9825 12486
rect 9517 12475 9825 12484
rect 9680 12436 9732 12442
rect 9876 12434 9904 14776
rect 9968 14006 9996 19332
rect 10060 19310 10088 19654
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 10152 19009 10180 19774
rect 10138 19000 10194 19009
rect 10138 18935 10194 18944
rect 10152 18766 10180 18935
rect 10140 18760 10192 18766
rect 10046 18728 10102 18737
rect 10140 18702 10192 18708
rect 10046 18663 10102 18672
rect 10060 18630 10088 18663
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10140 17128 10192 17134
rect 10244 17116 10272 20998
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10192 17088 10272 17116
rect 10140 17070 10192 17076
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10060 16250 10088 17002
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10152 16130 10180 16458
rect 10060 16102 10180 16130
rect 10060 14498 10088 16102
rect 10244 15065 10272 17088
rect 10230 15056 10286 15065
rect 10230 14991 10286 15000
rect 10244 14958 10272 14991
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 10152 14618 10180 14826
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10230 14512 10286 14521
rect 10060 14470 10180 14498
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9956 14000 10008 14006
rect 9956 13942 10008 13948
rect 10060 13870 10088 14282
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9954 13424 10010 13433
rect 9954 13359 10010 13368
rect 9968 12646 9996 13359
rect 10152 13190 10180 14470
rect 10230 14447 10286 14456
rect 10244 14414 10272 14447
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13258 10272 14350
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9680 12378 9732 12384
rect 9784 12406 9904 12434
rect 9692 12345 9720 12378
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9784 12102 9812 12406
rect 9954 12200 10010 12209
rect 9954 12135 10010 12144
rect 9968 12102 9996 12135
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9784 11694 9812 12038
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9517 11452 9825 11461
rect 9517 11450 9523 11452
rect 9579 11450 9603 11452
rect 9659 11450 9683 11452
rect 9739 11450 9763 11452
rect 9819 11450 9825 11452
rect 9579 11398 9581 11450
rect 9761 11398 9763 11450
rect 9517 11396 9523 11398
rect 9579 11396 9603 11398
rect 9659 11396 9683 11398
rect 9739 11396 9763 11398
rect 9819 11396 9825 11398
rect 9517 11387 9825 11396
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9692 10606 9720 11290
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9517 10364 9825 10373
rect 9517 10362 9523 10364
rect 9579 10362 9603 10364
rect 9659 10362 9683 10364
rect 9739 10362 9763 10364
rect 9819 10362 9825 10364
rect 9579 10310 9581 10362
rect 9761 10310 9763 10362
rect 9517 10308 9523 10310
rect 9579 10308 9603 10310
rect 9659 10308 9683 10310
rect 9739 10308 9763 10310
rect 9819 10308 9825 10310
rect 9517 10299 9825 10308
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9402 10160 9458 10169
rect 9402 10095 9458 10104
rect 9220 9998 9272 10004
rect 9310 10024 9366 10033
rect 9310 9959 9366 9968
rect 9416 9518 9444 10095
rect 9876 9586 9904 11698
rect 9968 10577 9996 12038
rect 10152 11898 10180 13126
rect 10336 12424 10364 20878
rect 10428 19310 10456 23616
rect 10612 21554 10640 24142
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10704 22778 10732 23802
rect 10692 22772 10744 22778
rect 10692 22714 10744 22720
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10704 21554 10732 22170
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10416 19304 10468 19310
rect 10508 19304 10560 19310
rect 10416 19246 10468 19252
rect 10506 19272 10508 19281
rect 10692 19304 10744 19310
rect 10560 19272 10562 19281
rect 10428 15473 10456 19246
rect 10692 19246 10744 19252
rect 10506 19207 10562 19216
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10520 18193 10548 19110
rect 10704 18970 10732 19246
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10796 18850 10824 28494
rect 10888 28150 10916 28966
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10980 28218 11008 28494
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 10876 28144 10928 28150
rect 10876 28086 10928 28092
rect 10876 27464 10928 27470
rect 10876 27406 10928 27412
rect 10888 25158 10916 27406
rect 11072 27130 11100 29582
rect 11060 27124 11112 27130
rect 11060 27066 11112 27072
rect 11164 27010 11192 30110
rect 11624 29889 11652 30126
rect 11610 29880 11666 29889
rect 11610 29815 11666 29824
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11230 29404 11538 29413
rect 11230 29402 11236 29404
rect 11292 29402 11316 29404
rect 11372 29402 11396 29404
rect 11452 29402 11476 29404
rect 11532 29402 11538 29404
rect 11292 29350 11294 29402
rect 11474 29350 11476 29402
rect 11230 29348 11236 29350
rect 11292 29348 11316 29350
rect 11372 29348 11396 29350
rect 11452 29348 11476 29350
rect 11532 29348 11538 29350
rect 11230 29339 11538 29348
rect 11230 28316 11538 28325
rect 11230 28314 11236 28316
rect 11292 28314 11316 28316
rect 11372 28314 11396 28316
rect 11452 28314 11476 28316
rect 11532 28314 11538 28316
rect 11292 28262 11294 28314
rect 11474 28262 11476 28314
rect 11230 28260 11236 28262
rect 11292 28260 11316 28262
rect 11372 28260 11396 28262
rect 11452 28260 11476 28262
rect 11532 28260 11538 28262
rect 11230 28251 11538 28260
rect 11230 27228 11538 27237
rect 11230 27226 11236 27228
rect 11292 27226 11316 27228
rect 11372 27226 11396 27228
rect 11452 27226 11476 27228
rect 11532 27226 11538 27228
rect 11292 27174 11294 27226
rect 11474 27174 11476 27226
rect 11230 27172 11236 27174
rect 11292 27172 11316 27174
rect 11372 27172 11396 27174
rect 11452 27172 11476 27174
rect 11532 27172 11538 27174
rect 11230 27163 11538 27172
rect 10980 26982 11192 27010
rect 10980 26246 11008 26982
rect 11152 26512 11204 26518
rect 11152 26454 11204 26460
rect 10968 26240 11020 26246
rect 10968 26182 11020 26188
rect 10980 25378 11008 26182
rect 11164 25838 11192 26454
rect 11230 26140 11538 26149
rect 11230 26138 11236 26140
rect 11292 26138 11316 26140
rect 11372 26138 11396 26140
rect 11452 26138 11476 26140
rect 11532 26138 11538 26140
rect 11292 26086 11294 26138
rect 11474 26086 11476 26138
rect 11230 26084 11236 26086
rect 11292 26084 11316 26086
rect 11372 26084 11396 26086
rect 11452 26084 11476 26086
rect 11532 26084 11538 26086
rect 11230 26075 11538 26084
rect 11152 25832 11204 25838
rect 11152 25774 11204 25780
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11072 25498 11100 25638
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 10980 25350 11100 25378
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 10888 24274 10916 24550
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10980 24154 11008 25230
rect 10888 24126 11008 24154
rect 10888 23526 10916 24126
rect 10968 24064 11020 24070
rect 10968 24006 11020 24012
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10876 22976 10928 22982
rect 10876 22918 10928 22924
rect 10888 21078 10916 22918
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10704 18822 10824 18850
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 10506 18184 10562 18193
rect 10506 18119 10562 18128
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10520 17134 10548 18022
rect 10612 17882 10640 18566
rect 10704 18358 10732 18822
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18358 10824 18566
rect 10888 18358 10916 20742
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10704 17882 10732 18294
rect 10784 18216 10836 18222
rect 10784 18158 10836 18164
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10796 17746 10824 18158
rect 10980 18154 11008 24006
rect 11072 23100 11100 25350
rect 11230 25052 11538 25061
rect 11230 25050 11236 25052
rect 11292 25050 11316 25052
rect 11372 25050 11396 25052
rect 11452 25050 11476 25052
rect 11532 25050 11538 25052
rect 11292 24998 11294 25050
rect 11474 24998 11476 25050
rect 11230 24996 11236 24998
rect 11292 24996 11316 24998
rect 11372 24996 11396 24998
rect 11452 24996 11476 24998
rect 11532 24996 11538 24998
rect 11230 24987 11538 24996
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11520 24608 11572 24614
rect 11520 24550 11572 24556
rect 11164 23322 11192 24550
rect 11532 24274 11560 24550
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11230 23964 11538 23973
rect 11230 23962 11236 23964
rect 11292 23962 11316 23964
rect 11372 23962 11396 23964
rect 11452 23962 11476 23964
rect 11532 23962 11538 23964
rect 11292 23910 11294 23962
rect 11474 23910 11476 23962
rect 11230 23908 11236 23910
rect 11292 23908 11316 23910
rect 11372 23908 11396 23910
rect 11452 23908 11476 23910
rect 11532 23908 11538 23910
rect 11230 23899 11538 23908
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11164 23225 11192 23258
rect 11150 23216 11206 23225
rect 11150 23151 11206 23160
rect 11152 23112 11204 23118
rect 11072 23072 11152 23100
rect 11152 23054 11204 23060
rect 11230 22876 11538 22885
rect 11230 22874 11236 22876
rect 11292 22874 11316 22876
rect 11372 22874 11396 22876
rect 11452 22874 11476 22876
rect 11532 22874 11538 22876
rect 11292 22822 11294 22874
rect 11474 22822 11476 22874
rect 11230 22820 11236 22822
rect 11292 22820 11316 22822
rect 11372 22820 11396 22822
rect 11452 22820 11476 22822
rect 11532 22820 11538 22822
rect 11230 22811 11538 22820
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11058 21448 11114 21457
rect 11058 21383 11114 21392
rect 11072 20942 11100 21383
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 11072 18034 11100 20878
rect 11164 18970 11192 22714
rect 11230 21788 11538 21797
rect 11230 21786 11236 21788
rect 11292 21786 11316 21788
rect 11372 21786 11396 21788
rect 11452 21786 11476 21788
rect 11532 21786 11538 21788
rect 11292 21734 11294 21786
rect 11474 21734 11476 21786
rect 11230 21732 11236 21734
rect 11292 21732 11316 21734
rect 11372 21732 11396 21734
rect 11452 21732 11476 21734
rect 11532 21732 11538 21734
rect 11230 21723 11538 21732
rect 11244 21344 11296 21350
rect 11244 21286 11296 21292
rect 11256 20942 11284 21286
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 20806 11284 20878
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11230 20700 11538 20709
rect 11230 20698 11236 20700
rect 11292 20698 11316 20700
rect 11372 20698 11396 20700
rect 11452 20698 11476 20700
rect 11532 20698 11538 20700
rect 11292 20646 11294 20698
rect 11474 20646 11476 20698
rect 11230 20644 11236 20646
rect 11292 20644 11316 20646
rect 11372 20644 11396 20646
rect 11452 20644 11476 20646
rect 11532 20644 11538 20646
rect 11230 20635 11538 20644
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 11256 19825 11284 20402
rect 11532 19922 11560 20470
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 19825 11560 19858
rect 11242 19816 11298 19825
rect 11242 19751 11298 19760
rect 11518 19816 11574 19825
rect 11518 19751 11574 19760
rect 11230 19612 11538 19621
rect 11230 19610 11236 19612
rect 11292 19610 11316 19612
rect 11372 19610 11396 19612
rect 11452 19610 11476 19612
rect 11532 19610 11538 19612
rect 11292 19558 11294 19610
rect 11474 19558 11476 19610
rect 11230 19556 11236 19558
rect 11292 19556 11316 19558
rect 11372 19556 11396 19558
rect 11452 19556 11476 19558
rect 11532 19556 11538 19558
rect 11230 19547 11538 19556
rect 11518 19408 11574 19417
rect 11518 19343 11574 19352
rect 11532 19292 11560 19343
rect 11440 19264 11560 19292
rect 11440 19174 11468 19264
rect 11428 19168 11480 19174
rect 11242 19136 11298 19145
rect 11428 19110 11480 19116
rect 11242 19071 11298 19080
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11256 18714 11284 19071
rect 11440 18834 11468 19110
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 10888 18006 11100 18034
rect 11164 18686 11284 18714
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10508 17128 10560 17134
rect 10508 17070 10560 17076
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10414 15464 10470 15473
rect 10414 15399 10470 15408
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10428 13938 10456 15302
rect 10520 14958 10548 17070
rect 10612 16794 10640 17070
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10796 16697 10824 16934
rect 10888 16833 10916 18006
rect 11058 17912 11114 17921
rect 11058 17847 11114 17856
rect 11072 17678 11100 17847
rect 11060 17672 11112 17678
rect 10980 17632 11060 17660
rect 10874 16824 10930 16833
rect 10874 16759 10930 16768
rect 10782 16688 10838 16697
rect 10782 16623 10838 16632
rect 10888 16572 10916 16759
rect 10796 16544 10916 16572
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15026 10732 15302
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10508 14952 10560 14958
rect 10560 14912 10640 14940
rect 10508 14894 10560 14900
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13326 10456 13874
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10612 12646 10640 14912
rect 10796 14278 10824 16544
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10888 13274 10916 15302
rect 10980 14346 11008 17632
rect 11060 17614 11112 17620
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 11072 13376 11100 17478
rect 11164 14929 11192 18686
rect 11230 18524 11538 18533
rect 11230 18522 11236 18524
rect 11292 18522 11316 18524
rect 11372 18522 11396 18524
rect 11452 18522 11476 18524
rect 11532 18522 11538 18524
rect 11292 18470 11294 18522
rect 11474 18470 11476 18522
rect 11230 18468 11236 18470
rect 11292 18468 11316 18470
rect 11372 18468 11396 18470
rect 11452 18468 11476 18470
rect 11532 18468 11538 18470
rect 11230 18459 11538 18468
rect 11244 18284 11296 18290
rect 11244 18226 11296 18232
rect 11256 17785 11284 18226
rect 11242 17776 11298 17785
rect 11242 17711 11298 17720
rect 11426 17776 11482 17785
rect 11426 17711 11482 17720
rect 11440 17610 11468 17711
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11230 17436 11538 17445
rect 11230 17434 11236 17436
rect 11292 17434 11316 17436
rect 11372 17434 11396 17436
rect 11452 17434 11476 17436
rect 11532 17434 11538 17436
rect 11292 17382 11294 17434
rect 11474 17382 11476 17434
rect 11230 17380 11236 17382
rect 11292 17380 11316 17382
rect 11372 17380 11396 17382
rect 11452 17380 11476 17382
rect 11532 17380 11538 17382
rect 11230 17371 11538 17380
rect 11624 17134 11652 29582
rect 11716 28218 11744 31622
rect 11808 31226 11836 31622
rect 11900 31362 11928 33458
rect 11992 31482 12020 33612
rect 12176 32994 12204 33918
rect 12360 33522 12388 35090
rect 12452 34474 12480 35566
rect 12820 35550 12940 35578
rect 13176 35624 13228 35630
rect 13280 35601 13308 37198
rect 13372 36650 13400 38286
rect 13464 38185 13492 38898
rect 13636 38752 13688 38758
rect 13636 38694 13688 38700
rect 14188 38752 14240 38758
rect 14384 38729 14412 39238
rect 14657 39196 14965 39205
rect 14657 39194 14663 39196
rect 14719 39194 14743 39196
rect 14799 39194 14823 39196
rect 14879 39194 14903 39196
rect 14959 39194 14965 39196
rect 14719 39142 14721 39194
rect 14901 39142 14903 39194
rect 14657 39140 14663 39142
rect 14719 39140 14743 39142
rect 14799 39140 14823 39142
rect 14879 39140 14903 39142
rect 14959 39140 14965 39142
rect 14657 39131 14965 39140
rect 14464 38752 14516 38758
rect 14188 38694 14240 38700
rect 14370 38720 14426 38729
rect 13648 38457 13676 38694
rect 14200 38457 14228 38694
rect 14464 38694 14516 38700
rect 14370 38655 14426 38664
rect 13634 38448 13690 38457
rect 13634 38383 13690 38392
rect 14186 38448 14242 38457
rect 14186 38383 14242 38392
rect 13820 38208 13872 38214
rect 13450 38176 13506 38185
rect 13820 38150 13872 38156
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 13450 38111 13506 38120
rect 13832 37913 13860 38150
rect 13818 37904 13874 37913
rect 13818 37839 13874 37848
rect 13544 37664 13596 37670
rect 13544 37606 13596 37612
rect 13636 37664 13688 37670
rect 13636 37606 13688 37612
rect 14188 37664 14240 37670
rect 14384 37641 14412 38150
rect 14188 37606 14240 37612
rect 14370 37632 14426 37641
rect 13556 37194 13584 37606
rect 13648 37233 13676 37606
rect 14200 37369 14228 37606
rect 14370 37567 14426 37576
rect 14186 37360 14242 37369
rect 14186 37295 14242 37304
rect 13634 37224 13690 37233
rect 13544 37188 13596 37194
rect 13634 37159 13690 37168
rect 13544 37130 13596 37136
rect 13636 37120 13688 37126
rect 13636 37062 13688 37068
rect 14372 37120 14424 37126
rect 14372 37062 14424 37068
rect 13648 36825 13676 37062
rect 13634 36816 13690 36825
rect 13452 36780 13504 36786
rect 13504 36740 13584 36768
rect 13634 36751 13690 36760
rect 13452 36722 13504 36728
rect 13360 36644 13412 36650
rect 13360 36586 13412 36592
rect 13452 36644 13504 36650
rect 13452 36586 13504 36592
rect 13464 36378 13492 36586
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13452 36168 13504 36174
rect 13452 36110 13504 36116
rect 13360 36032 13412 36038
rect 13360 35974 13412 35980
rect 13176 35566 13228 35572
rect 13266 35592 13322 35601
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12440 34468 12492 34474
rect 12440 34410 12492 34416
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 12544 33266 12572 35430
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12360 33238 12572 33266
rect 12176 32966 12296 32994
rect 12072 32836 12124 32842
rect 12072 32778 12124 32784
rect 11980 31476 12032 31482
rect 11980 31418 12032 31424
rect 11900 31334 12020 31362
rect 11808 31198 11928 31226
rect 11796 31136 11848 31142
rect 11796 31078 11848 31084
rect 11808 30938 11836 31078
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11796 30184 11848 30190
rect 11796 30126 11848 30132
rect 11808 29578 11836 30126
rect 11900 30122 11928 31198
rect 11888 30116 11940 30122
rect 11888 30058 11940 30064
rect 11796 29572 11848 29578
rect 11796 29514 11848 29520
rect 11808 29170 11836 29514
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11888 29096 11940 29102
rect 11888 29038 11940 29044
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 11704 28212 11756 28218
rect 11704 28154 11756 28160
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11716 26586 11744 27950
rect 11808 27849 11836 28970
rect 11794 27840 11850 27849
rect 11794 27775 11850 27784
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 11704 26580 11756 26586
rect 11704 26522 11756 26528
rect 11704 25968 11756 25974
rect 11704 25910 11756 25916
rect 11716 25294 11744 25910
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11716 23662 11744 25230
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11808 23118 11836 27406
rect 11900 24410 11928 29038
rect 11992 29016 12020 31334
rect 12084 30938 12112 32778
rect 12164 32428 12216 32434
rect 12164 32370 12216 32376
rect 12176 32026 12204 32370
rect 12164 32020 12216 32026
rect 12164 31962 12216 31968
rect 12268 31686 12296 32966
rect 12256 31680 12308 31686
rect 12256 31622 12308 31628
rect 12164 31408 12216 31414
rect 12164 31350 12216 31356
rect 12072 30932 12124 30938
rect 12072 30874 12124 30880
rect 12072 30048 12124 30054
rect 12072 29990 12124 29996
rect 12084 29730 12112 29990
rect 12176 29850 12204 31350
rect 12268 31278 12296 31622
rect 12256 31272 12308 31278
rect 12256 31214 12308 31220
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12164 29844 12216 29850
rect 12164 29786 12216 29792
rect 12268 29782 12296 31078
rect 12256 29776 12308 29782
rect 12084 29714 12204 29730
rect 12256 29718 12308 29724
rect 12084 29708 12216 29714
rect 12084 29702 12164 29708
rect 12164 29650 12216 29656
rect 12176 29594 12204 29650
rect 12176 29566 12296 29594
rect 11992 28988 12204 29016
rect 11978 28928 12034 28937
rect 11978 28863 12034 28872
rect 11992 28150 12020 28863
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 12084 28082 12112 28494
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11992 27130 12020 27270
rect 11980 27124 12032 27130
rect 11980 27066 12032 27072
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11992 25294 12020 25638
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11900 23066 11928 24142
rect 11992 23730 12020 25230
rect 12084 24970 12112 27406
rect 12176 27112 12204 28988
rect 12268 28966 12296 29566
rect 12256 28960 12308 28966
rect 12256 28902 12308 28908
rect 12268 28762 12296 28902
rect 12256 28756 12308 28762
rect 12256 28698 12308 28704
rect 12360 28694 12388 33238
rect 12636 33153 12664 35022
rect 12716 34536 12768 34542
rect 12716 34478 12768 34484
rect 12728 33862 12756 34478
rect 12820 34474 12848 35550
rect 13266 35527 13322 35536
rect 12944 35388 13252 35397
rect 12944 35386 12950 35388
rect 13006 35386 13030 35388
rect 13086 35386 13110 35388
rect 13166 35386 13190 35388
rect 13246 35386 13252 35388
rect 13006 35334 13008 35386
rect 13188 35334 13190 35386
rect 12944 35332 12950 35334
rect 13006 35332 13030 35334
rect 13086 35332 13110 35334
rect 13166 35332 13190 35334
rect 13246 35332 13252 35334
rect 12944 35323 13252 35332
rect 12900 34944 12952 34950
rect 12900 34886 12952 34892
rect 13176 34944 13228 34950
rect 13176 34886 13228 34892
rect 12912 34746 12940 34886
rect 13188 34746 13216 34886
rect 12900 34740 12952 34746
rect 12900 34682 12952 34688
rect 13176 34740 13228 34746
rect 13176 34682 13228 34688
rect 12808 34468 12860 34474
rect 12808 34410 12860 34416
rect 13268 34400 13320 34406
rect 13268 34342 13320 34348
rect 12944 34300 13252 34309
rect 12944 34298 12950 34300
rect 13006 34298 13030 34300
rect 13086 34298 13110 34300
rect 13166 34298 13190 34300
rect 13246 34298 13252 34300
rect 13006 34246 13008 34298
rect 13188 34246 13190 34298
rect 12944 34244 12950 34246
rect 13006 34244 13030 34246
rect 13086 34244 13110 34246
rect 13166 34244 13190 34246
rect 13246 34244 13252 34246
rect 12944 34235 13252 34244
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12716 33516 12768 33522
rect 12716 33458 12768 33464
rect 12622 33144 12678 33153
rect 12622 33079 12678 33088
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12440 32496 12492 32502
rect 12440 32438 12492 32444
rect 12452 32026 12480 32438
rect 12440 32020 12492 32026
rect 12440 31962 12492 31968
rect 12636 31906 12664 32710
rect 12728 32366 12756 33458
rect 13188 33402 13216 33934
rect 13280 33658 13308 34342
rect 13372 33998 13400 35974
rect 13464 35766 13492 36110
rect 13452 35760 13504 35766
rect 13452 35702 13504 35708
rect 13556 35136 13584 36740
rect 13636 36712 13688 36718
rect 13636 36654 13688 36660
rect 13648 35290 13676 36654
rect 13820 36576 13872 36582
rect 14384 36553 14412 37062
rect 13820 36518 13872 36524
rect 14370 36544 14426 36553
rect 13832 36281 13860 36518
rect 14370 36479 14426 36488
rect 13818 36272 13874 36281
rect 13818 36207 13874 36216
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13740 35737 13768 35974
rect 13726 35728 13782 35737
rect 13726 35663 13782 35672
rect 14004 35692 14056 35698
rect 14004 35634 14056 35640
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13636 35284 13688 35290
rect 13636 35226 13688 35232
rect 13832 35193 13860 35430
rect 13818 35184 13874 35193
rect 13556 35108 13676 35136
rect 13818 35119 13874 35128
rect 13542 35048 13598 35057
rect 13542 34983 13544 34992
rect 13596 34983 13598 34992
rect 13544 34954 13596 34960
rect 13452 34604 13504 34610
rect 13452 34546 13504 34552
rect 13360 33992 13412 33998
rect 13360 33934 13412 33940
rect 13268 33652 13320 33658
rect 13268 33594 13320 33600
rect 13464 33454 13492 34546
rect 13648 34490 13676 35108
rect 13728 35080 13780 35086
rect 13728 35022 13780 35028
rect 13556 34462 13676 34490
rect 13452 33448 13504 33454
rect 13188 33374 13308 33402
rect 13452 33390 13504 33396
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12716 32360 12768 32366
rect 12716 32302 12768 32308
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12544 31890 12664 31906
rect 12532 31884 12664 31890
rect 12584 31878 12664 31884
rect 12532 31826 12584 31832
rect 12624 31816 12676 31822
rect 12622 31784 12624 31793
rect 12676 31784 12678 31793
rect 12622 31719 12678 31728
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12452 31113 12480 31622
rect 12624 31136 12676 31142
rect 12438 31104 12494 31113
rect 12624 31078 12676 31084
rect 12438 31039 12494 31048
rect 12636 30938 12664 31078
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 12440 30728 12492 30734
rect 12728 30682 12756 32166
rect 12440 30670 12492 30676
rect 12452 29510 12480 30670
rect 12636 30654 12756 30682
rect 12636 30054 12664 30654
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12624 29640 12676 29646
rect 12624 29582 12676 29588
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12636 28914 12664 29582
rect 12728 29306 12756 30534
rect 12820 30258 12848 33254
rect 12944 33212 13252 33221
rect 12944 33210 12950 33212
rect 13006 33210 13030 33212
rect 13086 33210 13110 33212
rect 13166 33210 13190 33212
rect 13246 33210 13252 33212
rect 13006 33158 13008 33210
rect 13188 33158 13190 33210
rect 12944 33156 12950 33158
rect 13006 33156 13030 33158
rect 13086 33156 13110 33158
rect 13166 33156 13190 33158
rect 13246 33156 13252 33158
rect 12944 33147 13252 33156
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 12912 32416 12940 32846
rect 13280 32570 13308 33374
rect 13360 32904 13412 32910
rect 13360 32846 13412 32852
rect 13268 32564 13320 32570
rect 13268 32506 13320 32512
rect 12912 32388 13308 32416
rect 12944 32124 13252 32133
rect 12944 32122 12950 32124
rect 13006 32122 13030 32124
rect 13086 32122 13110 32124
rect 13166 32122 13190 32124
rect 13246 32122 13252 32124
rect 13006 32070 13008 32122
rect 13188 32070 13190 32122
rect 12944 32068 12950 32070
rect 13006 32068 13030 32070
rect 13086 32068 13110 32070
rect 13166 32068 13190 32070
rect 13246 32068 13252 32070
rect 12944 32059 13252 32068
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 13004 31385 13032 31758
rect 12990 31376 13046 31385
rect 12990 31311 13046 31320
rect 13280 31210 13308 32388
rect 13372 32314 13400 32846
rect 13556 32337 13584 34462
rect 13636 34400 13688 34406
rect 13636 34342 13688 34348
rect 13648 34105 13676 34342
rect 13740 34134 13768 35022
rect 13912 35012 13964 35018
rect 13912 34954 13964 34960
rect 13924 34649 13952 34954
rect 13910 34640 13966 34649
rect 13910 34575 13966 34584
rect 13728 34128 13780 34134
rect 13634 34096 13690 34105
rect 13728 34070 13780 34076
rect 13634 34031 13690 34040
rect 13820 34060 13872 34066
rect 13820 34002 13872 34008
rect 13728 33584 13780 33590
rect 13728 33526 13780 33532
rect 13636 33312 13688 33318
rect 13636 33254 13688 33260
rect 13648 33017 13676 33254
rect 13740 33114 13768 33526
rect 13728 33108 13780 33114
rect 13728 33050 13780 33056
rect 13634 33008 13690 33017
rect 13634 32943 13690 32952
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13636 32360 13688 32366
rect 13542 32328 13598 32337
rect 13372 32286 13492 32314
rect 13360 31680 13412 31686
rect 13360 31622 13412 31628
rect 13268 31204 13320 31210
rect 13268 31146 13320 31152
rect 13372 31113 13400 31622
rect 13464 31249 13492 32286
rect 13636 32302 13688 32308
rect 13542 32263 13598 32272
rect 13450 31240 13506 31249
rect 13648 31226 13676 32302
rect 13740 31929 13768 32370
rect 13726 31920 13782 31929
rect 13726 31855 13782 31864
rect 13648 31198 13768 31226
rect 13450 31175 13506 31184
rect 13544 31136 13596 31142
rect 13358 31104 13414 31113
rect 13544 31078 13596 31084
rect 13636 31136 13688 31142
rect 13636 31078 13688 31084
rect 12944 31036 13252 31045
rect 13358 31039 13414 31048
rect 12944 31034 12950 31036
rect 13006 31034 13030 31036
rect 13086 31034 13110 31036
rect 13166 31034 13190 31036
rect 13246 31034 13252 31036
rect 13006 30982 13008 31034
rect 13188 30982 13190 31034
rect 12944 30980 12950 30982
rect 13006 30980 13030 30982
rect 13086 30980 13110 30982
rect 13166 30980 13190 30982
rect 13246 30980 13252 30982
rect 12944 30971 13252 30980
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 12900 30660 12952 30666
rect 12900 30602 12952 30608
rect 12992 30660 13044 30666
rect 12992 30602 13044 30608
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 12912 30297 12940 30602
rect 12898 30288 12954 30297
rect 12808 30252 12860 30258
rect 12898 30223 12954 30232
rect 12808 30194 12860 30200
rect 13004 30036 13032 30602
rect 13372 30297 13400 30602
rect 13358 30288 13414 30297
rect 13358 30223 13414 30232
rect 13360 30184 13412 30190
rect 13360 30126 13412 30132
rect 12820 30008 13032 30036
rect 12820 29306 12848 30008
rect 12944 29948 13252 29957
rect 12944 29946 12950 29948
rect 13006 29946 13030 29948
rect 13086 29946 13110 29948
rect 13166 29946 13190 29948
rect 13246 29946 13252 29948
rect 13006 29894 13008 29946
rect 13188 29894 13190 29946
rect 12944 29892 12950 29894
rect 13006 29892 13030 29894
rect 13086 29892 13110 29894
rect 13166 29892 13190 29894
rect 13246 29892 13252 29894
rect 12944 29883 13252 29892
rect 12716 29300 12768 29306
rect 12716 29242 12768 29248
rect 12808 29300 12860 29306
rect 12808 29242 12860 29248
rect 12898 29200 12954 29209
rect 12898 29135 12900 29144
rect 12952 29135 12954 29144
rect 12992 29164 13044 29170
rect 12900 29106 12952 29112
rect 12992 29106 13044 29112
rect 13004 29016 13032 29106
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 12820 28988 13032 29016
rect 12636 28886 12756 28914
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12348 28688 12400 28694
rect 12348 28630 12400 28636
rect 12636 28558 12664 28698
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 12348 28416 12400 28422
rect 12348 28358 12400 28364
rect 12360 27470 12388 28358
rect 12624 28076 12676 28082
rect 12544 28036 12624 28064
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12544 27146 12572 28036
rect 12624 28018 12676 28024
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12360 27130 12572 27146
rect 12636 27130 12664 27270
rect 12348 27124 12572 27130
rect 12176 27084 12296 27112
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12176 26489 12204 26930
rect 12162 26480 12218 26489
rect 12162 26415 12218 26424
rect 12268 25106 12296 27084
rect 12400 27118 12572 27124
rect 12624 27124 12676 27130
rect 12348 27066 12400 27072
rect 12624 27066 12676 27072
rect 12530 27024 12586 27033
rect 12530 26959 12586 26968
rect 12348 26920 12400 26926
rect 12400 26868 12480 26874
rect 12348 26862 12480 26868
rect 12360 26846 12480 26862
rect 12348 26784 12400 26790
rect 12348 26726 12400 26732
rect 12360 25945 12388 26726
rect 12452 26042 12480 26846
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12346 25936 12402 25945
rect 12346 25871 12402 25880
rect 12544 25838 12572 26959
rect 12728 26330 12756 28886
rect 12820 27878 12848 28988
rect 12944 28860 13252 28869
rect 12944 28858 12950 28860
rect 13006 28858 13030 28860
rect 13086 28858 13110 28860
rect 13166 28858 13190 28860
rect 13246 28858 13252 28860
rect 13006 28806 13008 28858
rect 13188 28806 13190 28858
rect 12944 28804 12950 28806
rect 13006 28804 13030 28806
rect 13086 28804 13110 28806
rect 13166 28804 13190 28806
rect 13246 28804 13252 28806
rect 12944 28795 13252 28804
rect 12900 28552 12952 28558
rect 12900 28494 12952 28500
rect 12912 28218 12940 28494
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 12944 27772 13252 27781
rect 12944 27770 12950 27772
rect 13006 27770 13030 27772
rect 13086 27770 13110 27772
rect 13166 27770 13190 27772
rect 13246 27770 13252 27772
rect 13006 27718 13008 27770
rect 13188 27718 13190 27770
rect 12944 27716 12950 27718
rect 13006 27716 13030 27718
rect 13086 27716 13110 27718
rect 13166 27716 13190 27718
rect 13246 27716 13252 27718
rect 12944 27707 13252 27716
rect 13084 27464 13136 27470
rect 12636 26302 12756 26330
rect 12820 27424 13084 27452
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12532 25832 12584 25838
rect 12532 25774 12584 25780
rect 12452 25498 12480 25774
rect 12544 25702 12572 25774
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12636 25514 12664 26302
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12728 25906 12756 26182
rect 12820 26081 12848 27424
rect 13084 27406 13136 27412
rect 12900 27328 12952 27334
rect 12900 27270 12952 27276
rect 12990 27296 13046 27305
rect 12912 27130 12940 27270
rect 12990 27231 13046 27240
rect 12900 27124 12952 27130
rect 13004 27112 13032 27231
rect 13084 27124 13136 27130
rect 13004 27084 13084 27112
rect 12900 27066 12952 27072
rect 13084 27066 13136 27072
rect 13280 26874 13308 29038
rect 13372 27033 13400 30126
rect 13464 29850 13492 30738
rect 13452 29844 13504 29850
rect 13452 29786 13504 29792
rect 13556 28914 13584 31078
rect 13648 29753 13676 31078
rect 13740 30394 13768 31198
rect 13728 30388 13780 30394
rect 13728 30330 13780 30336
rect 13832 29782 13860 34002
rect 14016 33930 14044 35634
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14096 34944 14148 34950
rect 14096 34886 14148 34892
rect 13912 33924 13964 33930
rect 13912 33866 13964 33872
rect 14004 33924 14056 33930
rect 14004 33866 14056 33872
rect 13924 33561 13952 33866
rect 13910 33552 13966 33561
rect 13910 33487 13966 33496
rect 14108 32910 14136 34886
rect 14188 34400 14240 34406
rect 14384 34377 14412 35430
rect 14188 34342 14240 34348
rect 14370 34368 14426 34377
rect 14200 34105 14228 34342
rect 14370 34303 14426 34312
rect 14186 34096 14242 34105
rect 14186 34031 14242 34040
rect 14372 33856 14424 33862
rect 14372 33798 14424 33804
rect 14280 33380 14332 33386
rect 14280 33322 14332 33328
rect 14188 33312 14240 33318
rect 14188 33254 14240 33260
rect 14200 33017 14228 33254
rect 14186 33008 14242 33017
rect 14186 32943 14242 32952
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 14292 32858 14320 33322
rect 14384 33289 14412 33798
rect 14370 33280 14426 33289
rect 14370 33215 14426 33224
rect 14292 32830 14412 32858
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14292 32473 14320 32710
rect 14278 32464 14334 32473
rect 14188 32428 14240 32434
rect 14278 32399 14334 32408
rect 14188 32370 14240 32376
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 13924 31929 13952 32166
rect 13910 31920 13966 31929
rect 13910 31855 13966 31864
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13924 30841 13952 31622
rect 14016 31385 14044 32166
rect 14200 32026 14228 32370
rect 14384 32314 14412 32830
rect 14292 32286 14412 32314
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14188 31680 14240 31686
rect 14188 31622 14240 31628
rect 14002 31376 14058 31385
rect 14002 31311 14058 31320
rect 13910 30832 13966 30841
rect 13910 30767 13966 30776
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13820 29776 13872 29782
rect 13634 29744 13690 29753
rect 13820 29718 13872 29724
rect 13634 29679 13690 29688
rect 13820 29640 13872 29646
rect 13924 29617 13952 30058
rect 13820 29582 13872 29588
rect 13910 29608 13966 29617
rect 13464 28886 13584 28914
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13464 27554 13492 28886
rect 13648 28665 13676 28902
rect 13832 28762 13860 29582
rect 13910 29543 13966 29552
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13634 28656 13690 28665
rect 13634 28591 13690 28600
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 13556 27674 13584 28494
rect 13820 28416 13872 28422
rect 13820 28358 13872 28364
rect 13832 28121 13860 28358
rect 13924 28150 13952 29446
rect 14016 29170 14044 30194
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 14004 29164 14056 29170
rect 14004 29106 14056 29112
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 13912 28144 13964 28150
rect 13818 28112 13874 28121
rect 13912 28086 13964 28092
rect 13818 28047 13874 28056
rect 13636 27872 13688 27878
rect 13636 27814 13688 27820
rect 13544 27668 13596 27674
rect 13544 27610 13596 27616
rect 13648 27577 13676 27814
rect 13634 27568 13690 27577
rect 13464 27526 13584 27554
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13464 27062 13492 27406
rect 13452 27056 13504 27062
rect 13358 27024 13414 27033
rect 13452 26998 13504 27004
rect 13358 26959 13414 26968
rect 13280 26846 13492 26874
rect 13268 26784 13320 26790
rect 13268 26726 13320 26732
rect 12944 26684 13252 26693
rect 12944 26682 12950 26684
rect 13006 26682 13030 26684
rect 13086 26682 13110 26684
rect 13166 26682 13190 26684
rect 13246 26682 13252 26684
rect 13006 26630 13008 26682
rect 13188 26630 13190 26682
rect 12944 26628 12950 26630
rect 13006 26628 13030 26630
rect 13086 26628 13110 26630
rect 13166 26628 13190 26630
rect 13246 26628 13252 26630
rect 12944 26619 13252 26628
rect 13280 26217 13308 26726
rect 13266 26208 13322 26217
rect 13266 26143 13322 26152
rect 12806 26072 12862 26081
rect 13464 26058 13492 26846
rect 13556 26382 13584 27526
rect 13634 27503 13690 27512
rect 13636 27396 13688 27402
rect 13636 27338 13688 27344
rect 13912 27396 13964 27402
rect 13912 27338 13964 27344
rect 13544 26376 13596 26382
rect 13544 26318 13596 26324
rect 13648 26330 13676 27338
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13740 26586 13768 27270
rect 13924 27033 13952 27338
rect 13910 27024 13966 27033
rect 14016 26994 14044 28494
rect 14108 27470 14136 29446
rect 14200 29238 14228 31622
rect 14292 31414 14320 32286
rect 14372 32224 14424 32230
rect 14370 32192 14372 32201
rect 14424 32192 14426 32201
rect 14370 32127 14426 32136
rect 14280 31408 14332 31414
rect 14280 31350 14332 31356
rect 14280 30048 14332 30054
rect 14280 29990 14332 29996
rect 14188 29232 14240 29238
rect 14292 29209 14320 29990
rect 14372 29572 14424 29578
rect 14372 29514 14424 29520
rect 14188 29174 14240 29180
rect 14278 29200 14334 29209
rect 14278 29135 14334 29144
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14200 28665 14228 28902
rect 14186 28656 14242 28665
rect 14186 28591 14242 28600
rect 14384 28558 14412 29514
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14372 28416 14424 28422
rect 14372 28358 14424 28364
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14200 27577 14228 27814
rect 14186 27568 14242 27577
rect 14186 27503 14242 27512
rect 14096 27464 14148 27470
rect 14096 27406 14148 27412
rect 14292 27282 14320 28154
rect 14384 27849 14412 28358
rect 14370 27840 14426 27849
rect 14370 27775 14426 27784
rect 14108 27254 14320 27282
rect 13910 26959 13966 26968
rect 14004 26988 14056 26994
rect 14004 26930 14056 26936
rect 13820 26784 13872 26790
rect 13818 26752 13820 26761
rect 13872 26752 13874 26761
rect 13818 26687 13874 26696
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 13648 26302 13768 26330
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13464 26030 13584 26058
rect 12806 26007 12862 26016
rect 13452 25968 13504 25974
rect 13452 25910 13504 25916
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 13360 25900 13412 25906
rect 13360 25842 13412 25848
rect 12944 25596 13252 25605
rect 12944 25594 12950 25596
rect 13006 25594 13030 25596
rect 13086 25594 13110 25596
rect 13166 25594 13190 25596
rect 13246 25594 13252 25596
rect 13006 25542 13008 25594
rect 13188 25542 13190 25594
rect 12944 25540 12950 25542
rect 13006 25540 13030 25542
rect 13086 25540 13110 25542
rect 13166 25540 13190 25542
rect 13246 25540 13252 25542
rect 12944 25531 13252 25540
rect 12440 25492 12492 25498
rect 12636 25486 12756 25514
rect 12440 25434 12492 25440
rect 12268 25078 12388 25106
rect 12084 24942 12296 24970
rect 12072 24812 12124 24818
rect 12072 24754 12124 24760
rect 12084 23905 12112 24754
rect 12070 23896 12126 23905
rect 12070 23831 12126 23840
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11900 23038 12020 23066
rect 11888 22976 11940 22982
rect 11888 22918 11940 22924
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11796 22024 11848 22030
rect 11796 21966 11848 21972
rect 11716 21350 11744 21966
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11808 20777 11836 21966
rect 11900 21010 11928 22918
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11888 20800 11940 20806
rect 11794 20768 11850 20777
rect 11888 20742 11940 20748
rect 11794 20703 11850 20712
rect 11900 20618 11928 20742
rect 11716 20590 11928 20618
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 16590 11284 16934
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11230 16348 11538 16357
rect 11230 16346 11236 16348
rect 11292 16346 11316 16348
rect 11372 16346 11396 16348
rect 11452 16346 11476 16348
rect 11532 16346 11538 16348
rect 11292 16294 11294 16346
rect 11474 16294 11476 16346
rect 11230 16292 11236 16294
rect 11292 16292 11316 16294
rect 11372 16292 11396 16294
rect 11452 16292 11476 16294
rect 11532 16292 11538 16294
rect 11230 16283 11538 16292
rect 11624 16232 11652 17070
rect 11532 16204 11652 16232
rect 11532 15609 11560 16204
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15638 11652 15846
rect 11612 15632 11664 15638
rect 11518 15600 11574 15609
rect 11612 15574 11664 15580
rect 11518 15535 11574 15544
rect 11230 15260 11538 15269
rect 11230 15258 11236 15260
rect 11292 15258 11316 15260
rect 11372 15258 11396 15260
rect 11452 15258 11476 15260
rect 11532 15258 11538 15260
rect 11292 15206 11294 15258
rect 11474 15206 11476 15258
rect 11230 15204 11236 15206
rect 11292 15204 11316 15206
rect 11372 15204 11396 15206
rect 11452 15204 11476 15206
rect 11532 15204 11538 15206
rect 11230 15195 11538 15204
rect 11150 14920 11206 14929
rect 11150 14855 11206 14864
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11164 14074 11192 14282
rect 11230 14172 11538 14181
rect 11230 14170 11236 14172
rect 11292 14170 11316 14172
rect 11372 14170 11396 14172
rect 11452 14170 11476 14172
rect 11532 14170 11538 14172
rect 11292 14118 11294 14170
rect 11474 14118 11476 14170
rect 11230 14116 11236 14118
rect 11292 14116 11316 14118
rect 11372 14116 11396 14118
rect 11452 14116 11476 14118
rect 11532 14116 11538 14118
rect 11230 14107 11538 14116
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11072 13348 11192 13376
rect 10888 13246 11100 13274
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10520 12434 10548 12582
rect 10244 12396 10364 12424
rect 10428 12406 10548 12434
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9954 10568 10010 10577
rect 9954 10503 10010 10512
rect 9968 9722 9996 10503
rect 10244 10305 10272 12396
rect 10428 12322 10456 12406
rect 10336 12306 10456 12322
rect 10324 12300 10456 12306
rect 10376 12294 10456 12300
rect 10324 12242 10376 12248
rect 10704 12186 10732 13126
rect 10782 12336 10838 12345
rect 10782 12271 10838 12280
rect 10876 12300 10928 12306
rect 10428 12170 10732 12186
rect 10796 12170 10824 12271
rect 10876 12242 10928 12248
rect 10416 12164 10732 12170
rect 10468 12158 10732 12164
rect 10784 12164 10836 12170
rect 10416 12106 10468 12112
rect 10784 12106 10836 12112
rect 10888 12102 10916 12242
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10704 11762 10732 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10230 10296 10286 10305
rect 10230 10231 10286 10240
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 10244 9625 10272 10231
rect 10428 10198 10456 11086
rect 10416 10192 10468 10198
rect 10416 10134 10468 10140
rect 10428 10044 10456 10134
rect 10336 10016 10456 10044
rect 10508 10056 10560 10062
rect 10230 9616 10286 9625
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9968 9574 10230 9602
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 8956 8996 9076 9024
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8864 6322 8892 8910
rect 8956 6322 8984 8996
rect 9048 8906 9076 8996
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 9140 8090 9168 9454
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9048 7410 9076 7754
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9140 7342 9168 7822
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 5234 8984 6258
rect 9140 5914 9168 7278
rect 9324 6254 9352 8774
rect 9416 7886 9444 9454
rect 9517 9276 9825 9285
rect 9517 9274 9523 9276
rect 9579 9274 9603 9276
rect 9659 9274 9683 9276
rect 9739 9274 9763 9276
rect 9819 9274 9825 9276
rect 9579 9222 9581 9274
rect 9761 9222 9763 9274
rect 9517 9220 9523 9222
rect 9579 9220 9603 9222
rect 9659 9220 9683 9222
rect 9739 9220 9763 9222
rect 9819 9220 9825 9222
rect 9517 9211 9825 9220
rect 9968 9160 9996 9574
rect 10230 9551 10286 9560
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 10140 9444 10192 9450
rect 10140 9386 10192 9392
rect 10152 9178 10180 9386
rect 9784 9132 9996 9160
rect 10140 9172 10192 9178
rect 9678 8936 9734 8945
rect 9678 8871 9734 8880
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9508 8498 9536 8735
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9692 8430 9720 8871
rect 9784 8498 9812 9132
rect 10140 9114 10192 9120
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9517 8188 9825 8197
rect 9517 8186 9523 8188
rect 9579 8186 9603 8188
rect 9659 8186 9683 8188
rect 9739 8186 9763 8188
rect 9819 8186 9825 8188
rect 9579 8134 9581 8186
rect 9761 8134 9763 8186
rect 9517 8132 9523 8134
rect 9579 8132 9603 8134
rect 9659 8132 9683 8134
rect 9739 8132 9763 8134
rect 9819 8132 9825 8134
rect 9517 8123 9825 8132
rect 9770 7984 9826 7993
rect 9770 7919 9772 7928
rect 9824 7919 9826 7928
rect 9772 7890 9824 7896
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9586 7848 9642 7857
rect 9586 7783 9642 7792
rect 9600 7546 9628 7783
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9517 7100 9825 7109
rect 9517 7098 9523 7100
rect 9579 7098 9603 7100
rect 9659 7098 9683 7100
rect 9739 7098 9763 7100
rect 9819 7098 9825 7100
rect 9579 7046 9581 7098
rect 9761 7046 9763 7098
rect 9517 7044 9523 7046
rect 9579 7044 9603 7046
rect 9659 7044 9683 7046
rect 9739 7044 9763 7046
rect 9819 7044 9825 7046
rect 9517 7035 9825 7044
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9324 5710 9352 6190
rect 9416 6186 9444 6802
rect 9876 6798 9904 8978
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9968 8838 9996 8910
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9968 8022 9996 8570
rect 10152 8537 10180 9114
rect 10244 8838 10272 9454
rect 10336 9217 10364 10016
rect 10508 9998 10560 10004
rect 10520 9897 10548 9998
rect 10506 9888 10562 9897
rect 10506 9823 10562 9832
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10428 9353 10456 9658
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10520 9382 10548 9454
rect 10508 9376 10560 9382
rect 10414 9344 10470 9353
rect 10508 9318 10560 9324
rect 10414 9279 10470 9288
rect 10322 9208 10378 9217
rect 10322 9143 10378 9152
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10244 8634 10272 8774
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10336 8548 10364 8978
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 10302 8520 10364 8548
rect 10048 8356 10100 8362
rect 10302 8344 10330 8520
rect 10428 8498 10456 9279
rect 10612 8498 10640 11494
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10704 9722 10732 11290
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 9042 10732 9522
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8809 10732 8842
rect 10690 8800 10746 8809
rect 10690 8735 10746 8744
rect 10796 8514 10824 11834
rect 10888 11830 10916 12038
rect 10876 11824 10928 11830
rect 10876 11766 10928 11772
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 9738 10916 11630
rect 11072 10062 11100 13246
rect 11164 11898 11192 13348
rect 11440 13297 11468 13670
rect 11532 13394 11560 13806
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11426 13288 11482 13297
rect 11426 13223 11482 13232
rect 11230 13084 11538 13093
rect 11230 13082 11236 13084
rect 11292 13082 11316 13084
rect 11372 13082 11396 13084
rect 11452 13082 11476 13084
rect 11532 13082 11538 13084
rect 11292 13030 11294 13082
rect 11474 13030 11476 13082
rect 11230 13028 11236 13030
rect 11292 13028 11316 13030
rect 11372 13028 11396 13030
rect 11452 13028 11476 13030
rect 11532 13028 11538 13030
rect 11230 13019 11538 13028
rect 11624 12442 11652 15574
rect 11716 15026 11744 20590
rect 11992 20482 12020 23038
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12084 22001 12112 22034
rect 12070 21992 12126 22001
rect 12070 21927 12126 21936
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11900 20454 12020 20482
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11808 19145 11836 19994
rect 11900 19854 11928 20454
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11794 19136 11850 19145
rect 11794 19071 11850 19080
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11808 18290 11836 18906
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11808 17184 11836 18226
rect 11900 17610 11928 19790
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11992 17338 12020 20334
rect 12084 20330 12112 21286
rect 12268 20466 12296 24942
rect 12360 23866 12388 25078
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12452 23712 12480 24754
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12452 23684 12572 23712
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12360 22148 12388 23598
rect 12544 22216 12572 23684
rect 12636 23662 12664 24006
rect 12624 23656 12676 23662
rect 12624 23598 12676 23604
rect 12728 23338 12756 25486
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12636 23310 12756 23338
rect 12820 25276 12848 25434
rect 12900 25288 12952 25294
rect 12820 25248 12900 25276
rect 12820 23644 12848 25248
rect 12900 25230 12952 25236
rect 13372 24614 13400 25842
rect 13268 24608 13320 24614
rect 13268 24550 13320 24556
rect 13360 24608 13412 24614
rect 13360 24550 13412 24556
rect 12944 24508 13252 24517
rect 12944 24506 12950 24508
rect 13006 24506 13030 24508
rect 13086 24506 13110 24508
rect 13166 24506 13190 24508
rect 13246 24506 13252 24508
rect 13006 24454 13008 24506
rect 13188 24454 13190 24506
rect 12944 24452 12950 24454
rect 13006 24452 13030 24454
rect 13086 24452 13110 24454
rect 13166 24452 13190 24454
rect 13246 24452 13252 24454
rect 12944 24443 13252 24452
rect 13280 23746 13308 24550
rect 13464 24342 13492 25910
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13188 23730 13308 23746
rect 13176 23724 13308 23730
rect 13228 23718 13308 23724
rect 13176 23666 13228 23672
rect 12992 23656 13044 23662
rect 12820 23616 12992 23644
rect 12636 22438 12664 23310
rect 12820 23202 12848 23616
rect 12992 23598 13044 23604
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13360 23520 13412 23526
rect 13360 23462 13412 23468
rect 12944 23420 13252 23429
rect 12944 23418 12950 23420
rect 13006 23418 13030 23420
rect 13086 23418 13110 23420
rect 13166 23418 13190 23420
rect 13246 23418 13252 23420
rect 13006 23366 13008 23418
rect 13188 23366 13190 23418
rect 12944 23364 12950 23366
rect 13006 23364 13030 23366
rect 13086 23364 13110 23366
rect 13166 23364 13190 23366
rect 13246 23364 13252 23366
rect 12944 23355 13252 23364
rect 12728 23174 12848 23202
rect 12624 22432 12676 22438
rect 12624 22374 12676 22380
rect 12544 22188 12664 22216
rect 12360 22120 12572 22148
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12072 20324 12124 20330
rect 12072 20266 12124 20272
rect 12084 18766 12112 20266
rect 12176 19514 12204 20402
rect 12360 19854 12388 21490
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12452 20534 12480 20878
rect 12440 20528 12492 20534
rect 12440 20470 12492 20476
rect 12440 20392 12492 20398
rect 12438 20360 12440 20369
rect 12492 20360 12494 20369
rect 12438 20295 12494 20304
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 20058 12480 20198
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12254 19408 12310 19417
rect 12254 19343 12310 19352
rect 12440 19372 12492 19378
rect 12268 18970 12296 19343
rect 12440 19314 12492 19320
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18442 12112 18702
rect 12084 18414 12296 18442
rect 12164 18352 12216 18358
rect 12084 18312 12164 18340
rect 12084 17746 12112 18312
rect 12164 18294 12216 18300
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11806 17156 11836 17184
rect 11806 17082 11834 17156
rect 11806 17054 12020 17082
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11900 16658 11928 16934
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11794 15872 11850 15881
rect 11794 15807 11850 15816
rect 11808 15570 11836 15807
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11704 13864 11756 13870
rect 11704 13806 11756 13812
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11610 12336 11666 12345
rect 11610 12271 11612 12280
rect 11664 12271 11666 12280
rect 11612 12242 11664 12248
rect 11230 11996 11538 12005
rect 11230 11994 11236 11996
rect 11292 11994 11316 11996
rect 11372 11994 11396 11996
rect 11452 11994 11476 11996
rect 11532 11994 11538 11996
rect 11292 11942 11294 11994
rect 11474 11942 11476 11994
rect 11230 11940 11236 11942
rect 11292 11940 11316 11942
rect 11372 11940 11396 11942
rect 11452 11940 11476 11942
rect 11532 11940 11538 11942
rect 11230 11931 11538 11940
rect 11624 11898 11652 12242
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10888 9710 11100 9738
rect 10966 9616 11022 9625
rect 10966 9551 11022 9560
rect 10980 9042 11008 9551
rect 11072 9353 11100 9710
rect 11164 9450 11192 11630
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11256 11150 11284 11290
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11716 11014 11744 13806
rect 11808 13326 11836 15370
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12345 11836 12786
rect 11794 12336 11850 12345
rect 11794 12271 11850 12280
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11230 10908 11538 10917
rect 11230 10906 11236 10908
rect 11292 10906 11316 10908
rect 11372 10906 11396 10908
rect 11452 10906 11476 10908
rect 11532 10906 11538 10908
rect 11292 10854 11294 10906
rect 11474 10854 11476 10906
rect 11230 10852 11236 10854
rect 11292 10852 11316 10854
rect 11372 10852 11396 10854
rect 11452 10852 11476 10854
rect 11532 10852 11538 10854
rect 11230 10843 11538 10852
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11230 9820 11538 9829
rect 11230 9818 11236 9820
rect 11292 9818 11316 9820
rect 11372 9818 11396 9820
rect 11452 9818 11476 9820
rect 11532 9818 11538 9820
rect 11292 9766 11294 9818
rect 11474 9766 11476 9818
rect 11230 9764 11236 9766
rect 11292 9764 11316 9766
rect 11372 9764 11396 9766
rect 11452 9764 11476 9766
rect 11532 9764 11538 9766
rect 11230 9755 11538 9764
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11334 9616 11390 9625
rect 11334 9551 11336 9560
rect 11388 9551 11390 9560
rect 11336 9522 11388 9528
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 11058 9344 11114 9353
rect 11058 9279 11114 9288
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10888 8634 10916 8842
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10600 8492 10652 8498
rect 10796 8486 11008 8514
rect 10600 8434 10652 8440
rect 10302 8316 10364 8344
rect 10048 8298 10100 8304
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 10060 7954 10088 8298
rect 10336 8265 10364 8316
rect 10416 8288 10468 8294
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10322 8256 10378 8265
rect 10416 8230 10468 8236
rect 10322 8191 10378 8200
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9968 7002 9996 7414
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10060 6934 10088 7890
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6322 9720 6666
rect 9784 6610 9812 6734
rect 9956 6656 10008 6662
rect 9784 6582 9904 6610
rect 9956 6598 10008 6604
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 9416 4010 9444 6122
rect 9517 6012 9825 6021
rect 9517 6010 9523 6012
rect 9579 6010 9603 6012
rect 9659 6010 9683 6012
rect 9739 6010 9763 6012
rect 9819 6010 9825 6012
rect 9579 5958 9581 6010
rect 9761 5958 9763 6010
rect 9517 5956 9523 5958
rect 9579 5956 9603 5958
rect 9659 5956 9683 5958
rect 9739 5956 9763 5958
rect 9819 5956 9825 5958
rect 9517 5947 9825 5956
rect 9772 5772 9824 5778
rect 9876 5760 9904 6582
rect 9968 5778 9996 6598
rect 10152 5778 10180 8191
rect 10336 6118 10364 8191
rect 10428 7886 10456 8230
rect 10612 7954 10640 8434
rect 10980 8276 11008 8486
rect 11164 8294 11192 9386
rect 11532 9353 11560 9658
rect 11334 9344 11390 9353
rect 11334 9279 11390 9288
rect 11518 9344 11574 9353
rect 11518 9279 11574 9288
rect 11244 8968 11296 8974
rect 11242 8936 11244 8945
rect 11348 8956 11376 9279
rect 11296 8936 11376 8956
rect 11298 8928 11376 8936
rect 11242 8871 11298 8880
rect 11230 8732 11538 8741
rect 11230 8730 11236 8732
rect 11292 8730 11316 8732
rect 11372 8730 11396 8732
rect 11452 8730 11476 8732
rect 11532 8730 11538 8732
rect 11292 8678 11294 8730
rect 11474 8678 11476 8730
rect 11230 8676 11236 8678
rect 11292 8676 11316 8678
rect 11372 8676 11396 8678
rect 11452 8676 11476 8678
rect 11532 8676 11538 8678
rect 11230 8667 11538 8676
rect 11428 8492 11480 8498
rect 11428 8434 11480 8440
rect 11440 8362 11468 8434
rect 11624 8430 11652 10406
rect 11702 9888 11758 9897
rect 11702 9823 11758 9832
rect 11716 9450 11744 9823
rect 11794 9752 11850 9761
rect 11794 9687 11850 9696
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11808 9330 11836 9687
rect 11716 9302 11836 9330
rect 11716 9081 11744 9302
rect 11900 9160 11928 16594
rect 11992 16436 12020 17054
rect 12084 16794 12112 17546
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12176 17134 12204 17478
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12268 16561 12296 18414
rect 12070 16552 12126 16561
rect 12254 16552 12310 16561
rect 12126 16510 12204 16538
rect 12070 16487 12126 16496
rect 11992 16408 12112 16436
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11992 14958 12020 15506
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11992 13802 12020 14894
rect 12084 14414 12112 16408
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12176 14074 12204 16510
rect 12254 16487 12310 16496
rect 12360 16250 12388 19246
rect 12452 18086 12480 19314
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12544 17882 12572 22120
rect 12636 20942 12664 22188
rect 12624 20936 12676 20942
rect 12622 20904 12624 20913
rect 12676 20904 12678 20913
rect 12622 20839 12678 20848
rect 12728 20466 12756 23174
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12728 20058 12756 20266
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17202 12480 17682
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12346 15600 12402 15609
rect 12346 15535 12402 15544
rect 12360 15434 12388 15535
rect 12348 15428 12400 15434
rect 12348 15370 12400 15376
rect 12452 15201 12480 17138
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12438 15192 12494 15201
rect 12438 15127 12494 15136
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 14822 12388 14962
rect 12348 14816 12400 14822
rect 12544 14770 12572 17070
rect 12636 16658 12664 19110
rect 12714 19000 12770 19009
rect 12714 18935 12770 18944
rect 12728 18766 12756 18935
rect 12820 18873 12848 23054
rect 12944 22332 13252 22341
rect 12944 22330 12950 22332
rect 13006 22330 13030 22332
rect 13086 22330 13110 22332
rect 13166 22330 13190 22332
rect 13246 22330 13252 22332
rect 13006 22278 13008 22330
rect 13188 22278 13190 22330
rect 12944 22276 12950 22278
rect 13006 22276 13030 22278
rect 13086 22276 13110 22278
rect 13166 22276 13190 22278
rect 13246 22276 13252 22278
rect 12944 22267 13252 22276
rect 13176 22228 13228 22234
rect 13280 22216 13308 23462
rect 13372 23118 13400 23462
rect 13360 23112 13412 23118
rect 13452 23112 13504 23118
rect 13360 23054 13412 23060
rect 13450 23080 13452 23089
rect 13504 23080 13506 23089
rect 13450 23015 13506 23024
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13360 22500 13412 22506
rect 13360 22442 13412 22448
rect 13228 22188 13308 22216
rect 13176 22170 13228 22176
rect 12900 22024 12952 22030
rect 12900 21966 12952 21972
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 12912 21894 12940 21966
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 13004 21690 13032 21966
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13096 21554 13124 21830
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 12944 21244 13252 21253
rect 12944 21242 12950 21244
rect 13006 21242 13030 21244
rect 13086 21242 13110 21244
rect 13166 21242 13190 21244
rect 13246 21242 13252 21244
rect 13006 21190 13008 21242
rect 13188 21190 13190 21242
rect 12944 21188 12950 21190
rect 13006 21188 13030 21190
rect 13086 21188 13110 21190
rect 13166 21188 13190 21190
rect 13246 21188 13252 21190
rect 12944 21179 13252 21188
rect 13280 20466 13308 22188
rect 13372 22094 13400 22442
rect 13464 22273 13492 22578
rect 13450 22264 13506 22273
rect 13556 22234 13584 26030
rect 13648 25362 13676 26182
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 13740 25294 13768 26302
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13832 25401 13860 25638
rect 13818 25392 13874 25401
rect 13818 25327 13874 25336
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13820 25220 13872 25226
rect 13820 25162 13872 25168
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13740 24721 13768 24754
rect 13726 24712 13782 24721
rect 13726 24647 13782 24656
rect 13832 24290 13860 25162
rect 13636 24268 13688 24274
rect 13636 24210 13688 24216
rect 13740 24262 13860 24290
rect 13648 23254 13676 24210
rect 13740 24138 13768 24262
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13740 23322 13768 23734
rect 13728 23316 13780 23322
rect 13728 23258 13780 23264
rect 13636 23248 13688 23254
rect 13636 23190 13688 23196
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13648 22778 13676 23054
rect 13636 22772 13688 22778
rect 13636 22714 13688 22720
rect 13728 22636 13780 22642
rect 13728 22578 13780 22584
rect 13740 22409 13768 22578
rect 13726 22400 13782 22409
rect 13726 22335 13782 22344
rect 13832 22250 13860 24142
rect 13912 23044 13964 23050
rect 13912 22986 13964 22992
rect 13924 22642 13952 22986
rect 14108 22794 14136 27254
rect 14476 27146 14504 38694
rect 14657 38108 14965 38117
rect 14657 38106 14663 38108
rect 14719 38106 14743 38108
rect 14799 38106 14823 38108
rect 14879 38106 14903 38108
rect 14959 38106 14965 38108
rect 14719 38054 14721 38106
rect 14901 38054 14903 38106
rect 14657 38052 14663 38054
rect 14719 38052 14743 38054
rect 14799 38052 14823 38054
rect 14879 38052 14903 38054
rect 14959 38052 14965 38054
rect 14657 38043 14965 38052
rect 14657 37020 14965 37029
rect 14657 37018 14663 37020
rect 14719 37018 14743 37020
rect 14799 37018 14823 37020
rect 14879 37018 14903 37020
rect 14959 37018 14965 37020
rect 14719 36966 14721 37018
rect 14901 36966 14903 37018
rect 14657 36964 14663 36966
rect 14719 36964 14743 36966
rect 14799 36964 14823 36966
rect 14879 36964 14903 36966
rect 14959 36964 14965 36966
rect 14657 36955 14965 36964
rect 14657 35932 14965 35941
rect 14657 35930 14663 35932
rect 14719 35930 14743 35932
rect 14799 35930 14823 35932
rect 14879 35930 14903 35932
rect 14959 35930 14965 35932
rect 14719 35878 14721 35930
rect 14901 35878 14903 35930
rect 14657 35876 14663 35878
rect 14719 35876 14743 35878
rect 14799 35876 14823 35878
rect 14879 35876 14903 35878
rect 14959 35876 14965 35878
rect 14657 35867 14965 35876
rect 14657 34844 14965 34853
rect 14657 34842 14663 34844
rect 14719 34842 14743 34844
rect 14799 34842 14823 34844
rect 14879 34842 14903 34844
rect 14959 34842 14965 34844
rect 14719 34790 14721 34842
rect 14901 34790 14903 34842
rect 14657 34788 14663 34790
rect 14719 34788 14743 34790
rect 14799 34788 14823 34790
rect 14879 34788 14903 34790
rect 14959 34788 14965 34790
rect 14657 34779 14965 34788
rect 14657 33756 14965 33765
rect 14657 33754 14663 33756
rect 14719 33754 14743 33756
rect 14799 33754 14823 33756
rect 14879 33754 14903 33756
rect 14959 33754 14965 33756
rect 14719 33702 14721 33754
rect 14901 33702 14903 33754
rect 14657 33700 14663 33702
rect 14719 33700 14743 33702
rect 14799 33700 14823 33702
rect 14879 33700 14903 33702
rect 14959 33700 14965 33702
rect 14657 33691 14965 33700
rect 14657 32668 14965 32677
rect 14657 32666 14663 32668
rect 14719 32666 14743 32668
rect 14799 32666 14823 32668
rect 14879 32666 14903 32668
rect 14959 32666 14965 32668
rect 14719 32614 14721 32666
rect 14901 32614 14903 32666
rect 14657 32612 14663 32614
rect 14719 32612 14743 32614
rect 14799 32612 14823 32614
rect 14879 32612 14903 32614
rect 14959 32612 14965 32614
rect 14657 32603 14965 32612
rect 14657 31580 14965 31589
rect 14657 31578 14663 31580
rect 14719 31578 14743 31580
rect 14799 31578 14823 31580
rect 14879 31578 14903 31580
rect 14959 31578 14965 31580
rect 14719 31526 14721 31578
rect 14901 31526 14903 31578
rect 14657 31524 14663 31526
rect 14719 31524 14743 31526
rect 14799 31524 14823 31526
rect 14879 31524 14903 31526
rect 14959 31524 14965 31526
rect 14657 31515 14965 31524
rect 14556 30660 14608 30666
rect 14556 30602 14608 30608
rect 14568 28937 14596 30602
rect 14657 30492 14965 30501
rect 14657 30490 14663 30492
rect 14719 30490 14743 30492
rect 14799 30490 14823 30492
rect 14879 30490 14903 30492
rect 14959 30490 14965 30492
rect 14719 30438 14721 30490
rect 14901 30438 14903 30490
rect 14657 30436 14663 30438
rect 14719 30436 14743 30438
rect 14799 30436 14823 30438
rect 14879 30436 14903 30438
rect 14959 30436 14965 30438
rect 14657 30427 14965 30436
rect 14657 29404 14965 29413
rect 14657 29402 14663 29404
rect 14719 29402 14743 29404
rect 14799 29402 14823 29404
rect 14879 29402 14903 29404
rect 14959 29402 14965 29404
rect 14719 29350 14721 29402
rect 14901 29350 14903 29402
rect 14657 29348 14663 29350
rect 14719 29348 14743 29350
rect 14799 29348 14823 29350
rect 14879 29348 14903 29350
rect 14959 29348 14965 29350
rect 14657 29339 14965 29348
rect 14554 28928 14610 28937
rect 14554 28863 14610 28872
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14292 27118 14504 27146
rect 14292 24750 14320 27118
rect 14464 27056 14516 27062
rect 14464 26998 14516 27004
rect 14372 26240 14424 26246
rect 14372 26182 14424 26188
rect 14384 25265 14412 26182
rect 14370 25256 14426 25265
rect 14370 25191 14426 25200
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14188 24608 14240 24614
rect 14186 24576 14188 24585
rect 14240 24576 14242 24585
rect 14186 24511 14242 24520
rect 14384 24313 14412 25094
rect 14370 24304 14426 24313
rect 14370 24239 14426 24248
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23769 14412 24006
rect 14370 23760 14426 23769
rect 14370 23695 14426 23704
rect 14372 23520 14424 23526
rect 14370 23488 14372 23497
rect 14424 23488 14426 23497
rect 14370 23423 14426 23432
rect 14372 23248 14424 23254
rect 14370 23216 14372 23225
rect 14424 23216 14426 23225
rect 14370 23151 14426 23160
rect 14280 23112 14332 23118
rect 14280 23054 14332 23060
rect 14108 22766 14228 22794
rect 14292 22778 14320 23054
rect 14096 22704 14148 22710
rect 14096 22646 14148 22652
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 14004 22568 14056 22574
rect 13450 22199 13506 22208
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13648 22222 13860 22250
rect 13924 22516 14004 22522
rect 13924 22510 14056 22516
rect 13924 22494 14044 22510
rect 13372 22066 13492 22094
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13372 20602 13400 21490
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13360 20392 13412 20398
rect 13360 20334 13412 20340
rect 12944 20156 13252 20165
rect 12944 20154 12950 20156
rect 13006 20154 13030 20156
rect 13086 20154 13110 20156
rect 13166 20154 13190 20156
rect 13246 20154 13252 20156
rect 13006 20102 13008 20154
rect 13188 20102 13190 20154
rect 12944 20100 12950 20102
rect 13006 20100 13030 20102
rect 13086 20100 13110 20102
rect 13166 20100 13190 20102
rect 13246 20100 13252 20102
rect 12944 20091 13252 20100
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 12944 19068 13252 19077
rect 12944 19066 12950 19068
rect 13006 19066 13030 19068
rect 13086 19066 13110 19068
rect 13166 19066 13190 19068
rect 13246 19066 13252 19068
rect 13006 19014 13008 19066
rect 13188 19014 13190 19066
rect 12944 19012 12950 19014
rect 13006 19012 13030 19014
rect 13086 19012 13110 19014
rect 13166 19012 13190 19014
rect 13246 19012 13252 19014
rect 12944 19003 13252 19012
rect 12806 18864 12862 18873
rect 13280 18850 13308 19858
rect 12806 18799 12862 18808
rect 13096 18822 13308 18850
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 13096 18170 13124 18822
rect 13174 18728 13230 18737
rect 13174 18663 13230 18672
rect 13188 18290 13216 18663
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13174 18184 13230 18193
rect 13096 18142 13174 18170
rect 13174 18119 13230 18128
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12728 17202 12756 18022
rect 12820 17678 12848 18022
rect 12944 17980 13252 17989
rect 12944 17978 12950 17980
rect 13006 17978 13030 17980
rect 13086 17978 13110 17980
rect 13166 17978 13190 17980
rect 13246 17978 13252 17980
rect 13006 17926 13008 17978
rect 13188 17926 13190 17978
rect 12944 17924 12950 17926
rect 13006 17924 13030 17926
rect 13086 17924 13110 17926
rect 13166 17924 13190 17926
rect 13246 17924 13252 17926
rect 12944 17915 13252 17924
rect 12808 17672 12860 17678
rect 12808 17614 12860 17620
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 13096 17134 13124 17614
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 12944 16892 13252 16901
rect 12944 16890 12950 16892
rect 13006 16890 13030 16892
rect 13086 16890 13110 16892
rect 13166 16890 13190 16892
rect 13246 16890 13252 16892
rect 13006 16838 13008 16890
rect 13188 16838 13190 16890
rect 12944 16836 12950 16838
rect 13006 16836 13030 16838
rect 13086 16836 13110 16838
rect 13166 16836 13190 16838
rect 13246 16836 13252 16838
rect 12714 16824 12770 16833
rect 12944 16827 13252 16836
rect 12714 16759 12716 16768
rect 12768 16759 12770 16768
rect 12716 16730 12768 16736
rect 12990 16688 13046 16697
rect 12624 16652 12676 16658
rect 13046 16658 13124 16674
rect 13280 16658 13308 18566
rect 13372 18426 13400 20334
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13464 18358 13492 22066
rect 13648 21842 13676 22222
rect 13924 22094 13952 22494
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13832 22066 13952 22094
rect 13832 22012 13860 22066
rect 14016 22030 14044 22374
rect 14108 22098 14136 22646
rect 14096 22092 14148 22098
rect 14096 22034 14148 22040
rect 13912 22024 13964 22030
rect 13832 21984 13912 22012
rect 13912 21966 13964 21972
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14004 21888 14056 21894
rect 13648 21814 13952 21842
rect 14004 21830 14056 21836
rect 13820 21344 13872 21350
rect 13726 21312 13782 21321
rect 13820 21286 13872 21292
rect 13726 21247 13782 21256
rect 13542 21176 13598 21185
rect 13598 21134 13676 21162
rect 13542 21111 13598 21120
rect 13544 20800 13596 20806
rect 13544 20742 13596 20748
rect 13556 20466 13584 20742
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13648 20346 13676 21134
rect 13556 20318 13676 20346
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13452 18080 13504 18086
rect 13358 18048 13414 18057
rect 13452 18022 13504 18028
rect 13358 17983 13414 17992
rect 13372 17882 13400 17983
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13464 17762 13492 18022
rect 13372 17734 13492 17762
rect 13046 16652 13136 16658
rect 13046 16646 13084 16652
rect 12990 16623 13046 16632
rect 12624 16594 12676 16600
rect 13084 16594 13136 16600
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12714 16144 12770 16153
rect 12820 16114 12848 16390
rect 12348 14758 12400 14764
rect 12452 14742 12572 14770
rect 12636 16088 12714 16096
rect 12636 16068 12716 16088
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12268 13870 12296 14554
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11992 12782 12020 13738
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 11132 12020 12718
rect 12084 11558 12112 13262
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12072 11144 12124 11150
rect 11992 11104 12072 11132
rect 12072 11086 12124 11092
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 10441 12020 10542
rect 12084 10470 12112 11086
rect 12072 10464 12124 10470
rect 11978 10432 12034 10441
rect 12072 10406 12124 10412
rect 11978 10367 12034 10376
rect 12084 10266 12112 10406
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11978 10160 12034 10169
rect 12176 10146 12204 13262
rect 12268 12617 12296 13806
rect 12346 13288 12402 13297
rect 12346 13223 12402 13232
rect 12360 12918 12388 13223
rect 12452 12986 12480 14742
rect 12532 13864 12584 13870
rect 12530 13832 12532 13841
rect 12584 13832 12586 13841
rect 12530 13767 12586 13776
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12254 12608 12310 12617
rect 12254 12543 12310 12552
rect 12452 12322 12480 12922
rect 12544 12458 12572 13767
rect 12636 12900 12664 16068
rect 12768 16079 12770 16088
rect 12808 16108 12860 16114
rect 12716 16050 12768 16056
rect 12808 16050 12860 16056
rect 13004 15994 13032 16526
rect 13082 16280 13138 16289
rect 13082 16215 13138 16224
rect 12820 15978 13032 15994
rect 12808 15972 13032 15978
rect 12860 15966 13032 15972
rect 12808 15914 12860 15920
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12728 14929 12756 14962
rect 12714 14920 12770 14929
rect 12714 14855 12770 14864
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12728 13938 12756 14214
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12716 13388 12768 13394
rect 12716 13330 12768 13336
rect 12728 12986 12756 13330
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12634 12872 12664 12900
rect 12634 12832 12662 12872
rect 12634 12804 12756 12832
rect 12622 12472 12678 12481
rect 12544 12430 12622 12458
rect 12622 12407 12678 12416
rect 12256 12300 12308 12306
rect 12452 12294 12664 12322
rect 12256 12242 12308 12248
rect 12268 11354 12296 12242
rect 12636 12238 12664 12294
rect 12622 12232 12674 12238
rect 12622 12174 12674 12180
rect 12622 11792 12678 11801
rect 12348 11756 12400 11762
rect 12622 11727 12678 11736
rect 12348 11698 12400 11704
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12360 11257 12388 11698
rect 12346 11248 12402 11257
rect 12346 11183 12402 11192
rect 12636 11150 12664 11727
rect 12728 11626 12756 12804
rect 12820 12434 12848 15914
rect 13096 15910 13124 16215
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13084 15904 13136 15910
rect 13084 15846 13136 15852
rect 12944 15804 13252 15813
rect 12944 15802 12950 15804
rect 13006 15802 13030 15804
rect 13086 15802 13110 15804
rect 13166 15802 13190 15804
rect 13246 15802 13252 15804
rect 13006 15750 13008 15802
rect 13188 15750 13190 15802
rect 12944 15748 12950 15750
rect 13006 15748 13030 15750
rect 13086 15748 13110 15750
rect 13166 15748 13190 15750
rect 13246 15748 13252 15750
rect 12944 15739 13252 15748
rect 13280 15706 13308 15982
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 12898 15056 12954 15065
rect 12898 14991 12954 15000
rect 12912 14822 12940 14991
rect 12900 14816 12952 14822
rect 13188 14804 13216 15302
rect 13372 15162 13400 17734
rect 13556 17320 13584 20318
rect 13634 20224 13690 20233
rect 13634 20159 13690 20168
rect 13648 19836 13676 20159
rect 13740 20058 13768 21247
rect 13832 21049 13860 21286
rect 13818 21040 13874 21049
rect 13818 20975 13874 20984
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13648 19808 13768 19836
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13648 18902 13676 19382
rect 13636 18896 13688 18902
rect 13636 18838 13688 18844
rect 13740 17954 13768 19808
rect 13832 18358 13860 19926
rect 13924 18902 13952 21814
rect 14016 19990 14044 21830
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14108 20602 14136 21490
rect 14200 21486 14228 22766
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 14476 22556 14504 26998
rect 14292 22528 14504 22556
rect 14292 21842 14320 22528
rect 14462 22400 14518 22409
rect 14462 22335 14518 22344
rect 14476 22234 14504 22335
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14462 22128 14518 22137
rect 14462 22063 14518 22072
rect 14292 21814 14412 21842
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 14292 21593 14320 21626
rect 14278 21584 14334 21593
rect 14278 21519 14334 21528
rect 14188 21480 14240 21486
rect 14384 21468 14412 21814
rect 14476 21690 14504 22063
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14188 21422 14240 21428
rect 14292 21440 14412 21468
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14094 20496 14150 20505
rect 14094 20431 14150 20440
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 14004 19848 14056 19854
rect 14004 19790 14056 19796
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13912 18760 13964 18766
rect 13912 18702 13964 18708
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13464 17292 13584 17320
rect 13648 17926 13768 17954
rect 13648 17320 13676 17926
rect 13728 17808 13780 17814
rect 13780 17756 13860 17762
rect 13728 17750 13860 17756
rect 13740 17734 13860 17750
rect 13648 17292 13768 17320
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13188 14776 13308 14804
rect 12900 14758 12952 14764
rect 12944 14716 13252 14725
rect 12944 14714 12950 14716
rect 13006 14714 13030 14716
rect 13086 14714 13110 14716
rect 13166 14714 13190 14716
rect 13246 14714 13252 14716
rect 13006 14662 13008 14714
rect 13188 14662 13190 14714
rect 12944 14660 12950 14662
rect 13006 14660 13030 14662
rect 13086 14660 13110 14662
rect 13166 14660 13190 14662
rect 13246 14660 13252 14662
rect 12944 14651 13252 14660
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13188 13734 13216 14418
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 12944 13628 13252 13637
rect 12944 13626 12950 13628
rect 13006 13626 13030 13628
rect 13086 13626 13110 13628
rect 13166 13626 13190 13628
rect 13246 13626 13252 13628
rect 13006 13574 13008 13626
rect 13188 13574 13190 13626
rect 12944 13572 12950 13574
rect 13006 13572 13030 13574
rect 13086 13572 13110 13574
rect 13166 13572 13190 13574
rect 13246 13572 13252 13574
rect 12944 13563 13252 13572
rect 13280 13512 13308 14776
rect 13464 14278 13492 17292
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13556 16153 13584 17138
rect 13648 17105 13676 17138
rect 13634 17096 13690 17105
rect 13634 17031 13690 17040
rect 13542 16144 13598 16153
rect 13542 16079 13598 16088
rect 13636 16040 13688 16046
rect 13740 16028 13768 17292
rect 13832 16969 13860 17734
rect 13818 16960 13874 16969
rect 13818 16895 13874 16904
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16289 13860 16390
rect 13818 16280 13874 16289
rect 13818 16215 13874 16224
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13688 16000 13768 16028
rect 13636 15982 13688 15988
rect 13542 15328 13598 15337
rect 13542 15263 13598 15272
rect 13556 14550 13584 15263
rect 13648 14940 13676 15982
rect 13726 15872 13782 15881
rect 13726 15807 13782 15816
rect 13740 15094 13768 15807
rect 13832 15162 13860 16050
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13648 14912 13860 14940
rect 13634 14648 13690 14657
rect 13634 14583 13690 14592
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13004 13484 13308 13512
rect 13004 13394 13032 13484
rect 13082 13424 13138 13433
rect 12992 13388 13044 13394
rect 13138 13368 13216 13376
rect 13082 13359 13084 13368
rect 12992 13330 13044 13336
rect 13136 13348 13216 13368
rect 13084 13330 13136 13336
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 13096 12889 13124 13223
rect 13188 12918 13216 13348
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 13161 13308 13262
rect 13266 13152 13322 13161
rect 13266 13087 13322 13096
rect 13176 12912 13228 12918
rect 13082 12880 13138 12889
rect 13176 12854 13228 12860
rect 13082 12815 13138 12824
rect 12944 12540 13252 12549
rect 12944 12538 12950 12540
rect 13006 12538 13030 12540
rect 13086 12538 13110 12540
rect 13166 12538 13190 12540
rect 13246 12538 13252 12540
rect 13006 12486 13008 12538
rect 13188 12486 13190 12538
rect 12944 12484 12950 12486
rect 13006 12484 13030 12486
rect 13086 12484 13110 12486
rect 13166 12484 13190 12486
rect 13246 12484 13252 12486
rect 12944 12475 13252 12484
rect 12820 12406 12940 12434
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 11620 12768 11626
rect 12716 11562 12768 11568
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12728 11014 12756 11562
rect 12820 11354 12848 12174
rect 12912 11558 12940 12406
rect 13372 12306 13400 13670
rect 13556 13002 13584 14486
rect 13648 14482 13676 14583
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13648 14006 13676 14214
rect 13636 14000 13688 14006
rect 13636 13942 13688 13948
rect 13636 13864 13688 13870
rect 13728 13864 13780 13870
rect 13636 13806 13688 13812
rect 13726 13832 13728 13841
rect 13780 13832 13782 13841
rect 13648 13705 13676 13806
rect 13726 13767 13782 13776
rect 13634 13696 13690 13705
rect 13634 13631 13690 13640
rect 13556 12974 13676 13002
rect 13648 12866 13676 12974
rect 13648 12838 13768 12866
rect 13544 12708 13596 12714
rect 13544 12650 13596 12656
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13268 11620 13320 11626
rect 13268 11562 13320 11568
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12944 11452 13252 11461
rect 12944 11450 12950 11452
rect 13006 11450 13030 11452
rect 13086 11450 13110 11452
rect 13166 11450 13190 11452
rect 13246 11450 13252 11452
rect 13006 11398 13008 11450
rect 13188 11398 13190 11450
rect 12944 11396 12950 11398
rect 13006 11396 13030 11398
rect 13086 11396 13110 11398
rect 13166 11396 13190 11398
rect 13246 11396 13252 11398
rect 12944 11387 13252 11396
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 11978 10095 12034 10104
rect 12084 10118 12204 10146
rect 11992 9586 12020 10095
rect 12084 9636 12112 10118
rect 12268 10062 12296 10474
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12084 9608 12204 9636
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11808 9132 11928 9160
rect 11978 9208 12034 9217
rect 12084 9178 12112 9386
rect 11978 9143 12034 9152
rect 12072 9172 12124 9178
rect 11702 9072 11758 9081
rect 11702 9007 11758 9016
rect 11716 8820 11744 9007
rect 11808 8888 11836 9132
rect 11992 8974 12020 9143
rect 12072 9114 12124 9120
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11808 8860 11928 8888
rect 11716 8792 11836 8820
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11428 8356 11480 8362
rect 11428 8298 11480 8304
rect 11152 8288 11204 8294
rect 10980 8248 11100 8276
rect 10600 7948 10652 7954
rect 10652 7908 11008 7936
rect 10600 7890 10652 7896
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10598 7848 10654 7857
rect 10428 7206 10456 7822
rect 10598 7783 10654 7792
rect 10612 7478 10640 7783
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 9824 5732 9904 5760
rect 9956 5772 10008 5778
rect 9772 5714 9824 5720
rect 9956 5714 10008 5720
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 9784 5681 9812 5714
rect 9770 5672 9826 5681
rect 9770 5607 9826 5616
rect 10152 5370 10180 5714
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 9517 4924 9825 4933
rect 9517 4922 9523 4924
rect 9579 4922 9603 4924
rect 9659 4922 9683 4924
rect 9739 4922 9763 4924
rect 9819 4922 9825 4924
rect 9579 4870 9581 4922
rect 9761 4870 9763 4922
rect 9517 4868 9523 4870
rect 9579 4868 9603 4870
rect 9659 4868 9683 4870
rect 9739 4868 9763 4870
rect 9819 4868 9825 4870
rect 9517 4859 9825 4868
rect 10612 4214 10640 7414
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10704 6390 10732 6734
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10704 5778 10732 6326
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 10796 5166 10824 7346
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10888 5710 10916 6938
rect 10980 6866 11008 7908
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6322 11008 6802
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10980 5778 11008 6122
rect 10968 5772 11020 5778
rect 10968 5714 11020 5720
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10888 5250 10916 5646
rect 10966 5264 11022 5273
rect 10888 5222 10966 5250
rect 10966 5199 11022 5208
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 11072 4622 11100 8248
rect 11152 8230 11204 8236
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11244 8016 11296 8022
rect 11242 7984 11244 7993
rect 11296 7984 11298 7993
rect 11152 7948 11204 7954
rect 11242 7919 11298 7928
rect 11152 7890 11204 7896
rect 11164 6338 11192 7890
rect 11230 7644 11538 7653
rect 11230 7642 11236 7644
rect 11292 7642 11316 7644
rect 11372 7642 11396 7644
rect 11452 7642 11476 7644
rect 11532 7642 11538 7644
rect 11292 7590 11294 7642
rect 11474 7590 11476 7642
rect 11230 7588 11236 7590
rect 11292 7588 11316 7590
rect 11372 7588 11396 7590
rect 11452 7588 11476 7590
rect 11532 7588 11538 7590
rect 11230 7579 11538 7588
rect 11624 6866 11652 8230
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11230 6556 11538 6565
rect 11230 6554 11236 6556
rect 11292 6554 11316 6556
rect 11372 6554 11396 6556
rect 11452 6554 11476 6556
rect 11532 6554 11538 6556
rect 11292 6502 11294 6554
rect 11474 6502 11476 6554
rect 11230 6500 11236 6502
rect 11292 6500 11316 6502
rect 11372 6500 11396 6502
rect 11452 6500 11476 6502
rect 11532 6500 11538 6502
rect 11230 6491 11538 6500
rect 11164 6310 11284 6338
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11164 5914 11192 6054
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11256 5794 11284 6310
rect 11164 5766 11284 5794
rect 11164 4690 11192 5766
rect 11716 5574 11744 8366
rect 11808 8090 11836 8792
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11900 7546 11928 8860
rect 11978 8256 12034 8265
rect 12084 8242 12112 8910
rect 12034 8214 12112 8242
rect 11978 8191 12034 8200
rect 12072 7880 12124 7886
rect 11992 7840 12072 7868
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11808 5642 11836 6734
rect 11900 6089 11928 7278
rect 11992 6458 12020 7840
rect 12072 7822 12124 7828
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11886 6080 11942 6089
rect 11886 6015 11942 6024
rect 11886 5944 11942 5953
rect 11886 5879 11942 5888
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11230 5468 11538 5477
rect 11230 5466 11236 5468
rect 11292 5466 11316 5468
rect 11372 5466 11396 5468
rect 11452 5466 11476 5468
rect 11532 5466 11538 5468
rect 11292 5414 11294 5466
rect 11474 5414 11476 5466
rect 11230 5412 11236 5414
rect 11292 5412 11316 5414
rect 11372 5412 11396 5414
rect 11452 5412 11476 5414
rect 11532 5412 11538 5414
rect 11230 5403 11538 5412
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11230 4380 11538 4389
rect 11230 4378 11236 4380
rect 11292 4378 11316 4380
rect 11372 4378 11396 4380
rect 11452 4378 11476 4380
rect 11532 4378 11538 4380
rect 11292 4326 11294 4378
rect 11474 4326 11476 4378
rect 11230 4324 11236 4326
rect 11292 4324 11316 4326
rect 11372 4324 11396 4326
rect 11452 4324 11476 4326
rect 11532 4324 11538 4326
rect 11230 4315 11538 4324
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 11900 4146 11928 5879
rect 12084 5846 12112 6598
rect 12176 6497 12204 9608
rect 12254 9480 12310 9489
rect 12254 9415 12310 9424
rect 12268 7410 12296 9415
rect 12360 7546 12388 10950
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12438 10296 12494 10305
rect 12438 10231 12494 10240
rect 12452 9722 12480 10231
rect 12544 9761 12572 10610
rect 12530 9752 12586 9761
rect 12440 9716 12492 9722
rect 12530 9687 12586 9696
rect 12440 9658 12492 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 9042 12480 9318
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12544 8838 12572 9522
rect 12636 9432 12664 10746
rect 12944 10364 13252 10373
rect 12944 10362 12950 10364
rect 13006 10362 13030 10364
rect 13086 10362 13110 10364
rect 13166 10362 13190 10364
rect 13246 10362 13252 10364
rect 13006 10310 13008 10362
rect 13188 10310 13190 10362
rect 12944 10308 12950 10310
rect 13006 10308 13030 10310
rect 13086 10308 13110 10310
rect 13166 10308 13190 10310
rect 13246 10308 13252 10310
rect 12944 10299 13252 10308
rect 13280 10266 13308 11562
rect 13372 10266 13400 11834
rect 13464 11762 13492 12242
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13556 11694 13584 12650
rect 13740 12434 13768 12838
rect 13832 12714 13860 14912
rect 13924 13530 13952 18702
rect 14016 14618 14044 19790
rect 14108 19514 14136 20431
rect 14200 19854 14228 20742
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 17678 14136 18566
rect 14200 18086 14228 19654
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14292 17864 14320 21440
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14370 20224 14426 20233
rect 14370 20159 14426 20168
rect 14384 19514 14412 20159
rect 14476 19718 14504 20402
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14370 19136 14426 19145
rect 14370 19071 14426 19080
rect 14384 18426 14412 19071
rect 14476 18873 14504 19178
rect 14462 18864 14518 18873
rect 14462 18799 14518 18808
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14200 17836 14320 17864
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14094 17232 14150 17241
rect 14094 17167 14150 17176
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14002 13696 14058 13705
rect 14002 13631 14058 13640
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13910 13424 13966 13433
rect 13910 13359 13966 13368
rect 13924 12850 13952 13359
rect 14016 12850 14044 13631
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13910 12744 13966 12753
rect 13820 12708 13872 12714
rect 13910 12679 13966 12688
rect 13820 12650 13872 12656
rect 13648 12406 13768 12434
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13452 11552 13504 11558
rect 13452 11494 13504 11500
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 12714 10160 12770 10169
rect 13464 10146 13492 11494
rect 13556 11286 13584 11630
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 12770 10118 12848 10146
rect 12714 10095 12770 10104
rect 12716 9648 12768 9654
rect 12714 9616 12716 9625
rect 12768 9616 12770 9625
rect 12714 9551 12770 9560
rect 12820 9518 12848 10118
rect 13372 10118 13492 10146
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 12808 9512 12860 9518
rect 13280 9489 13308 9862
rect 12808 9454 12860 9460
rect 13266 9480 13322 9489
rect 12636 9404 12756 9432
rect 12622 9208 12678 9217
rect 12622 9143 12678 9152
rect 12532 8832 12584 8838
rect 12438 8800 12494 8809
rect 12532 8774 12584 8780
rect 12438 8735 12494 8744
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12162 6488 12218 6497
rect 12162 6423 12218 6432
rect 12176 6390 12204 6423
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12268 5846 12296 6802
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 12256 5840 12308 5846
rect 12256 5782 12308 5788
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 11992 4826 12020 5714
rect 12070 5128 12126 5137
rect 12070 5063 12072 5072
rect 12124 5063 12126 5072
rect 12072 5034 12124 5040
rect 12084 4826 12112 5034
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9517 3836 9825 3845
rect 9517 3834 9523 3836
rect 9579 3834 9603 3836
rect 9659 3834 9683 3836
rect 9739 3834 9763 3836
rect 9819 3834 9825 3836
rect 9579 3782 9581 3834
rect 9761 3782 9763 3834
rect 9517 3780 9523 3782
rect 9579 3780 9603 3782
rect 9659 3780 9683 3782
rect 9739 3780 9763 3782
rect 9819 3780 9825 3782
rect 9517 3771 9825 3780
rect 11164 3534 11192 4082
rect 12084 3942 12112 4762
rect 12360 3942 12388 6190
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12084 3602 12112 3878
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11230 3292 11538 3301
rect 11230 3290 11236 3292
rect 11292 3290 11316 3292
rect 11372 3290 11396 3292
rect 11452 3290 11476 3292
rect 11532 3290 11538 3292
rect 11292 3238 11294 3290
rect 11474 3238 11476 3290
rect 11230 3236 11236 3238
rect 11292 3236 11316 3238
rect 11372 3236 11396 3238
rect 11452 3236 11476 3238
rect 11532 3236 11538 3238
rect 11230 3227 11538 3236
rect 9517 2748 9825 2757
rect 9517 2746 9523 2748
rect 9579 2746 9603 2748
rect 9659 2746 9683 2748
rect 9739 2746 9763 2748
rect 9819 2746 9825 2748
rect 9579 2694 9581 2746
rect 9761 2694 9763 2746
rect 9517 2692 9523 2694
rect 9579 2692 9603 2694
rect 9659 2692 9683 2694
rect 9739 2692 9763 2694
rect 9819 2692 9825 2694
rect 9517 2683 9825 2692
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 10888 2106 10916 2615
rect 11230 2204 11538 2213
rect 11230 2202 11236 2204
rect 11292 2202 11316 2204
rect 11372 2202 11396 2204
rect 11452 2202 11476 2204
rect 11532 2202 11538 2204
rect 11292 2150 11294 2202
rect 11474 2150 11476 2202
rect 11230 2148 11236 2150
rect 11292 2148 11316 2150
rect 11372 2148 11396 2150
rect 11452 2148 11476 2150
rect 11532 2148 11538 2150
rect 11230 2139 11538 2148
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 12084 2038 12112 3538
rect 12452 2106 12480 8735
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12544 8498 12572 8599
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 7936 12664 9143
rect 12728 8634 12756 9404
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12728 8090 12756 8366
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12716 7948 12768 7954
rect 12636 7908 12716 7936
rect 12716 7890 12768 7896
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 6730 12572 7142
rect 12532 6724 12584 6730
rect 12532 6666 12584 6672
rect 12544 5030 12572 6666
rect 12636 5760 12664 7686
rect 12820 7410 12848 9454
rect 13266 9415 13322 9424
rect 12944 9276 13252 9285
rect 12944 9274 12950 9276
rect 13006 9274 13030 9276
rect 13086 9274 13110 9276
rect 13166 9274 13190 9276
rect 13246 9274 13252 9276
rect 13006 9222 13008 9274
rect 13188 9222 13190 9274
rect 12944 9220 12950 9222
rect 13006 9220 13030 9222
rect 13086 9220 13110 9222
rect 13166 9220 13190 9222
rect 13246 9220 13252 9222
rect 12944 9211 13252 9220
rect 12992 9104 13044 9110
rect 13372 9058 13400 10118
rect 13450 10024 13506 10033
rect 13450 9959 13506 9968
rect 12992 9046 13044 9052
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 8294 12940 8842
rect 13004 8537 13032 9046
rect 13280 9030 13400 9058
rect 12990 8528 13046 8537
rect 12990 8463 13046 8472
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12944 8188 13252 8197
rect 12944 8186 12950 8188
rect 13006 8186 13030 8188
rect 13086 8186 13110 8188
rect 13166 8186 13190 8188
rect 13246 8186 13252 8188
rect 13006 8134 13008 8186
rect 13188 8134 13190 8186
rect 12944 8132 12950 8134
rect 13006 8132 13030 8134
rect 13086 8132 13110 8134
rect 13166 8132 13190 8134
rect 13246 8132 13252 8134
rect 12944 8123 13252 8132
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 12912 7857 12940 7958
rect 12898 7848 12954 7857
rect 12898 7783 12954 7792
rect 12900 7744 12952 7750
rect 13280 7732 13308 9030
rect 13360 8968 13412 8974
rect 13358 8936 13360 8945
rect 13412 8936 13414 8945
rect 13358 8871 13414 8880
rect 13464 8838 13492 9959
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13556 9586 13584 9658
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13556 8634 13584 9522
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 7993 13400 8230
rect 13358 7984 13414 7993
rect 13358 7919 13414 7928
rect 12952 7704 13308 7732
rect 12900 7686 12952 7692
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12716 7336 12768 7342
rect 12912 7290 12940 7686
rect 13556 7562 13584 8366
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13464 7534 13584 7562
rect 12716 7278 12768 7284
rect 12728 6730 12756 7278
rect 12820 7262 12940 7290
rect 12820 6798 12848 7262
rect 12944 7100 13252 7109
rect 12944 7098 12950 7100
rect 13006 7098 13030 7100
rect 13086 7098 13110 7100
rect 13166 7098 13190 7100
rect 13246 7098 13252 7100
rect 13006 7046 13008 7098
rect 13188 7046 13190 7098
rect 12944 7044 12950 7046
rect 13006 7044 13030 7046
rect 13086 7044 13110 7046
rect 13166 7044 13190 7046
rect 13246 7044 13252 7046
rect 12944 7035 13252 7044
rect 13280 6984 13308 7482
rect 13188 6956 13308 6984
rect 12898 6896 12954 6905
rect 12898 6831 12954 6840
rect 12912 6798 12940 6831
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12990 6488 13046 6497
rect 13188 6458 13216 6956
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 12990 6423 13046 6432
rect 13176 6452 13228 6458
rect 13004 6322 13032 6423
rect 13176 6394 13228 6400
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12714 6080 12770 6089
rect 12820 6066 12848 6258
rect 12770 6038 12848 6066
rect 12714 6015 12770 6024
rect 12944 6012 13252 6021
rect 12944 6010 12950 6012
rect 13006 6010 13030 6012
rect 13086 6010 13110 6012
rect 13166 6010 13190 6012
rect 13246 6010 13252 6012
rect 13006 5958 13008 6010
rect 13188 5958 13190 6010
rect 12944 5956 12950 5958
rect 13006 5956 13030 5958
rect 13086 5956 13110 5958
rect 13166 5956 13190 5958
rect 13246 5956 13252 5958
rect 12944 5947 13252 5956
rect 12716 5772 12768 5778
rect 12636 5732 12716 5760
rect 12716 5714 12768 5720
rect 12900 5704 12952 5710
rect 12622 5672 12678 5681
rect 12900 5646 12952 5652
rect 12622 5607 12678 5616
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12636 4554 12664 5607
rect 12912 5114 12940 5646
rect 12820 5086 12940 5114
rect 12716 4820 12768 4826
rect 12820 4808 12848 5086
rect 12944 4924 13252 4933
rect 12944 4922 12950 4924
rect 13006 4922 13030 4924
rect 13086 4922 13110 4924
rect 13166 4922 13190 4924
rect 13246 4922 13252 4924
rect 13006 4870 13008 4922
rect 13188 4870 13190 4922
rect 12944 4868 12950 4870
rect 13006 4868 13030 4870
rect 13086 4868 13110 4870
rect 13166 4868 13190 4870
rect 13246 4868 13252 4870
rect 12944 4859 13252 4868
rect 12768 4780 12848 4808
rect 12716 4762 12768 4768
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12636 4282 12664 4490
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 12072 2032 12124 2038
rect 12072 1974 12124 1980
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 10048 1964 10100 1970
rect 10048 1906 10100 1912
rect 10784 1964 10836 1970
rect 10784 1906 10836 1912
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 12256 1964 12308 1970
rect 12256 1906 12308 1912
rect 8588 1562 8616 1906
rect 9324 1562 9352 1906
rect 9517 1660 9825 1669
rect 9517 1658 9523 1660
rect 9579 1658 9603 1660
rect 9659 1658 9683 1660
rect 9739 1658 9763 1660
rect 9819 1658 9825 1660
rect 9579 1606 9581 1658
rect 9761 1606 9763 1658
rect 9517 1604 9523 1606
rect 9579 1604 9603 1606
rect 9659 1604 9683 1606
rect 9739 1604 9763 1606
rect 9819 1604 9825 1606
rect 9517 1595 9825 1604
rect 10060 1562 10088 1906
rect 10796 1562 10824 1906
rect 11624 1562 11652 1906
rect 11702 1864 11758 1873
rect 11702 1799 11758 1808
rect 11716 1766 11744 1799
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 12268 1562 12296 1906
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10784 1556 10836 1562
rect 10784 1498 10836 1504
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 11612 1352 11664 1358
rect 11612 1294 11664 1300
rect 12348 1352 12400 1358
rect 12348 1294 12400 1300
rect 8392 1012 8444 1018
rect 8392 954 8444 960
rect 8680 160 8708 1294
rect 9416 190 9536 218
rect 9416 160 9444 190
rect 7930 54 8248 82
rect 7194 0 7250 54
rect 7930 0 7986 54
rect 8666 0 8722 160
rect 9402 0 9458 160
rect 9508 82 9536 190
rect 9692 82 9720 1294
rect 9508 54 9720 82
rect 10138 82 10194 160
rect 10428 82 10456 1294
rect 10888 160 10916 1294
rect 11230 1116 11538 1125
rect 11230 1114 11236 1116
rect 11292 1114 11316 1116
rect 11372 1114 11396 1116
rect 11452 1114 11476 1116
rect 11532 1114 11538 1116
rect 11292 1062 11294 1114
rect 11474 1062 11476 1114
rect 11230 1060 11236 1062
rect 11292 1060 11316 1062
rect 11372 1060 11396 1062
rect 11452 1060 11476 1062
rect 11532 1060 11538 1062
rect 11230 1051 11538 1060
rect 11624 160 11652 1294
rect 12360 160 12388 1294
rect 12544 1290 12572 4014
rect 12944 3836 13252 3845
rect 12944 3834 12950 3836
rect 13006 3834 13030 3836
rect 13086 3834 13110 3836
rect 13166 3834 13190 3836
rect 13246 3834 13252 3836
rect 13006 3782 13008 3834
rect 13188 3782 13190 3834
rect 12944 3780 12950 3782
rect 13006 3780 13030 3782
rect 13086 3780 13110 3782
rect 13166 3780 13190 3782
rect 13246 3780 13252 3782
rect 12944 3771 13252 3780
rect 13280 3738 13308 6326
rect 13372 5370 13400 6802
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 13464 2774 13492 7534
rect 13544 7404 13596 7410
rect 13648 7392 13676 12406
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13740 10810 13768 11630
rect 13832 11218 13860 12038
rect 13924 11354 13952 12679
rect 14002 12472 14058 12481
rect 14108 12442 14136 17167
rect 14200 16726 14228 17836
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 14292 17241 14320 17682
rect 14278 17232 14334 17241
rect 14278 17167 14334 17176
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14278 16688 14334 16697
rect 14278 16623 14334 16632
rect 14292 16590 14320 16623
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14278 15056 14334 15065
rect 14188 15020 14240 15026
rect 14278 14991 14334 15000
rect 14188 14962 14240 14968
rect 14200 14521 14228 14962
rect 14186 14512 14242 14521
rect 14186 14447 14242 14456
rect 14292 14346 14320 14991
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14278 13832 14334 13841
rect 14278 13767 14334 13776
rect 14186 13560 14242 13569
rect 14186 13495 14242 13504
rect 14200 13025 14228 13495
rect 14186 13016 14242 13025
rect 14186 12951 14242 12960
rect 14200 12782 14228 12951
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14002 12407 14058 12416
rect 14096 12436 14148 12442
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13924 10266 13952 10950
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13820 10192 13872 10198
rect 13726 10160 13782 10169
rect 13820 10134 13872 10140
rect 13726 10095 13782 10104
rect 13740 8498 13768 10095
rect 13832 9586 13860 10134
rect 13910 9888 13966 9897
rect 13910 9823 13966 9832
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13818 9480 13874 9489
rect 13818 9415 13874 9424
rect 13832 9382 13860 9415
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13924 8537 13952 9823
rect 13910 8528 13966 8537
rect 13728 8492 13780 8498
rect 13910 8463 13966 8472
rect 13728 8434 13780 8440
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13740 7410 13768 8191
rect 13596 7364 13676 7392
rect 13728 7404 13780 7410
rect 13544 7346 13596 7352
rect 13728 7346 13780 7352
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13556 5914 13584 6287
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13648 4826 13676 6831
rect 13726 6352 13782 6361
rect 13726 6287 13782 6296
rect 13740 5234 13768 6287
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13832 3942 13860 7278
rect 14016 6798 14044 12407
rect 14096 12378 14148 12384
rect 14292 12238 14320 13767
rect 14384 13530 14412 18226
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14476 13410 14504 18634
rect 14384 13382 14504 13410
rect 14280 12232 14332 12238
rect 14280 12174 14332 12180
rect 14094 11792 14150 11801
rect 14094 11727 14150 11736
rect 14108 11150 14136 11727
rect 14278 11520 14334 11529
rect 14278 11455 14334 11464
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14188 10736 14240 10742
rect 14186 10704 14188 10713
rect 14240 10704 14242 10713
rect 14186 10639 14242 10648
rect 14094 10568 14150 10577
rect 14094 10503 14150 10512
rect 14108 10266 14136 10503
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14108 8430 14136 9658
rect 14292 8974 14320 11455
rect 14384 9654 14412 13382
rect 14464 13252 14516 13258
rect 14464 13194 14516 13200
rect 14476 12986 14504 13194
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14462 9344 14518 9353
rect 14462 9279 14518 9288
rect 14370 9072 14426 9081
rect 14476 9042 14504 9279
rect 14370 9007 14372 9016
rect 14424 9007 14426 9016
rect 14464 9036 14516 9042
rect 14372 8978 14424 8984
rect 14464 8978 14516 8984
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14292 8265 14320 8434
rect 14278 8256 14334 8265
rect 14278 8191 14334 8200
rect 14278 7984 14334 7993
rect 14568 7970 14596 28494
rect 14657 28316 14965 28325
rect 14657 28314 14663 28316
rect 14719 28314 14743 28316
rect 14799 28314 14823 28316
rect 14879 28314 14903 28316
rect 14959 28314 14965 28316
rect 14719 28262 14721 28314
rect 14901 28262 14903 28314
rect 14657 28260 14663 28262
rect 14719 28260 14743 28262
rect 14799 28260 14823 28262
rect 14879 28260 14903 28262
rect 14959 28260 14965 28262
rect 14657 28251 14965 28260
rect 14657 27228 14965 27237
rect 14657 27226 14663 27228
rect 14719 27226 14743 27228
rect 14799 27226 14823 27228
rect 14879 27226 14903 27228
rect 14959 27226 14965 27228
rect 14719 27174 14721 27226
rect 14901 27174 14903 27226
rect 14657 27172 14663 27174
rect 14719 27172 14743 27174
rect 14799 27172 14823 27174
rect 14879 27172 14903 27174
rect 14959 27172 14965 27174
rect 14657 27163 14965 27172
rect 14924 27124 14976 27130
rect 14924 27066 14976 27072
rect 14936 26489 14964 27066
rect 14922 26480 14978 26489
rect 14922 26415 14978 26424
rect 14657 26140 14965 26149
rect 14657 26138 14663 26140
rect 14719 26138 14743 26140
rect 14799 26138 14823 26140
rect 14879 26138 14903 26140
rect 14959 26138 14965 26140
rect 14719 26086 14721 26138
rect 14901 26086 14903 26138
rect 14657 26084 14663 26086
rect 14719 26084 14743 26086
rect 14799 26084 14823 26086
rect 14879 26084 14903 26086
rect 14959 26084 14965 26086
rect 14657 26075 14965 26084
rect 14657 25052 14965 25061
rect 14657 25050 14663 25052
rect 14719 25050 14743 25052
rect 14799 25050 14823 25052
rect 14879 25050 14903 25052
rect 14959 25050 14965 25052
rect 14719 24998 14721 25050
rect 14901 24998 14903 25050
rect 14657 24996 14663 24998
rect 14719 24996 14743 24998
rect 14799 24996 14823 24998
rect 14879 24996 14903 24998
rect 14959 24996 14965 24998
rect 14657 24987 14965 24996
rect 14657 23964 14965 23973
rect 14657 23962 14663 23964
rect 14719 23962 14743 23964
rect 14799 23962 14823 23964
rect 14879 23962 14903 23964
rect 14959 23962 14965 23964
rect 14719 23910 14721 23962
rect 14901 23910 14903 23962
rect 14657 23908 14663 23910
rect 14719 23908 14743 23910
rect 14799 23908 14823 23910
rect 14879 23908 14903 23910
rect 14959 23908 14965 23910
rect 14657 23899 14965 23908
rect 14657 22876 14965 22885
rect 14657 22874 14663 22876
rect 14719 22874 14743 22876
rect 14799 22874 14823 22876
rect 14879 22874 14903 22876
rect 14959 22874 14965 22876
rect 14719 22822 14721 22874
rect 14901 22822 14903 22874
rect 14657 22820 14663 22822
rect 14719 22820 14743 22822
rect 14799 22820 14823 22822
rect 14879 22820 14903 22822
rect 14959 22820 14965 22822
rect 14657 22811 14965 22820
rect 14924 22432 14976 22438
rect 14922 22400 14924 22409
rect 14976 22400 14978 22409
rect 14922 22335 14978 22344
rect 14657 21788 14965 21797
rect 14657 21786 14663 21788
rect 14719 21786 14743 21788
rect 14799 21786 14823 21788
rect 14879 21786 14903 21788
rect 14959 21786 14965 21788
rect 14719 21734 14721 21786
rect 14901 21734 14903 21786
rect 14657 21732 14663 21734
rect 14719 21732 14743 21734
rect 14799 21732 14823 21734
rect 14879 21732 14903 21734
rect 14959 21732 14965 21734
rect 14657 21723 14965 21732
rect 14657 20700 14965 20709
rect 14657 20698 14663 20700
rect 14719 20698 14743 20700
rect 14799 20698 14823 20700
rect 14879 20698 14903 20700
rect 14959 20698 14965 20700
rect 14719 20646 14721 20698
rect 14901 20646 14903 20698
rect 14657 20644 14663 20646
rect 14719 20644 14743 20646
rect 14799 20644 14823 20646
rect 14879 20644 14903 20646
rect 14959 20644 14965 20646
rect 14657 20635 14965 20644
rect 14646 19816 14702 19825
rect 14646 19751 14648 19760
rect 14700 19751 14702 19760
rect 14648 19722 14700 19728
rect 14657 19612 14965 19621
rect 14657 19610 14663 19612
rect 14719 19610 14743 19612
rect 14799 19610 14823 19612
rect 14879 19610 14903 19612
rect 14959 19610 14965 19612
rect 14719 19558 14721 19610
rect 14901 19558 14903 19610
rect 14657 19556 14663 19558
rect 14719 19556 14743 19558
rect 14799 19556 14823 19558
rect 14879 19556 14903 19558
rect 14959 19556 14965 19558
rect 14657 19547 14965 19556
rect 14657 18524 14965 18533
rect 14657 18522 14663 18524
rect 14719 18522 14743 18524
rect 14799 18522 14823 18524
rect 14879 18522 14903 18524
rect 14959 18522 14965 18524
rect 14719 18470 14721 18522
rect 14901 18470 14903 18522
rect 14657 18468 14663 18470
rect 14719 18468 14743 18470
rect 14799 18468 14823 18470
rect 14879 18468 14903 18470
rect 14959 18468 14965 18470
rect 14657 18459 14965 18468
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14660 17610 14688 18362
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14657 17436 14965 17445
rect 14657 17434 14663 17436
rect 14719 17434 14743 17436
rect 14799 17434 14823 17436
rect 14879 17434 14903 17436
rect 14959 17434 14965 17436
rect 14719 17382 14721 17434
rect 14901 17382 14903 17434
rect 14657 17380 14663 17382
rect 14719 17380 14743 17382
rect 14799 17380 14823 17382
rect 14879 17380 14903 17382
rect 14959 17380 14965 17382
rect 14657 17371 14965 17380
rect 14657 16348 14965 16357
rect 14657 16346 14663 16348
rect 14719 16346 14743 16348
rect 14799 16346 14823 16348
rect 14879 16346 14903 16348
rect 14959 16346 14965 16348
rect 14719 16294 14721 16346
rect 14901 16294 14903 16346
rect 14657 16292 14663 16294
rect 14719 16292 14743 16294
rect 14799 16292 14823 16294
rect 14879 16292 14903 16294
rect 14959 16292 14965 16294
rect 14657 16283 14965 16292
rect 14830 15600 14886 15609
rect 14830 15535 14886 15544
rect 14844 15502 14872 15535
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14657 15260 14965 15269
rect 14657 15258 14663 15260
rect 14719 15258 14743 15260
rect 14799 15258 14823 15260
rect 14879 15258 14903 15260
rect 14959 15258 14965 15260
rect 14719 15206 14721 15258
rect 14901 15206 14903 15258
rect 14657 15204 14663 15206
rect 14719 15204 14743 15206
rect 14799 15204 14823 15206
rect 14879 15204 14903 15206
rect 14959 15204 14965 15206
rect 14657 15195 14965 15204
rect 14830 14784 14886 14793
rect 14830 14719 14886 14728
rect 14844 14414 14872 14719
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14657 14172 14965 14181
rect 14657 14170 14663 14172
rect 14719 14170 14743 14172
rect 14799 14170 14823 14172
rect 14879 14170 14903 14172
rect 14959 14170 14965 14172
rect 14719 14118 14721 14170
rect 14901 14118 14903 14170
rect 14657 14116 14663 14118
rect 14719 14116 14743 14118
rect 14799 14116 14823 14118
rect 14879 14116 14903 14118
rect 14959 14116 14965 14118
rect 14657 14107 14965 14116
rect 14657 13084 14965 13093
rect 14657 13082 14663 13084
rect 14719 13082 14743 13084
rect 14799 13082 14823 13084
rect 14879 13082 14903 13084
rect 14959 13082 14965 13084
rect 14719 13030 14721 13082
rect 14901 13030 14903 13082
rect 14657 13028 14663 13030
rect 14719 13028 14743 13030
rect 14799 13028 14823 13030
rect 14879 13028 14903 13030
rect 14959 13028 14965 13030
rect 14657 13019 14965 13028
rect 14657 11996 14965 12005
rect 14657 11994 14663 11996
rect 14719 11994 14743 11996
rect 14799 11994 14823 11996
rect 14879 11994 14903 11996
rect 14959 11994 14965 11996
rect 14719 11942 14721 11994
rect 14901 11942 14903 11994
rect 14657 11940 14663 11942
rect 14719 11940 14743 11942
rect 14799 11940 14823 11942
rect 14879 11940 14903 11942
rect 14959 11940 14965 11942
rect 14657 11931 14965 11940
rect 14657 10908 14965 10917
rect 14657 10906 14663 10908
rect 14719 10906 14743 10908
rect 14799 10906 14823 10908
rect 14879 10906 14903 10908
rect 14959 10906 14965 10908
rect 14719 10854 14721 10906
rect 14901 10854 14903 10906
rect 14657 10852 14663 10854
rect 14719 10852 14743 10854
rect 14799 10852 14823 10854
rect 14879 10852 14903 10854
rect 14959 10852 14965 10854
rect 14657 10843 14965 10852
rect 14646 10432 14702 10441
rect 14646 10367 14702 10376
rect 14660 10130 14688 10367
rect 14648 10124 14700 10130
rect 14648 10066 14700 10072
rect 14657 9820 14965 9829
rect 14657 9818 14663 9820
rect 14719 9818 14743 9820
rect 14799 9818 14823 9820
rect 14879 9818 14903 9820
rect 14959 9818 14965 9820
rect 14719 9766 14721 9818
rect 14901 9766 14903 9818
rect 14657 9764 14663 9766
rect 14719 9764 14743 9766
rect 14799 9764 14823 9766
rect 14879 9764 14903 9766
rect 14959 9764 14965 9766
rect 14657 9755 14965 9764
rect 14657 8732 14965 8741
rect 14657 8730 14663 8732
rect 14719 8730 14743 8732
rect 14799 8730 14823 8732
rect 14879 8730 14903 8732
rect 14959 8730 14965 8732
rect 14719 8678 14721 8730
rect 14901 8678 14903 8730
rect 14657 8676 14663 8678
rect 14719 8676 14743 8678
rect 14799 8676 14823 8678
rect 14879 8676 14903 8678
rect 14959 8676 14965 8678
rect 14657 8667 14965 8676
rect 14278 7919 14334 7928
rect 14476 7942 14596 7970
rect 14292 7886 14320 7919
rect 14188 7880 14240 7886
rect 14186 7848 14188 7857
rect 14280 7880 14332 7886
rect 14240 7848 14242 7857
rect 14280 7822 14332 7828
rect 14186 7783 14242 7792
rect 14372 7200 14424 7206
rect 14278 7168 14334 7177
rect 14372 7142 14424 7148
rect 14278 7103 14334 7112
rect 14292 6798 14320 7103
rect 14384 7002 14412 7142
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14004 6792 14056 6798
rect 13910 6760 13966 6769
rect 14004 6734 14056 6740
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 13910 6695 13966 6704
rect 13924 6662 13952 6695
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13924 5545 13952 6258
rect 13910 5536 13966 5545
rect 13910 5471 13966 5480
rect 13924 4826 13952 5471
rect 14016 5273 14044 6734
rect 14476 6458 14504 7942
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14568 7449 14596 7754
rect 14657 7644 14965 7653
rect 14657 7642 14663 7644
rect 14719 7642 14743 7644
rect 14799 7642 14823 7644
rect 14879 7642 14903 7644
rect 14959 7642 14965 7644
rect 14719 7590 14721 7642
rect 14901 7590 14903 7642
rect 14657 7588 14663 7590
rect 14719 7588 14743 7590
rect 14799 7588 14823 7590
rect 14879 7588 14903 7590
rect 14959 7588 14965 7590
rect 14657 7579 14965 7588
rect 14554 7440 14610 7449
rect 14554 7375 14610 7384
rect 14657 6556 14965 6565
rect 14657 6554 14663 6556
rect 14719 6554 14743 6556
rect 14799 6554 14823 6556
rect 14879 6554 14903 6556
rect 14959 6554 14965 6556
rect 14719 6502 14721 6554
rect 14901 6502 14903 6554
rect 14657 6500 14663 6502
rect 14719 6500 14743 6502
rect 14799 6500 14823 6502
rect 14879 6500 14903 6502
rect 14959 6500 14965 6502
rect 14657 6491 14965 6500
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14370 6216 14426 6225
rect 14370 6151 14426 6160
rect 14384 5914 14412 6151
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14830 5808 14886 5817
rect 14830 5743 14886 5752
rect 14844 5710 14872 5743
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14292 5545 14320 5578
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14657 5468 14965 5477
rect 14657 5466 14663 5468
rect 14719 5466 14743 5468
rect 14799 5466 14823 5468
rect 14879 5466 14903 5468
rect 14959 5466 14965 5468
rect 14719 5414 14721 5466
rect 14901 5414 14903 5466
rect 14657 5412 14663 5414
rect 14719 5412 14743 5414
rect 14799 5412 14823 5414
rect 14879 5412 14903 5414
rect 14959 5412 14965 5414
rect 14657 5403 14965 5412
rect 14002 5264 14058 5273
rect 14002 5199 14004 5208
rect 14056 5199 14058 5208
rect 14004 5170 14056 5176
rect 14278 4992 14334 5001
rect 14278 4927 14334 4936
rect 13912 4820 13964 4826
rect 13912 4762 13964 4768
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 14292 3534 14320 4927
rect 14657 4380 14965 4389
rect 14657 4378 14663 4380
rect 14719 4378 14743 4380
rect 14799 4378 14823 4380
rect 14879 4378 14903 4380
rect 14959 4378 14965 4380
rect 14719 4326 14721 4378
rect 14901 4326 14903 4378
rect 14657 4324 14663 4326
rect 14719 4324 14743 4326
rect 14799 4324 14823 4326
rect 14879 4324 14903 4326
rect 14959 4324 14965 4326
rect 14657 4315 14965 4324
rect 14370 4040 14426 4049
rect 14370 3975 14426 3984
rect 14384 3738 14412 3975
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14657 3292 14965 3301
rect 14657 3290 14663 3292
rect 14719 3290 14743 3292
rect 14799 3290 14823 3292
rect 14879 3290 14903 3292
rect 14959 3290 14965 3292
rect 14719 3238 14721 3290
rect 14901 3238 14903 3290
rect 14657 3236 14663 3238
rect 14719 3236 14743 3238
rect 14799 3236 14823 3238
rect 14879 3236 14903 3238
rect 14959 3236 14965 3238
rect 14657 3227 14965 3236
rect 12944 2748 13252 2757
rect 12944 2746 12950 2748
rect 13006 2746 13030 2748
rect 13086 2746 13110 2748
rect 13166 2746 13190 2748
rect 13246 2746 13252 2748
rect 13006 2694 13008 2746
rect 13188 2694 13190 2746
rect 12944 2692 12950 2694
rect 13006 2692 13030 2694
rect 13086 2692 13110 2694
rect 13166 2692 13190 2694
rect 13246 2692 13252 2694
rect 12944 2683 13252 2692
rect 13372 2746 13492 2774
rect 13372 2106 13400 2746
rect 14657 2204 14965 2213
rect 14657 2202 14663 2204
rect 14719 2202 14743 2204
rect 14799 2202 14823 2204
rect 14879 2202 14903 2204
rect 14959 2202 14965 2204
rect 14719 2150 14721 2202
rect 14901 2150 14903 2202
rect 14657 2148 14663 2150
rect 14719 2148 14743 2150
rect 14799 2148 14823 2150
rect 14879 2148 14903 2150
rect 14959 2148 14965 2150
rect 14657 2139 14965 2148
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 15028 2038 15056 41618
rect 15120 41414 15148 41958
rect 15476 41608 15528 41614
rect 15476 41550 15528 41556
rect 15120 41386 15240 41414
rect 15108 36032 15160 36038
rect 15106 36000 15108 36009
rect 15160 36000 15162 36009
rect 15106 35935 15162 35944
rect 15108 35556 15160 35562
rect 15108 35498 15160 35504
rect 15120 34921 15148 35498
rect 15106 34912 15162 34921
rect 15106 34847 15162 34856
rect 15108 32836 15160 32842
rect 15108 32778 15160 32784
rect 15120 31657 15148 32778
rect 15106 31648 15162 31657
rect 15106 31583 15162 31592
rect 15108 30592 15160 30598
rect 15106 30560 15108 30569
rect 15160 30560 15162 30569
rect 15106 30495 15162 30504
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15120 25838 15148 27882
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 15120 24857 15148 25638
rect 15106 24848 15162 24857
rect 15106 24783 15162 24792
rect 15108 24132 15160 24138
rect 15108 24074 15160 24080
rect 15120 24041 15148 24074
rect 15106 24032 15162 24041
rect 15106 23967 15162 23976
rect 15108 22976 15160 22982
rect 15106 22944 15108 22953
rect 15160 22944 15162 22953
rect 15106 22879 15162 22888
rect 15212 22794 15240 41386
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15304 35601 15332 36518
rect 15290 35592 15346 35601
rect 15290 35527 15346 35536
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15304 29753 15332 31078
rect 15290 29744 15346 29753
rect 15290 29679 15346 29688
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15304 25673 15332 26726
rect 15290 25664 15346 25673
rect 15290 25599 15346 25608
rect 15292 25560 15344 25566
rect 15292 25502 15344 25508
rect 15120 22766 15240 22794
rect 15120 21962 15148 22766
rect 15304 22098 15332 25502
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15292 22092 15344 22098
rect 15292 22034 15344 22040
rect 15108 21956 15160 21962
rect 15108 21898 15160 21904
rect 15106 21856 15162 21865
rect 15106 21791 15162 21800
rect 15120 21146 15148 21791
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15120 18698 15148 19994
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15106 18592 15162 18601
rect 15106 18527 15162 18536
rect 15120 17882 15148 18527
rect 15212 18306 15240 22034
rect 15396 22001 15424 31282
rect 15382 21992 15438 22001
rect 15382 21927 15438 21936
rect 15384 21752 15436 21758
rect 15384 21694 15436 21700
rect 15290 20768 15346 20777
rect 15290 20703 15346 20712
rect 15304 18426 15332 20703
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15212 18278 15332 18306
rect 15198 18184 15254 18193
rect 15198 18119 15254 18128
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15212 17338 15240 18119
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15304 17270 15332 18278
rect 15292 17264 15344 17270
rect 15292 17206 15344 17212
rect 15198 16552 15254 16561
rect 15198 16487 15254 16496
rect 15106 16416 15162 16425
rect 15106 16351 15162 16360
rect 15120 15434 15148 16351
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15106 14240 15162 14249
rect 15106 14175 15162 14184
rect 15120 12850 15148 14175
rect 15212 13274 15240 16487
rect 15290 14376 15346 14385
rect 15290 14311 15346 14320
rect 15304 13394 15332 14311
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15212 13246 15332 13274
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15106 11928 15162 11937
rect 15106 11863 15162 11872
rect 15120 10674 15148 11863
rect 15212 11150 15240 13087
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15198 10976 15254 10985
rect 15198 10911 15254 10920
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15212 10062 15240 10911
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15120 9897 15148 9930
rect 15106 9888 15162 9897
rect 15106 9823 15162 9832
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15120 8809 15148 9114
rect 15106 8800 15162 8809
rect 15106 8735 15162 8744
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15120 6322 15148 6831
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15198 6216 15254 6225
rect 15198 6151 15254 6160
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15120 5302 15148 5471
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 15212 4622 15240 6151
rect 15304 5914 15332 13246
rect 15396 9722 15424 21694
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 15016 2032 15068 2038
rect 15016 1974 15068 1980
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 12944 1660 13252 1669
rect 12944 1658 12950 1660
rect 13006 1658 13030 1660
rect 13086 1658 13110 1660
rect 13166 1658 13190 1660
rect 13246 1658 13252 1660
rect 13006 1606 13008 1658
rect 13188 1606 13190 1658
rect 12944 1604 12950 1606
rect 13006 1604 13030 1606
rect 13086 1604 13110 1606
rect 13166 1604 13190 1606
rect 13246 1604 13252 1606
rect 12944 1595 13252 1604
rect 13280 1562 13308 1906
rect 13464 1562 13492 1974
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 13740 1562 13768 1906
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13452 1556 13504 1562
rect 13452 1498 13504 1504
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 15488 1358 15516 41550
rect 15568 33040 15620 33046
rect 15568 32982 15620 32988
rect 15580 25226 15608 32982
rect 15660 31816 15712 31822
rect 15660 31758 15712 31764
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15672 24818 15700 31758
rect 15764 31754 15792 42162
rect 15764 31726 15976 31754
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15764 24698 15792 29990
rect 15580 24670 15792 24698
rect 15580 20058 15608 24670
rect 15948 24290 15976 31726
rect 15764 24262 15976 24290
rect 15658 22264 15714 22273
rect 15658 22199 15714 22208
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15566 19952 15622 19961
rect 15566 19887 15622 19896
rect 15580 17882 15608 19887
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15580 11898 15608 17206
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 7546 15700 22199
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15764 2106 15792 24262
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15856 17678 15884 21830
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15856 10810 15884 13330
rect 15948 12442 15976 22986
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15752 2100 15804 2106
rect 15752 2042 15804 2048
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 13912 1352 13964 1358
rect 13912 1294 13964 1300
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 15476 1352 15528 1358
rect 15476 1294 15528 1300
rect 12532 1284 12584 1290
rect 12532 1226 12584 1232
rect 13096 1018 13124 1294
rect 13084 1012 13136 1018
rect 13084 954 13136 960
rect 13096 190 13216 218
rect 13096 160 13124 190
rect 10138 54 10456 82
rect 10138 0 10194 54
rect 10874 0 10930 160
rect 11610 0 11666 160
rect 12346 0 12402 160
rect 13082 0 13138 160
rect 13188 82 13216 190
rect 13372 82 13400 1294
rect 13188 54 13400 82
rect 13818 82 13874 160
rect 13924 82 13952 1294
rect 14568 160 14596 1294
rect 14657 1116 14965 1125
rect 14657 1114 14663 1116
rect 14719 1114 14743 1116
rect 14799 1114 14823 1116
rect 14879 1114 14903 1116
rect 14959 1114 14965 1116
rect 14719 1062 14721 1114
rect 14901 1062 14903 1114
rect 14657 1060 14663 1062
rect 14719 1060 14743 1062
rect 14799 1060 14823 1062
rect 14879 1060 14903 1062
rect 14959 1060 14965 1062
rect 14657 1051 14965 1060
rect 15292 1012 15344 1018
rect 15292 954 15344 960
rect 15304 160 15332 954
rect 13818 54 13952 82
rect 13818 0 13874 54
rect 14554 0 14610 160
rect 15290 0 15346 160
<< via2 >>
rect 754 40568 810 40624
rect 754 38936 810 38992
rect 754 38120 810 38176
rect 754 37304 810 37360
rect 754 36488 810 36544
rect 754 34856 810 34912
rect 754 33224 810 33280
rect 754 32408 810 32464
rect 754 30776 810 30832
rect 754 29960 810 30016
rect 754 29144 810 29200
rect 754 28328 810 28384
rect 754 26696 810 26752
rect 754 25064 810 25120
rect 754 24248 810 24304
rect 754 23432 810 23488
rect 754 22616 810 22672
rect 754 21800 810 21856
rect 754 20984 810 21040
rect 754 20168 810 20224
rect 754 19352 810 19408
rect 754 18536 810 18592
rect 754 16904 810 16960
rect 754 16088 810 16144
rect 846 15272 902 15328
rect 846 14456 902 14512
rect 846 12044 848 12064
rect 848 12044 900 12064
rect 900 12044 902 12064
rect 846 12008 902 12044
rect 846 11192 902 11248
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 938 9596 940 9616
rect 940 9596 992 9616
rect 992 9596 994 9616
rect 938 9560 994 9596
rect 846 7148 848 7168
rect 848 7148 900 7168
rect 900 7148 902 7168
rect 846 7112 902 7148
rect 846 6296 902 6352
rect 846 5480 902 5536
rect 938 4664 994 4720
rect 754 3848 810 3904
rect 1398 39888 1454 39944
rect 1398 35808 1454 35864
rect 4382 43546 4438 43548
rect 4462 43546 4518 43548
rect 4542 43546 4598 43548
rect 4622 43546 4678 43548
rect 4382 43494 4428 43546
rect 4428 43494 4438 43546
rect 4462 43494 4492 43546
rect 4492 43494 4504 43546
rect 4504 43494 4518 43546
rect 4542 43494 4556 43546
rect 4556 43494 4568 43546
rect 4568 43494 4598 43546
rect 4622 43494 4632 43546
rect 4632 43494 4678 43546
rect 4382 43492 4438 43494
rect 4462 43492 4518 43494
rect 4542 43492 4598 43494
rect 4622 43492 4678 43494
rect 7809 43546 7865 43548
rect 7889 43546 7945 43548
rect 7969 43546 8025 43548
rect 8049 43546 8105 43548
rect 7809 43494 7855 43546
rect 7855 43494 7865 43546
rect 7889 43494 7919 43546
rect 7919 43494 7931 43546
rect 7931 43494 7945 43546
rect 7969 43494 7983 43546
rect 7983 43494 7995 43546
rect 7995 43494 8025 43546
rect 8049 43494 8059 43546
rect 8059 43494 8105 43546
rect 7809 43492 7865 43494
rect 7889 43492 7945 43494
rect 7969 43492 8025 43494
rect 8049 43492 8105 43494
rect 11236 43546 11292 43548
rect 11316 43546 11372 43548
rect 11396 43546 11452 43548
rect 11476 43546 11532 43548
rect 11236 43494 11282 43546
rect 11282 43494 11292 43546
rect 11316 43494 11346 43546
rect 11346 43494 11358 43546
rect 11358 43494 11372 43546
rect 11396 43494 11410 43546
rect 11410 43494 11422 43546
rect 11422 43494 11452 43546
rect 11476 43494 11486 43546
rect 11486 43494 11532 43546
rect 11236 43492 11292 43494
rect 11316 43492 11372 43494
rect 11396 43492 11452 43494
rect 11476 43492 11532 43494
rect 1398 34448 1454 34504
rect 1398 31592 1454 31648
rect 1490 27512 1546 27568
rect 1674 27648 1730 27704
rect 1490 26152 1546 26208
rect 1582 21392 1638 21448
rect 1490 17856 1546 17912
rect 1674 14048 1730 14104
rect 1950 12960 2006 13016
rect 1398 9016 1454 9072
rect 1582 8336 1638 8392
rect 1858 8200 1914 8256
rect 2669 43002 2725 43004
rect 2749 43002 2805 43004
rect 2829 43002 2885 43004
rect 2909 43002 2965 43004
rect 2669 42950 2715 43002
rect 2715 42950 2725 43002
rect 2749 42950 2779 43002
rect 2779 42950 2791 43002
rect 2791 42950 2805 43002
rect 2829 42950 2843 43002
rect 2843 42950 2855 43002
rect 2855 42950 2885 43002
rect 2909 42950 2919 43002
rect 2919 42950 2965 43002
rect 2669 42948 2725 42950
rect 2749 42948 2805 42950
rect 2829 42948 2885 42950
rect 2909 42948 2965 42950
rect 2669 41914 2725 41916
rect 2749 41914 2805 41916
rect 2829 41914 2885 41916
rect 2909 41914 2965 41916
rect 2669 41862 2715 41914
rect 2715 41862 2725 41914
rect 2749 41862 2779 41914
rect 2779 41862 2791 41914
rect 2791 41862 2805 41914
rect 2829 41862 2843 41914
rect 2843 41862 2855 41914
rect 2855 41862 2885 41914
rect 2909 41862 2919 41914
rect 2919 41862 2965 41914
rect 2669 41860 2725 41862
rect 2749 41860 2805 41862
rect 2829 41860 2885 41862
rect 2909 41860 2965 41862
rect 2669 40826 2725 40828
rect 2749 40826 2805 40828
rect 2829 40826 2885 40828
rect 2909 40826 2965 40828
rect 2669 40774 2715 40826
rect 2715 40774 2725 40826
rect 2749 40774 2779 40826
rect 2779 40774 2791 40826
rect 2791 40774 2805 40826
rect 2829 40774 2843 40826
rect 2843 40774 2855 40826
rect 2855 40774 2885 40826
rect 2909 40774 2919 40826
rect 2919 40774 2965 40826
rect 2669 40772 2725 40774
rect 2749 40772 2805 40774
rect 2829 40772 2885 40774
rect 2909 40772 2965 40774
rect 2669 39738 2725 39740
rect 2749 39738 2805 39740
rect 2829 39738 2885 39740
rect 2909 39738 2965 39740
rect 2669 39686 2715 39738
rect 2715 39686 2725 39738
rect 2749 39686 2779 39738
rect 2779 39686 2791 39738
rect 2791 39686 2805 39738
rect 2829 39686 2843 39738
rect 2843 39686 2855 39738
rect 2855 39686 2885 39738
rect 2909 39686 2919 39738
rect 2919 39686 2965 39738
rect 2669 39684 2725 39686
rect 2749 39684 2805 39686
rect 2829 39684 2885 39686
rect 2909 39684 2965 39686
rect 2669 38650 2725 38652
rect 2749 38650 2805 38652
rect 2829 38650 2885 38652
rect 2909 38650 2965 38652
rect 2669 38598 2715 38650
rect 2715 38598 2725 38650
rect 2749 38598 2779 38650
rect 2779 38598 2791 38650
rect 2791 38598 2805 38650
rect 2829 38598 2843 38650
rect 2843 38598 2855 38650
rect 2855 38598 2885 38650
rect 2909 38598 2919 38650
rect 2919 38598 2965 38650
rect 2669 38596 2725 38598
rect 2749 38596 2805 38598
rect 2829 38596 2885 38598
rect 2909 38596 2965 38598
rect 2669 37562 2725 37564
rect 2749 37562 2805 37564
rect 2829 37562 2885 37564
rect 2909 37562 2965 37564
rect 2669 37510 2715 37562
rect 2715 37510 2725 37562
rect 2749 37510 2779 37562
rect 2779 37510 2791 37562
rect 2791 37510 2805 37562
rect 2829 37510 2843 37562
rect 2843 37510 2855 37562
rect 2855 37510 2885 37562
rect 2909 37510 2919 37562
rect 2919 37510 2965 37562
rect 2669 37508 2725 37510
rect 2749 37508 2805 37510
rect 2829 37508 2885 37510
rect 2909 37508 2965 37510
rect 2669 36474 2725 36476
rect 2749 36474 2805 36476
rect 2829 36474 2885 36476
rect 2909 36474 2965 36476
rect 2669 36422 2715 36474
rect 2715 36422 2725 36474
rect 2749 36422 2779 36474
rect 2779 36422 2791 36474
rect 2791 36422 2805 36474
rect 2829 36422 2843 36474
rect 2843 36422 2855 36474
rect 2855 36422 2885 36474
rect 2909 36422 2919 36474
rect 2919 36422 2965 36474
rect 2669 36420 2725 36422
rect 2749 36420 2805 36422
rect 2829 36420 2885 36422
rect 2909 36420 2965 36422
rect 2669 35386 2725 35388
rect 2749 35386 2805 35388
rect 2829 35386 2885 35388
rect 2909 35386 2965 35388
rect 2669 35334 2715 35386
rect 2715 35334 2725 35386
rect 2749 35334 2779 35386
rect 2779 35334 2791 35386
rect 2791 35334 2805 35386
rect 2829 35334 2843 35386
rect 2843 35334 2855 35386
rect 2855 35334 2885 35386
rect 2909 35334 2919 35386
rect 2919 35334 2965 35386
rect 2669 35332 2725 35334
rect 2749 35332 2805 35334
rect 2829 35332 2885 35334
rect 2909 35332 2965 35334
rect 2669 34298 2725 34300
rect 2749 34298 2805 34300
rect 2829 34298 2885 34300
rect 2909 34298 2965 34300
rect 2669 34246 2715 34298
rect 2715 34246 2725 34298
rect 2749 34246 2779 34298
rect 2779 34246 2791 34298
rect 2791 34246 2805 34298
rect 2829 34246 2843 34298
rect 2843 34246 2855 34298
rect 2855 34246 2885 34298
rect 2909 34246 2919 34298
rect 2919 34246 2965 34298
rect 2669 34244 2725 34246
rect 2749 34244 2805 34246
rect 2829 34244 2885 34246
rect 2909 34244 2965 34246
rect 2669 33210 2725 33212
rect 2749 33210 2805 33212
rect 2829 33210 2885 33212
rect 2909 33210 2965 33212
rect 2669 33158 2715 33210
rect 2715 33158 2725 33210
rect 2749 33158 2779 33210
rect 2779 33158 2791 33210
rect 2791 33158 2805 33210
rect 2829 33158 2843 33210
rect 2843 33158 2855 33210
rect 2855 33158 2885 33210
rect 2909 33158 2919 33210
rect 2919 33158 2965 33210
rect 2669 33156 2725 33158
rect 2749 33156 2805 33158
rect 2829 33156 2885 33158
rect 2909 33156 2965 33158
rect 2669 32122 2725 32124
rect 2749 32122 2805 32124
rect 2829 32122 2885 32124
rect 2909 32122 2965 32124
rect 2669 32070 2715 32122
rect 2715 32070 2725 32122
rect 2749 32070 2779 32122
rect 2779 32070 2791 32122
rect 2791 32070 2805 32122
rect 2829 32070 2843 32122
rect 2843 32070 2855 32122
rect 2855 32070 2885 32122
rect 2909 32070 2919 32122
rect 2919 32070 2965 32122
rect 2669 32068 2725 32070
rect 2749 32068 2805 32070
rect 2829 32068 2885 32070
rect 2909 32068 2965 32070
rect 2669 31034 2725 31036
rect 2749 31034 2805 31036
rect 2829 31034 2885 31036
rect 2909 31034 2965 31036
rect 2669 30982 2715 31034
rect 2715 30982 2725 31034
rect 2749 30982 2779 31034
rect 2779 30982 2791 31034
rect 2791 30982 2805 31034
rect 2829 30982 2843 31034
rect 2843 30982 2855 31034
rect 2855 30982 2885 31034
rect 2909 30982 2919 31034
rect 2919 30982 2965 31034
rect 2669 30980 2725 30982
rect 2749 30980 2805 30982
rect 2829 30980 2885 30982
rect 2909 30980 2965 30982
rect 2669 29946 2725 29948
rect 2749 29946 2805 29948
rect 2829 29946 2885 29948
rect 2909 29946 2965 29948
rect 2669 29894 2715 29946
rect 2715 29894 2725 29946
rect 2749 29894 2779 29946
rect 2779 29894 2791 29946
rect 2791 29894 2805 29946
rect 2829 29894 2843 29946
rect 2843 29894 2855 29946
rect 2855 29894 2885 29946
rect 2909 29894 2919 29946
rect 2919 29894 2965 29946
rect 2669 29892 2725 29894
rect 2749 29892 2805 29894
rect 2829 29892 2885 29894
rect 2909 29892 2965 29894
rect 2669 28858 2725 28860
rect 2749 28858 2805 28860
rect 2829 28858 2885 28860
rect 2909 28858 2965 28860
rect 2669 28806 2715 28858
rect 2715 28806 2725 28858
rect 2749 28806 2779 28858
rect 2779 28806 2791 28858
rect 2791 28806 2805 28858
rect 2829 28806 2843 28858
rect 2843 28806 2855 28858
rect 2855 28806 2885 28858
rect 2909 28806 2919 28858
rect 2919 28806 2965 28858
rect 2669 28804 2725 28806
rect 2749 28804 2805 28806
rect 2829 28804 2885 28806
rect 2909 28804 2965 28806
rect 2669 27770 2725 27772
rect 2749 27770 2805 27772
rect 2829 27770 2885 27772
rect 2909 27770 2965 27772
rect 2669 27718 2715 27770
rect 2715 27718 2725 27770
rect 2749 27718 2779 27770
rect 2779 27718 2791 27770
rect 2791 27718 2805 27770
rect 2829 27718 2843 27770
rect 2843 27718 2855 27770
rect 2855 27718 2885 27770
rect 2909 27718 2919 27770
rect 2919 27718 2965 27770
rect 2669 27716 2725 27718
rect 2749 27716 2805 27718
rect 2829 27716 2885 27718
rect 2909 27716 2965 27718
rect 2669 26682 2725 26684
rect 2749 26682 2805 26684
rect 2829 26682 2885 26684
rect 2909 26682 2965 26684
rect 2669 26630 2715 26682
rect 2715 26630 2725 26682
rect 2749 26630 2779 26682
rect 2779 26630 2791 26682
rect 2791 26630 2805 26682
rect 2829 26630 2843 26682
rect 2843 26630 2855 26682
rect 2855 26630 2885 26682
rect 2909 26630 2919 26682
rect 2919 26630 2965 26682
rect 2669 26628 2725 26630
rect 2749 26628 2805 26630
rect 2829 26628 2885 26630
rect 2909 26628 2965 26630
rect 2669 25594 2725 25596
rect 2749 25594 2805 25596
rect 2829 25594 2885 25596
rect 2909 25594 2965 25596
rect 2669 25542 2715 25594
rect 2715 25542 2725 25594
rect 2749 25542 2779 25594
rect 2779 25542 2791 25594
rect 2791 25542 2805 25594
rect 2829 25542 2843 25594
rect 2843 25542 2855 25594
rect 2855 25542 2885 25594
rect 2909 25542 2919 25594
rect 2919 25542 2965 25594
rect 2669 25540 2725 25542
rect 2749 25540 2805 25542
rect 2829 25540 2885 25542
rect 2909 25540 2965 25542
rect 2669 24506 2725 24508
rect 2749 24506 2805 24508
rect 2829 24506 2885 24508
rect 2909 24506 2965 24508
rect 2669 24454 2715 24506
rect 2715 24454 2725 24506
rect 2749 24454 2779 24506
rect 2779 24454 2791 24506
rect 2791 24454 2805 24506
rect 2829 24454 2843 24506
rect 2843 24454 2855 24506
rect 2855 24454 2885 24506
rect 2909 24454 2919 24506
rect 2919 24454 2965 24506
rect 2669 24452 2725 24454
rect 2749 24452 2805 24454
rect 2829 24452 2885 24454
rect 2909 24452 2965 24454
rect 2669 23418 2725 23420
rect 2749 23418 2805 23420
rect 2829 23418 2885 23420
rect 2909 23418 2965 23420
rect 2669 23366 2715 23418
rect 2715 23366 2725 23418
rect 2749 23366 2779 23418
rect 2779 23366 2791 23418
rect 2791 23366 2805 23418
rect 2829 23366 2843 23418
rect 2843 23366 2855 23418
rect 2855 23366 2885 23418
rect 2909 23366 2919 23418
rect 2919 23366 2965 23418
rect 2669 23364 2725 23366
rect 2749 23364 2805 23366
rect 2829 23364 2885 23366
rect 2909 23364 2965 23366
rect 2669 22330 2725 22332
rect 2749 22330 2805 22332
rect 2829 22330 2885 22332
rect 2909 22330 2965 22332
rect 2669 22278 2715 22330
rect 2715 22278 2725 22330
rect 2749 22278 2779 22330
rect 2779 22278 2791 22330
rect 2791 22278 2805 22330
rect 2829 22278 2843 22330
rect 2843 22278 2855 22330
rect 2855 22278 2885 22330
rect 2909 22278 2919 22330
rect 2919 22278 2965 22330
rect 2669 22276 2725 22278
rect 2749 22276 2805 22278
rect 2829 22276 2885 22278
rect 2909 22276 2965 22278
rect 2669 21242 2725 21244
rect 2749 21242 2805 21244
rect 2829 21242 2885 21244
rect 2909 21242 2965 21244
rect 2669 21190 2715 21242
rect 2715 21190 2725 21242
rect 2749 21190 2779 21242
rect 2779 21190 2791 21242
rect 2791 21190 2805 21242
rect 2829 21190 2843 21242
rect 2843 21190 2855 21242
rect 2855 21190 2885 21242
rect 2909 21190 2919 21242
rect 2919 21190 2965 21242
rect 2669 21188 2725 21190
rect 2749 21188 2805 21190
rect 2829 21188 2885 21190
rect 2909 21188 2965 21190
rect 2669 20154 2725 20156
rect 2749 20154 2805 20156
rect 2829 20154 2885 20156
rect 2909 20154 2965 20156
rect 2669 20102 2715 20154
rect 2715 20102 2725 20154
rect 2749 20102 2779 20154
rect 2779 20102 2791 20154
rect 2791 20102 2805 20154
rect 2829 20102 2843 20154
rect 2843 20102 2855 20154
rect 2855 20102 2885 20154
rect 2909 20102 2919 20154
rect 2919 20102 2965 20154
rect 2669 20100 2725 20102
rect 2749 20100 2805 20102
rect 2829 20100 2885 20102
rect 2909 20100 2965 20102
rect 2669 19066 2725 19068
rect 2749 19066 2805 19068
rect 2829 19066 2885 19068
rect 2909 19066 2965 19068
rect 2669 19014 2715 19066
rect 2715 19014 2725 19066
rect 2749 19014 2779 19066
rect 2779 19014 2791 19066
rect 2791 19014 2805 19066
rect 2829 19014 2843 19066
rect 2843 19014 2855 19066
rect 2855 19014 2885 19066
rect 2909 19014 2919 19066
rect 2919 19014 2965 19066
rect 2669 19012 2725 19014
rect 2749 19012 2805 19014
rect 2829 19012 2885 19014
rect 2909 19012 2965 19014
rect 2669 17978 2725 17980
rect 2749 17978 2805 17980
rect 2829 17978 2885 17980
rect 2909 17978 2965 17980
rect 2669 17926 2715 17978
rect 2715 17926 2725 17978
rect 2749 17926 2779 17978
rect 2779 17926 2791 17978
rect 2791 17926 2805 17978
rect 2829 17926 2843 17978
rect 2843 17926 2855 17978
rect 2855 17926 2885 17978
rect 2909 17926 2919 17978
rect 2919 17926 2965 17978
rect 2669 17924 2725 17926
rect 2749 17924 2805 17926
rect 2829 17924 2885 17926
rect 2909 17924 2965 17926
rect 2669 16890 2725 16892
rect 2749 16890 2805 16892
rect 2829 16890 2885 16892
rect 2909 16890 2965 16892
rect 2669 16838 2715 16890
rect 2715 16838 2725 16890
rect 2749 16838 2779 16890
rect 2779 16838 2791 16890
rect 2791 16838 2805 16890
rect 2829 16838 2843 16890
rect 2843 16838 2855 16890
rect 2855 16838 2885 16890
rect 2909 16838 2919 16890
rect 2919 16838 2965 16890
rect 2669 16836 2725 16838
rect 2749 16836 2805 16838
rect 2829 16836 2885 16838
rect 2909 16836 2965 16838
rect 2669 15802 2725 15804
rect 2749 15802 2805 15804
rect 2829 15802 2885 15804
rect 2909 15802 2965 15804
rect 2669 15750 2715 15802
rect 2715 15750 2725 15802
rect 2749 15750 2779 15802
rect 2779 15750 2791 15802
rect 2791 15750 2805 15802
rect 2829 15750 2843 15802
rect 2843 15750 2855 15802
rect 2855 15750 2885 15802
rect 2909 15750 2919 15802
rect 2919 15750 2965 15802
rect 2669 15748 2725 15750
rect 2749 15748 2805 15750
rect 2829 15748 2885 15750
rect 2909 15748 2965 15750
rect 2669 14714 2725 14716
rect 2749 14714 2805 14716
rect 2829 14714 2885 14716
rect 2909 14714 2965 14716
rect 2669 14662 2715 14714
rect 2715 14662 2725 14714
rect 2749 14662 2779 14714
rect 2779 14662 2791 14714
rect 2791 14662 2805 14714
rect 2829 14662 2843 14714
rect 2843 14662 2855 14714
rect 2855 14662 2885 14714
rect 2909 14662 2919 14714
rect 2919 14662 2965 14714
rect 2669 14660 2725 14662
rect 2749 14660 2805 14662
rect 2829 14660 2885 14662
rect 2909 14660 2965 14662
rect 2502 13676 2504 13696
rect 2504 13676 2556 13696
rect 2556 13676 2558 13696
rect 2502 13640 2558 13676
rect 2669 13626 2725 13628
rect 2749 13626 2805 13628
rect 2829 13626 2885 13628
rect 2909 13626 2965 13628
rect 2669 13574 2715 13626
rect 2715 13574 2725 13626
rect 2749 13574 2779 13626
rect 2779 13574 2791 13626
rect 2791 13574 2805 13626
rect 2829 13574 2843 13626
rect 2843 13574 2855 13626
rect 2855 13574 2885 13626
rect 2909 13574 2919 13626
rect 2919 13574 2965 13626
rect 2669 13572 2725 13574
rect 2749 13572 2805 13574
rect 2829 13572 2885 13574
rect 2909 13572 2965 13574
rect 2669 12538 2725 12540
rect 2749 12538 2805 12540
rect 2829 12538 2885 12540
rect 2909 12538 2965 12540
rect 2669 12486 2715 12538
rect 2715 12486 2725 12538
rect 2749 12486 2779 12538
rect 2779 12486 2791 12538
rect 2791 12486 2805 12538
rect 2829 12486 2843 12538
rect 2843 12486 2855 12538
rect 2855 12486 2885 12538
rect 2909 12486 2919 12538
rect 2919 12486 2965 12538
rect 2669 12484 2725 12486
rect 2749 12484 2805 12486
rect 2829 12484 2885 12486
rect 2909 12484 2965 12486
rect 2669 11450 2725 11452
rect 2749 11450 2805 11452
rect 2829 11450 2885 11452
rect 2909 11450 2965 11452
rect 2669 11398 2715 11450
rect 2715 11398 2725 11450
rect 2749 11398 2779 11450
rect 2779 11398 2791 11450
rect 2791 11398 2805 11450
rect 2829 11398 2843 11450
rect 2843 11398 2855 11450
rect 2855 11398 2885 11450
rect 2909 11398 2919 11450
rect 2919 11398 2965 11450
rect 2669 11396 2725 11398
rect 2749 11396 2805 11398
rect 2829 11396 2885 11398
rect 2909 11396 2965 11398
rect 2669 10362 2725 10364
rect 2749 10362 2805 10364
rect 2829 10362 2885 10364
rect 2909 10362 2965 10364
rect 2669 10310 2715 10362
rect 2715 10310 2725 10362
rect 2749 10310 2779 10362
rect 2779 10310 2791 10362
rect 2791 10310 2805 10362
rect 2829 10310 2843 10362
rect 2843 10310 2855 10362
rect 2855 10310 2885 10362
rect 2909 10310 2919 10362
rect 2919 10310 2965 10362
rect 2669 10308 2725 10310
rect 2749 10308 2805 10310
rect 2829 10308 2885 10310
rect 2909 10308 2965 10310
rect 2669 9274 2725 9276
rect 2749 9274 2805 9276
rect 2829 9274 2885 9276
rect 2909 9274 2965 9276
rect 2669 9222 2715 9274
rect 2715 9222 2725 9274
rect 2749 9222 2779 9274
rect 2779 9222 2791 9274
rect 2791 9222 2805 9274
rect 2829 9222 2843 9274
rect 2843 9222 2855 9274
rect 2855 9222 2885 9274
rect 2909 9222 2919 9274
rect 2919 9222 2965 9274
rect 2669 9220 2725 9222
rect 2749 9220 2805 9222
rect 2829 9220 2885 9222
rect 2909 9220 2965 9222
rect 2669 8186 2725 8188
rect 2749 8186 2805 8188
rect 2829 8186 2885 8188
rect 2909 8186 2965 8188
rect 2669 8134 2715 8186
rect 2715 8134 2725 8186
rect 2749 8134 2779 8186
rect 2779 8134 2791 8186
rect 2791 8134 2805 8186
rect 2829 8134 2843 8186
rect 2843 8134 2855 8186
rect 2855 8134 2885 8186
rect 2909 8134 2919 8186
rect 2919 8134 2965 8186
rect 2669 8132 2725 8134
rect 2749 8132 2805 8134
rect 2829 8132 2885 8134
rect 2909 8132 2965 8134
rect 2669 7098 2725 7100
rect 2749 7098 2805 7100
rect 2829 7098 2885 7100
rect 2909 7098 2965 7100
rect 2669 7046 2715 7098
rect 2715 7046 2725 7098
rect 2749 7046 2779 7098
rect 2779 7046 2791 7098
rect 2791 7046 2805 7098
rect 2829 7046 2843 7098
rect 2843 7046 2855 7098
rect 2855 7046 2885 7098
rect 2909 7046 2919 7098
rect 2919 7046 2965 7098
rect 2669 7044 2725 7046
rect 2749 7044 2805 7046
rect 2829 7044 2885 7046
rect 2909 7044 2965 7046
rect 2669 6010 2725 6012
rect 2749 6010 2805 6012
rect 2829 6010 2885 6012
rect 2909 6010 2965 6012
rect 2669 5958 2715 6010
rect 2715 5958 2725 6010
rect 2749 5958 2779 6010
rect 2779 5958 2791 6010
rect 2791 5958 2805 6010
rect 2829 5958 2843 6010
rect 2843 5958 2855 6010
rect 2855 5958 2885 6010
rect 2909 5958 2919 6010
rect 2919 5958 2965 6010
rect 2669 5956 2725 5958
rect 2749 5956 2805 5958
rect 2829 5956 2885 5958
rect 2909 5956 2965 5958
rect 2669 4922 2725 4924
rect 2749 4922 2805 4924
rect 2829 4922 2885 4924
rect 2909 4922 2965 4924
rect 2669 4870 2715 4922
rect 2715 4870 2725 4922
rect 2749 4870 2779 4922
rect 2779 4870 2791 4922
rect 2791 4870 2805 4922
rect 2829 4870 2843 4922
rect 2843 4870 2855 4922
rect 2855 4870 2885 4922
rect 2909 4870 2919 4922
rect 2919 4870 2965 4922
rect 2669 4868 2725 4870
rect 2749 4868 2805 4870
rect 2829 4868 2885 4870
rect 2909 4868 2965 4870
rect 2669 3834 2725 3836
rect 2749 3834 2805 3836
rect 2829 3834 2885 3836
rect 2909 3834 2965 3836
rect 2669 3782 2715 3834
rect 2715 3782 2725 3834
rect 2749 3782 2779 3834
rect 2779 3782 2791 3834
rect 2791 3782 2805 3834
rect 2829 3782 2843 3834
rect 2843 3782 2855 3834
rect 2855 3782 2885 3834
rect 2909 3782 2919 3834
rect 2919 3782 2965 3834
rect 2669 3780 2725 3782
rect 2749 3780 2805 3782
rect 2829 3780 2885 3782
rect 2909 3780 2965 3782
rect 2669 2746 2725 2748
rect 2749 2746 2805 2748
rect 2829 2746 2885 2748
rect 2909 2746 2965 2748
rect 2669 2694 2715 2746
rect 2715 2694 2725 2746
rect 2749 2694 2779 2746
rect 2779 2694 2791 2746
rect 2791 2694 2805 2746
rect 2829 2694 2843 2746
rect 2843 2694 2855 2746
rect 2855 2694 2885 2746
rect 2909 2694 2919 2746
rect 2919 2694 2965 2746
rect 2669 2692 2725 2694
rect 2749 2692 2805 2694
rect 2829 2692 2885 2694
rect 2909 2692 2965 2694
rect 4382 42458 4438 42460
rect 4462 42458 4518 42460
rect 4542 42458 4598 42460
rect 4622 42458 4678 42460
rect 4382 42406 4428 42458
rect 4428 42406 4438 42458
rect 4462 42406 4492 42458
rect 4492 42406 4504 42458
rect 4504 42406 4518 42458
rect 4542 42406 4556 42458
rect 4556 42406 4568 42458
rect 4568 42406 4598 42458
rect 4622 42406 4632 42458
rect 4632 42406 4678 42458
rect 4382 42404 4438 42406
rect 4462 42404 4518 42406
rect 4542 42404 4598 42406
rect 4622 42404 4678 42406
rect 3330 6160 3386 6216
rect 4382 41370 4438 41372
rect 4462 41370 4518 41372
rect 4542 41370 4598 41372
rect 4622 41370 4678 41372
rect 4382 41318 4428 41370
rect 4428 41318 4438 41370
rect 4462 41318 4492 41370
rect 4492 41318 4504 41370
rect 4504 41318 4518 41370
rect 4542 41318 4556 41370
rect 4556 41318 4568 41370
rect 4568 41318 4598 41370
rect 4622 41318 4632 41370
rect 4632 41318 4678 41370
rect 4382 41316 4438 41318
rect 4462 41316 4518 41318
rect 4542 41316 4598 41318
rect 4622 41316 4678 41318
rect 4382 40282 4438 40284
rect 4462 40282 4518 40284
rect 4542 40282 4598 40284
rect 4622 40282 4678 40284
rect 4382 40230 4428 40282
rect 4428 40230 4438 40282
rect 4462 40230 4492 40282
rect 4492 40230 4504 40282
rect 4504 40230 4518 40282
rect 4542 40230 4556 40282
rect 4556 40230 4568 40282
rect 4568 40230 4598 40282
rect 4622 40230 4632 40282
rect 4632 40230 4678 40282
rect 4382 40228 4438 40230
rect 4462 40228 4518 40230
rect 4542 40228 4598 40230
rect 4622 40228 4678 40230
rect 4382 39194 4438 39196
rect 4462 39194 4518 39196
rect 4542 39194 4598 39196
rect 4622 39194 4678 39196
rect 4382 39142 4428 39194
rect 4428 39142 4438 39194
rect 4462 39142 4492 39194
rect 4492 39142 4504 39194
rect 4504 39142 4518 39194
rect 4542 39142 4556 39194
rect 4556 39142 4568 39194
rect 4568 39142 4598 39194
rect 4622 39142 4632 39194
rect 4632 39142 4678 39194
rect 4382 39140 4438 39142
rect 4462 39140 4518 39142
rect 4542 39140 4598 39142
rect 4622 39140 4678 39142
rect 6096 43002 6152 43004
rect 6176 43002 6232 43004
rect 6256 43002 6312 43004
rect 6336 43002 6392 43004
rect 6096 42950 6142 43002
rect 6142 42950 6152 43002
rect 6176 42950 6206 43002
rect 6206 42950 6218 43002
rect 6218 42950 6232 43002
rect 6256 42950 6270 43002
rect 6270 42950 6282 43002
rect 6282 42950 6312 43002
rect 6336 42950 6346 43002
rect 6346 42950 6392 43002
rect 6096 42948 6152 42950
rect 6176 42948 6232 42950
rect 6256 42948 6312 42950
rect 6336 42948 6392 42950
rect 9523 43002 9579 43004
rect 9603 43002 9659 43004
rect 9683 43002 9739 43004
rect 9763 43002 9819 43004
rect 9523 42950 9569 43002
rect 9569 42950 9579 43002
rect 9603 42950 9633 43002
rect 9633 42950 9645 43002
rect 9645 42950 9659 43002
rect 9683 42950 9697 43002
rect 9697 42950 9709 43002
rect 9709 42950 9739 43002
rect 9763 42950 9773 43002
rect 9773 42950 9819 43002
rect 9523 42948 9579 42950
rect 9603 42948 9659 42950
rect 9683 42948 9739 42950
rect 9763 42948 9819 42950
rect 12950 43002 13006 43004
rect 13030 43002 13086 43004
rect 13110 43002 13166 43004
rect 13190 43002 13246 43004
rect 12950 42950 12996 43002
rect 12996 42950 13006 43002
rect 13030 42950 13060 43002
rect 13060 42950 13072 43002
rect 13072 42950 13086 43002
rect 13110 42950 13124 43002
rect 13124 42950 13136 43002
rect 13136 42950 13166 43002
rect 13190 42950 13200 43002
rect 13200 42950 13246 43002
rect 12950 42948 13006 42950
rect 13030 42948 13086 42950
rect 13110 42948 13166 42950
rect 13190 42948 13246 42950
rect 14663 43546 14719 43548
rect 14743 43546 14799 43548
rect 14823 43546 14879 43548
rect 14903 43546 14959 43548
rect 14663 43494 14709 43546
rect 14709 43494 14719 43546
rect 14743 43494 14773 43546
rect 14773 43494 14785 43546
rect 14785 43494 14799 43546
rect 14823 43494 14837 43546
rect 14837 43494 14849 43546
rect 14849 43494 14879 43546
rect 14903 43494 14913 43546
rect 14913 43494 14959 43546
rect 14663 43492 14719 43494
rect 14743 43492 14799 43494
rect 14823 43492 14879 43494
rect 14903 43492 14959 43494
rect 7809 42458 7865 42460
rect 7889 42458 7945 42460
rect 7969 42458 8025 42460
rect 8049 42458 8105 42460
rect 7809 42406 7855 42458
rect 7855 42406 7865 42458
rect 7889 42406 7919 42458
rect 7919 42406 7931 42458
rect 7931 42406 7945 42458
rect 7969 42406 7983 42458
rect 7983 42406 7995 42458
rect 7995 42406 8025 42458
rect 8049 42406 8059 42458
rect 8059 42406 8105 42458
rect 7809 42404 7865 42406
rect 7889 42404 7945 42406
rect 7969 42404 8025 42406
rect 8049 42404 8105 42406
rect 11236 42458 11292 42460
rect 11316 42458 11372 42460
rect 11396 42458 11452 42460
rect 11476 42458 11532 42460
rect 11236 42406 11282 42458
rect 11282 42406 11292 42458
rect 11316 42406 11346 42458
rect 11346 42406 11358 42458
rect 11358 42406 11372 42458
rect 11396 42406 11410 42458
rect 11410 42406 11422 42458
rect 11422 42406 11452 42458
rect 11476 42406 11486 42458
rect 11486 42406 11532 42458
rect 11236 42404 11292 42406
rect 11316 42404 11372 42406
rect 11396 42404 11452 42406
rect 11476 42404 11532 42406
rect 14663 42458 14719 42460
rect 14743 42458 14799 42460
rect 14823 42458 14879 42460
rect 14903 42458 14959 42460
rect 14663 42406 14709 42458
rect 14709 42406 14719 42458
rect 14743 42406 14773 42458
rect 14773 42406 14785 42458
rect 14785 42406 14799 42458
rect 14823 42406 14837 42458
rect 14837 42406 14849 42458
rect 14849 42406 14879 42458
rect 14903 42406 14913 42458
rect 14913 42406 14959 42458
rect 14663 42404 14719 42406
rect 14743 42404 14799 42406
rect 14823 42404 14879 42406
rect 14903 42404 14959 42406
rect 6096 41914 6152 41916
rect 6176 41914 6232 41916
rect 6256 41914 6312 41916
rect 6336 41914 6392 41916
rect 6096 41862 6142 41914
rect 6142 41862 6152 41914
rect 6176 41862 6206 41914
rect 6206 41862 6218 41914
rect 6218 41862 6232 41914
rect 6256 41862 6270 41914
rect 6270 41862 6282 41914
rect 6282 41862 6312 41914
rect 6336 41862 6346 41914
rect 6346 41862 6392 41914
rect 6096 41860 6152 41862
rect 6176 41860 6232 41862
rect 6256 41860 6312 41862
rect 6336 41860 6392 41862
rect 5722 41792 5778 41848
rect 6550 41792 6606 41848
rect 9523 41914 9579 41916
rect 9603 41914 9659 41916
rect 9683 41914 9739 41916
rect 9763 41914 9819 41916
rect 9523 41862 9569 41914
rect 9569 41862 9579 41914
rect 9603 41862 9633 41914
rect 9633 41862 9645 41914
rect 9645 41862 9659 41914
rect 9683 41862 9697 41914
rect 9697 41862 9709 41914
rect 9709 41862 9739 41914
rect 9763 41862 9773 41914
rect 9773 41862 9819 41914
rect 9523 41860 9579 41862
rect 9603 41860 9659 41862
rect 9683 41860 9739 41862
rect 9763 41860 9819 41862
rect 11702 42064 11758 42120
rect 8114 41792 8170 41848
rect 10966 41792 11022 41848
rect 12950 41914 13006 41916
rect 13030 41914 13086 41916
rect 13110 41914 13166 41916
rect 13190 41914 13246 41916
rect 12950 41862 12996 41914
rect 12996 41862 13006 41914
rect 13030 41862 13060 41914
rect 13060 41862 13072 41914
rect 13072 41862 13086 41914
rect 13110 41862 13124 41914
rect 13124 41862 13136 41914
rect 13136 41862 13166 41914
rect 13190 41862 13200 41914
rect 13200 41862 13246 41914
rect 12950 41860 13006 41862
rect 13030 41860 13086 41862
rect 13110 41860 13166 41862
rect 13190 41860 13246 41862
rect 6096 40826 6152 40828
rect 6176 40826 6232 40828
rect 6256 40826 6312 40828
rect 6336 40826 6392 40828
rect 6096 40774 6142 40826
rect 6142 40774 6152 40826
rect 6176 40774 6206 40826
rect 6206 40774 6218 40826
rect 6218 40774 6232 40826
rect 6256 40774 6270 40826
rect 6270 40774 6282 40826
rect 6282 40774 6312 40826
rect 6336 40774 6346 40826
rect 6346 40774 6392 40826
rect 6096 40772 6152 40774
rect 6176 40772 6232 40774
rect 6256 40772 6312 40774
rect 6336 40772 6392 40774
rect 6096 39738 6152 39740
rect 6176 39738 6232 39740
rect 6256 39738 6312 39740
rect 6336 39738 6392 39740
rect 6096 39686 6142 39738
rect 6142 39686 6152 39738
rect 6176 39686 6206 39738
rect 6206 39686 6218 39738
rect 6218 39686 6232 39738
rect 6256 39686 6270 39738
rect 6270 39686 6282 39738
rect 6282 39686 6312 39738
rect 6336 39686 6346 39738
rect 6346 39686 6392 39738
rect 6096 39684 6152 39686
rect 6176 39684 6232 39686
rect 6256 39684 6312 39686
rect 6336 39684 6392 39686
rect 6096 38650 6152 38652
rect 6176 38650 6232 38652
rect 6256 38650 6312 38652
rect 6336 38650 6392 38652
rect 6096 38598 6142 38650
rect 6142 38598 6152 38650
rect 6176 38598 6206 38650
rect 6206 38598 6218 38650
rect 6218 38598 6232 38650
rect 6256 38598 6270 38650
rect 6270 38598 6282 38650
rect 6282 38598 6312 38650
rect 6336 38598 6346 38650
rect 6346 38598 6392 38650
rect 6096 38596 6152 38598
rect 6176 38596 6232 38598
rect 6256 38596 6312 38598
rect 6336 38596 6392 38598
rect 4382 38106 4438 38108
rect 4462 38106 4518 38108
rect 4542 38106 4598 38108
rect 4622 38106 4678 38108
rect 4382 38054 4428 38106
rect 4428 38054 4438 38106
rect 4462 38054 4492 38106
rect 4492 38054 4504 38106
rect 4504 38054 4518 38106
rect 4542 38054 4556 38106
rect 4556 38054 4568 38106
rect 4568 38054 4598 38106
rect 4622 38054 4632 38106
rect 4632 38054 4678 38106
rect 4382 38052 4438 38054
rect 4462 38052 4518 38054
rect 4542 38052 4598 38054
rect 4622 38052 4678 38054
rect 4382 37018 4438 37020
rect 4462 37018 4518 37020
rect 4542 37018 4598 37020
rect 4622 37018 4678 37020
rect 4382 36966 4428 37018
rect 4428 36966 4438 37018
rect 4462 36966 4492 37018
rect 4492 36966 4504 37018
rect 4504 36966 4518 37018
rect 4542 36966 4556 37018
rect 4556 36966 4568 37018
rect 4568 36966 4598 37018
rect 4622 36966 4632 37018
rect 4632 36966 4678 37018
rect 4382 36964 4438 36966
rect 4462 36964 4518 36966
rect 4542 36964 4598 36966
rect 4622 36964 4678 36966
rect 4382 35930 4438 35932
rect 4462 35930 4518 35932
rect 4542 35930 4598 35932
rect 4622 35930 4678 35932
rect 4382 35878 4428 35930
rect 4428 35878 4438 35930
rect 4462 35878 4492 35930
rect 4492 35878 4504 35930
rect 4504 35878 4518 35930
rect 4542 35878 4556 35930
rect 4556 35878 4568 35930
rect 4568 35878 4598 35930
rect 4622 35878 4632 35930
rect 4632 35878 4678 35930
rect 4382 35876 4438 35878
rect 4462 35876 4518 35878
rect 4542 35876 4598 35878
rect 4622 35876 4678 35878
rect 4382 34842 4438 34844
rect 4462 34842 4518 34844
rect 4542 34842 4598 34844
rect 4622 34842 4678 34844
rect 4382 34790 4428 34842
rect 4428 34790 4438 34842
rect 4462 34790 4492 34842
rect 4492 34790 4504 34842
rect 4504 34790 4518 34842
rect 4542 34790 4556 34842
rect 4556 34790 4568 34842
rect 4568 34790 4598 34842
rect 4622 34790 4632 34842
rect 4632 34790 4678 34842
rect 4382 34788 4438 34790
rect 4462 34788 4518 34790
rect 4542 34788 4598 34790
rect 4622 34788 4678 34790
rect 4382 33754 4438 33756
rect 4462 33754 4518 33756
rect 4542 33754 4598 33756
rect 4622 33754 4678 33756
rect 4382 33702 4428 33754
rect 4428 33702 4438 33754
rect 4462 33702 4492 33754
rect 4492 33702 4504 33754
rect 4504 33702 4518 33754
rect 4542 33702 4556 33754
rect 4556 33702 4568 33754
rect 4568 33702 4598 33754
rect 4622 33702 4632 33754
rect 4632 33702 4678 33754
rect 4382 33700 4438 33702
rect 4462 33700 4518 33702
rect 4542 33700 4598 33702
rect 4622 33700 4678 33702
rect 4382 32666 4438 32668
rect 4462 32666 4518 32668
rect 4542 32666 4598 32668
rect 4622 32666 4678 32668
rect 4382 32614 4428 32666
rect 4428 32614 4438 32666
rect 4462 32614 4492 32666
rect 4492 32614 4504 32666
rect 4504 32614 4518 32666
rect 4542 32614 4556 32666
rect 4556 32614 4568 32666
rect 4568 32614 4598 32666
rect 4622 32614 4632 32666
rect 4632 32614 4678 32666
rect 4382 32612 4438 32614
rect 4462 32612 4518 32614
rect 4542 32612 4598 32614
rect 4622 32612 4678 32614
rect 4382 31578 4438 31580
rect 4462 31578 4518 31580
rect 4542 31578 4598 31580
rect 4622 31578 4678 31580
rect 4382 31526 4428 31578
rect 4428 31526 4438 31578
rect 4462 31526 4492 31578
rect 4492 31526 4504 31578
rect 4504 31526 4518 31578
rect 4542 31526 4556 31578
rect 4556 31526 4568 31578
rect 4568 31526 4598 31578
rect 4622 31526 4632 31578
rect 4632 31526 4678 31578
rect 4382 31524 4438 31526
rect 4462 31524 4518 31526
rect 4542 31524 4598 31526
rect 4622 31524 4678 31526
rect 4382 30490 4438 30492
rect 4462 30490 4518 30492
rect 4542 30490 4598 30492
rect 4622 30490 4678 30492
rect 4382 30438 4428 30490
rect 4428 30438 4438 30490
rect 4462 30438 4492 30490
rect 4492 30438 4504 30490
rect 4504 30438 4518 30490
rect 4542 30438 4556 30490
rect 4556 30438 4568 30490
rect 4568 30438 4598 30490
rect 4622 30438 4632 30490
rect 4632 30438 4678 30490
rect 4382 30436 4438 30438
rect 4462 30436 4518 30438
rect 4542 30436 4598 30438
rect 4622 30436 4678 30438
rect 3698 18672 3754 18728
rect 4382 29402 4438 29404
rect 4462 29402 4518 29404
rect 4542 29402 4598 29404
rect 4622 29402 4678 29404
rect 4382 29350 4428 29402
rect 4428 29350 4438 29402
rect 4462 29350 4492 29402
rect 4492 29350 4504 29402
rect 4504 29350 4518 29402
rect 4542 29350 4556 29402
rect 4556 29350 4568 29402
rect 4568 29350 4598 29402
rect 4622 29350 4632 29402
rect 4632 29350 4678 29402
rect 4382 29348 4438 29350
rect 4462 29348 4518 29350
rect 4542 29348 4598 29350
rect 4622 29348 4678 29350
rect 3974 29144 4030 29200
rect 4382 28314 4438 28316
rect 4462 28314 4518 28316
rect 4542 28314 4598 28316
rect 4622 28314 4678 28316
rect 4382 28262 4428 28314
rect 4428 28262 4438 28314
rect 4462 28262 4492 28314
rect 4492 28262 4504 28314
rect 4504 28262 4518 28314
rect 4542 28262 4556 28314
rect 4556 28262 4568 28314
rect 4568 28262 4598 28314
rect 4622 28262 4632 28314
rect 4632 28262 4678 28314
rect 4382 28260 4438 28262
rect 4462 28260 4518 28262
rect 4542 28260 4598 28262
rect 4622 28260 4678 28262
rect 4382 27226 4438 27228
rect 4462 27226 4518 27228
rect 4542 27226 4598 27228
rect 4622 27226 4678 27228
rect 4382 27174 4428 27226
rect 4428 27174 4438 27226
rect 4462 27174 4492 27226
rect 4492 27174 4504 27226
rect 4504 27174 4518 27226
rect 4542 27174 4556 27226
rect 4556 27174 4568 27226
rect 4568 27174 4598 27226
rect 4622 27174 4632 27226
rect 4632 27174 4678 27226
rect 4382 27172 4438 27174
rect 4462 27172 4518 27174
rect 4542 27172 4598 27174
rect 4622 27172 4678 27174
rect 4382 26138 4438 26140
rect 4462 26138 4518 26140
rect 4542 26138 4598 26140
rect 4622 26138 4678 26140
rect 4382 26086 4428 26138
rect 4428 26086 4438 26138
rect 4462 26086 4492 26138
rect 4492 26086 4504 26138
rect 4504 26086 4518 26138
rect 4542 26086 4556 26138
rect 4556 26086 4568 26138
rect 4568 26086 4598 26138
rect 4622 26086 4632 26138
rect 4632 26086 4678 26138
rect 4382 26084 4438 26086
rect 4462 26084 4518 26086
rect 4542 26084 4598 26086
rect 4622 26084 4678 26086
rect 4382 25050 4438 25052
rect 4462 25050 4518 25052
rect 4542 25050 4598 25052
rect 4622 25050 4678 25052
rect 4382 24998 4428 25050
rect 4428 24998 4438 25050
rect 4462 24998 4492 25050
rect 4492 24998 4504 25050
rect 4504 24998 4518 25050
rect 4542 24998 4556 25050
rect 4556 24998 4568 25050
rect 4568 24998 4598 25050
rect 4622 24998 4632 25050
rect 4632 24998 4678 25050
rect 4382 24996 4438 24998
rect 4462 24996 4518 24998
rect 4542 24996 4598 24998
rect 4622 24996 4678 24998
rect 4382 23962 4438 23964
rect 4462 23962 4518 23964
rect 4542 23962 4598 23964
rect 4622 23962 4678 23964
rect 4382 23910 4428 23962
rect 4428 23910 4438 23962
rect 4462 23910 4492 23962
rect 4492 23910 4504 23962
rect 4504 23910 4518 23962
rect 4542 23910 4556 23962
rect 4556 23910 4568 23962
rect 4568 23910 4598 23962
rect 4622 23910 4632 23962
rect 4632 23910 4678 23962
rect 4382 23908 4438 23910
rect 4462 23908 4518 23910
rect 4542 23908 4598 23910
rect 4622 23908 4678 23910
rect 4382 22874 4438 22876
rect 4462 22874 4518 22876
rect 4542 22874 4598 22876
rect 4622 22874 4678 22876
rect 4382 22822 4428 22874
rect 4428 22822 4438 22874
rect 4462 22822 4492 22874
rect 4492 22822 4504 22874
rect 4504 22822 4518 22874
rect 4542 22822 4556 22874
rect 4556 22822 4568 22874
rect 4568 22822 4598 22874
rect 4622 22822 4632 22874
rect 4632 22822 4678 22874
rect 4382 22820 4438 22822
rect 4462 22820 4518 22822
rect 4542 22820 4598 22822
rect 4622 22820 4678 22822
rect 4382 21786 4438 21788
rect 4462 21786 4518 21788
rect 4542 21786 4598 21788
rect 4622 21786 4678 21788
rect 4382 21734 4428 21786
rect 4428 21734 4438 21786
rect 4462 21734 4492 21786
rect 4492 21734 4504 21786
rect 4504 21734 4518 21786
rect 4542 21734 4556 21786
rect 4556 21734 4568 21786
rect 4568 21734 4598 21786
rect 4622 21734 4632 21786
rect 4632 21734 4678 21786
rect 4382 21732 4438 21734
rect 4462 21732 4518 21734
rect 4542 21732 4598 21734
rect 4622 21732 4678 21734
rect 4382 20698 4438 20700
rect 4462 20698 4518 20700
rect 4542 20698 4598 20700
rect 4622 20698 4678 20700
rect 4382 20646 4428 20698
rect 4428 20646 4438 20698
rect 4462 20646 4492 20698
rect 4492 20646 4504 20698
rect 4504 20646 4518 20698
rect 4542 20646 4556 20698
rect 4556 20646 4568 20698
rect 4568 20646 4598 20698
rect 4622 20646 4632 20698
rect 4632 20646 4678 20698
rect 4382 20644 4438 20646
rect 4462 20644 4518 20646
rect 4542 20644 4598 20646
rect 4622 20644 4678 20646
rect 4382 19610 4438 19612
rect 4462 19610 4518 19612
rect 4542 19610 4598 19612
rect 4622 19610 4678 19612
rect 4382 19558 4428 19610
rect 4428 19558 4438 19610
rect 4462 19558 4492 19610
rect 4492 19558 4504 19610
rect 4504 19558 4518 19610
rect 4542 19558 4556 19610
rect 4556 19558 4568 19610
rect 4568 19558 4598 19610
rect 4622 19558 4632 19610
rect 4632 19558 4678 19610
rect 4382 19556 4438 19558
rect 4462 19556 4518 19558
rect 4542 19556 4598 19558
rect 4622 19556 4678 19558
rect 4382 18522 4438 18524
rect 4462 18522 4518 18524
rect 4542 18522 4598 18524
rect 4622 18522 4678 18524
rect 4382 18470 4428 18522
rect 4428 18470 4438 18522
rect 4462 18470 4492 18522
rect 4492 18470 4504 18522
rect 4504 18470 4518 18522
rect 4542 18470 4556 18522
rect 4556 18470 4568 18522
rect 4568 18470 4598 18522
rect 4622 18470 4632 18522
rect 4632 18470 4678 18522
rect 4382 18468 4438 18470
rect 4462 18468 4518 18470
rect 4542 18468 4598 18470
rect 4622 18468 4678 18470
rect 4382 17434 4438 17436
rect 4462 17434 4518 17436
rect 4542 17434 4598 17436
rect 4622 17434 4678 17436
rect 4382 17382 4428 17434
rect 4428 17382 4438 17434
rect 4462 17382 4492 17434
rect 4492 17382 4504 17434
rect 4504 17382 4518 17434
rect 4542 17382 4556 17434
rect 4556 17382 4568 17434
rect 4568 17382 4598 17434
rect 4622 17382 4632 17434
rect 4632 17382 4678 17434
rect 4382 17380 4438 17382
rect 4462 17380 4518 17382
rect 4542 17380 4598 17382
rect 4622 17380 4678 17382
rect 4382 16346 4438 16348
rect 4462 16346 4518 16348
rect 4542 16346 4598 16348
rect 4622 16346 4678 16348
rect 4382 16294 4428 16346
rect 4428 16294 4438 16346
rect 4462 16294 4492 16346
rect 4492 16294 4504 16346
rect 4504 16294 4518 16346
rect 4542 16294 4556 16346
rect 4556 16294 4568 16346
rect 4568 16294 4598 16346
rect 4622 16294 4632 16346
rect 4632 16294 4678 16346
rect 4382 16292 4438 16294
rect 4462 16292 4518 16294
rect 4542 16292 4598 16294
rect 4622 16292 4678 16294
rect 4382 15258 4438 15260
rect 4462 15258 4518 15260
rect 4542 15258 4598 15260
rect 4622 15258 4678 15260
rect 4382 15206 4428 15258
rect 4428 15206 4438 15258
rect 4462 15206 4492 15258
rect 4492 15206 4504 15258
rect 4504 15206 4518 15258
rect 4542 15206 4556 15258
rect 4556 15206 4568 15258
rect 4568 15206 4598 15258
rect 4622 15206 4632 15258
rect 4632 15206 4678 15258
rect 4382 15204 4438 15206
rect 4462 15204 4518 15206
rect 4542 15204 4598 15206
rect 4622 15204 4678 15206
rect 4382 14170 4438 14172
rect 4462 14170 4518 14172
rect 4542 14170 4598 14172
rect 4622 14170 4678 14172
rect 4382 14118 4428 14170
rect 4428 14118 4438 14170
rect 4462 14118 4492 14170
rect 4492 14118 4504 14170
rect 4504 14118 4518 14170
rect 4542 14118 4556 14170
rect 4556 14118 4568 14170
rect 4568 14118 4598 14170
rect 4622 14118 4632 14170
rect 4632 14118 4678 14170
rect 4382 14116 4438 14118
rect 4462 14116 4518 14118
rect 4542 14116 4598 14118
rect 4622 14116 4678 14118
rect 4382 13082 4438 13084
rect 4462 13082 4518 13084
rect 4542 13082 4598 13084
rect 4622 13082 4678 13084
rect 4382 13030 4428 13082
rect 4428 13030 4438 13082
rect 4462 13030 4492 13082
rect 4492 13030 4504 13082
rect 4504 13030 4518 13082
rect 4542 13030 4556 13082
rect 4556 13030 4568 13082
rect 4568 13030 4598 13082
rect 4622 13030 4632 13082
rect 4632 13030 4678 13082
rect 4382 13028 4438 13030
rect 4462 13028 4518 13030
rect 4542 13028 4598 13030
rect 4622 13028 4678 13030
rect 4382 11994 4438 11996
rect 4462 11994 4518 11996
rect 4542 11994 4598 11996
rect 4622 11994 4678 11996
rect 4382 11942 4428 11994
rect 4428 11942 4438 11994
rect 4462 11942 4492 11994
rect 4492 11942 4504 11994
rect 4504 11942 4518 11994
rect 4542 11942 4556 11994
rect 4556 11942 4568 11994
rect 4568 11942 4598 11994
rect 4622 11942 4632 11994
rect 4632 11942 4678 11994
rect 4382 11940 4438 11942
rect 4462 11940 4518 11942
rect 4542 11940 4598 11942
rect 4622 11940 4678 11942
rect 4382 10906 4438 10908
rect 4462 10906 4518 10908
rect 4542 10906 4598 10908
rect 4622 10906 4678 10908
rect 4382 10854 4428 10906
rect 4428 10854 4438 10906
rect 4462 10854 4492 10906
rect 4492 10854 4504 10906
rect 4504 10854 4518 10906
rect 4542 10854 4556 10906
rect 4556 10854 4568 10906
rect 4568 10854 4598 10906
rect 4622 10854 4632 10906
rect 4632 10854 4678 10906
rect 4382 10852 4438 10854
rect 4462 10852 4518 10854
rect 4542 10852 4598 10854
rect 4622 10852 4678 10854
rect 4382 9818 4438 9820
rect 4462 9818 4518 9820
rect 4542 9818 4598 9820
rect 4622 9818 4678 9820
rect 4382 9766 4428 9818
rect 4428 9766 4438 9818
rect 4462 9766 4492 9818
rect 4492 9766 4504 9818
rect 4504 9766 4518 9818
rect 4542 9766 4556 9818
rect 4556 9766 4568 9818
rect 4568 9766 4598 9818
rect 4622 9766 4632 9818
rect 4632 9766 4678 9818
rect 4382 9764 4438 9766
rect 4462 9764 4518 9766
rect 4542 9764 4598 9766
rect 4622 9764 4678 9766
rect 4382 8730 4438 8732
rect 4462 8730 4518 8732
rect 4542 8730 4598 8732
rect 4622 8730 4678 8732
rect 4382 8678 4428 8730
rect 4428 8678 4438 8730
rect 4462 8678 4492 8730
rect 4492 8678 4504 8730
rect 4504 8678 4518 8730
rect 4542 8678 4556 8730
rect 4556 8678 4568 8730
rect 4568 8678 4598 8730
rect 4622 8678 4632 8730
rect 4632 8678 4678 8730
rect 4382 8676 4438 8678
rect 4462 8676 4518 8678
rect 4542 8676 4598 8678
rect 4622 8676 4678 8678
rect 5446 35536 5502 35592
rect 6096 37562 6152 37564
rect 6176 37562 6232 37564
rect 6256 37562 6312 37564
rect 6336 37562 6392 37564
rect 6096 37510 6142 37562
rect 6142 37510 6152 37562
rect 6176 37510 6206 37562
rect 6206 37510 6218 37562
rect 6218 37510 6232 37562
rect 6256 37510 6270 37562
rect 6270 37510 6282 37562
rect 6282 37510 6312 37562
rect 6336 37510 6346 37562
rect 6346 37510 6392 37562
rect 6096 37508 6152 37510
rect 6176 37508 6232 37510
rect 6256 37508 6312 37510
rect 6336 37508 6392 37510
rect 6096 36474 6152 36476
rect 6176 36474 6232 36476
rect 6256 36474 6312 36476
rect 6336 36474 6392 36476
rect 6096 36422 6142 36474
rect 6142 36422 6152 36474
rect 6176 36422 6206 36474
rect 6206 36422 6218 36474
rect 6218 36422 6232 36474
rect 6256 36422 6270 36474
rect 6270 36422 6282 36474
rect 6282 36422 6312 36474
rect 6336 36422 6346 36474
rect 6346 36422 6392 36474
rect 6096 36420 6152 36422
rect 6176 36420 6232 36422
rect 6256 36420 6312 36422
rect 6336 36420 6392 36422
rect 6096 35386 6152 35388
rect 6176 35386 6232 35388
rect 6256 35386 6312 35388
rect 6336 35386 6392 35388
rect 6096 35334 6142 35386
rect 6142 35334 6152 35386
rect 6176 35334 6206 35386
rect 6206 35334 6218 35386
rect 6218 35334 6232 35386
rect 6256 35334 6270 35386
rect 6270 35334 6282 35386
rect 6282 35334 6312 35386
rect 6336 35334 6346 35386
rect 6346 35334 6392 35386
rect 6096 35332 6152 35334
rect 6176 35332 6232 35334
rect 6256 35332 6312 35334
rect 6336 35332 6392 35334
rect 5262 20440 5318 20496
rect 5446 19896 5502 19952
rect 5262 13368 5318 13424
rect 6096 34298 6152 34300
rect 6176 34298 6232 34300
rect 6256 34298 6312 34300
rect 6336 34298 6392 34300
rect 6096 34246 6142 34298
rect 6142 34246 6152 34298
rect 6176 34246 6206 34298
rect 6206 34246 6218 34298
rect 6218 34246 6232 34298
rect 6256 34246 6270 34298
rect 6270 34246 6282 34298
rect 6282 34246 6312 34298
rect 6336 34246 6346 34298
rect 6346 34246 6392 34298
rect 6096 34244 6152 34246
rect 6176 34244 6232 34246
rect 6256 34244 6312 34246
rect 6336 34244 6392 34246
rect 6096 33210 6152 33212
rect 6176 33210 6232 33212
rect 6256 33210 6312 33212
rect 6336 33210 6392 33212
rect 6096 33158 6142 33210
rect 6142 33158 6152 33210
rect 6176 33158 6206 33210
rect 6206 33158 6218 33210
rect 6218 33158 6232 33210
rect 6256 33158 6270 33210
rect 6270 33158 6282 33210
rect 6282 33158 6312 33210
rect 6336 33158 6346 33210
rect 6346 33158 6392 33210
rect 6096 33156 6152 33158
rect 6176 33156 6232 33158
rect 6256 33156 6312 33158
rect 6336 33156 6392 33158
rect 6096 32122 6152 32124
rect 6176 32122 6232 32124
rect 6256 32122 6312 32124
rect 6336 32122 6392 32124
rect 6096 32070 6142 32122
rect 6142 32070 6152 32122
rect 6176 32070 6206 32122
rect 6206 32070 6218 32122
rect 6218 32070 6232 32122
rect 6256 32070 6270 32122
rect 6270 32070 6282 32122
rect 6282 32070 6312 32122
rect 6336 32070 6346 32122
rect 6346 32070 6392 32122
rect 6096 32068 6152 32070
rect 6176 32068 6232 32070
rect 6256 32068 6312 32070
rect 6336 32068 6392 32070
rect 6096 31034 6152 31036
rect 6176 31034 6232 31036
rect 6256 31034 6312 31036
rect 6336 31034 6392 31036
rect 6096 30982 6142 31034
rect 6142 30982 6152 31034
rect 6176 30982 6206 31034
rect 6206 30982 6218 31034
rect 6218 30982 6232 31034
rect 6256 30982 6270 31034
rect 6270 30982 6282 31034
rect 6282 30982 6312 31034
rect 6336 30982 6346 31034
rect 6346 30982 6392 31034
rect 6096 30980 6152 30982
rect 6176 30980 6232 30982
rect 6256 30980 6312 30982
rect 6336 30980 6392 30982
rect 6096 29946 6152 29948
rect 6176 29946 6232 29948
rect 6256 29946 6312 29948
rect 6336 29946 6392 29948
rect 6096 29894 6142 29946
rect 6142 29894 6152 29946
rect 6176 29894 6206 29946
rect 6206 29894 6218 29946
rect 6218 29894 6232 29946
rect 6256 29894 6270 29946
rect 6270 29894 6282 29946
rect 6282 29894 6312 29946
rect 6336 29894 6346 29946
rect 6346 29894 6392 29946
rect 6096 29892 6152 29894
rect 6176 29892 6232 29894
rect 6256 29892 6312 29894
rect 6336 29892 6392 29894
rect 6096 28858 6152 28860
rect 6176 28858 6232 28860
rect 6256 28858 6312 28860
rect 6336 28858 6392 28860
rect 6096 28806 6142 28858
rect 6142 28806 6152 28858
rect 6176 28806 6206 28858
rect 6206 28806 6218 28858
rect 6218 28806 6232 28858
rect 6256 28806 6270 28858
rect 6270 28806 6282 28858
rect 6282 28806 6312 28858
rect 6336 28806 6346 28858
rect 6346 28806 6392 28858
rect 6096 28804 6152 28806
rect 6176 28804 6232 28806
rect 6256 28804 6312 28806
rect 6336 28804 6392 28806
rect 6096 27770 6152 27772
rect 6176 27770 6232 27772
rect 6256 27770 6312 27772
rect 6336 27770 6392 27772
rect 6096 27718 6142 27770
rect 6142 27718 6152 27770
rect 6176 27718 6206 27770
rect 6206 27718 6218 27770
rect 6218 27718 6232 27770
rect 6256 27718 6270 27770
rect 6270 27718 6282 27770
rect 6282 27718 6312 27770
rect 6336 27718 6346 27770
rect 6346 27718 6392 27770
rect 6096 27716 6152 27718
rect 6176 27716 6232 27718
rect 6256 27716 6312 27718
rect 6336 27716 6392 27718
rect 7286 41520 7342 41576
rect 12438 41520 12494 41576
rect 7809 41370 7865 41372
rect 7889 41370 7945 41372
rect 7969 41370 8025 41372
rect 8049 41370 8105 41372
rect 7809 41318 7855 41370
rect 7855 41318 7865 41370
rect 7889 41318 7919 41370
rect 7919 41318 7931 41370
rect 7931 41318 7945 41370
rect 7969 41318 7983 41370
rect 7983 41318 7995 41370
rect 7995 41318 8025 41370
rect 8049 41318 8059 41370
rect 8059 41318 8105 41370
rect 7809 41316 7865 41318
rect 7889 41316 7945 41318
rect 7969 41316 8025 41318
rect 8049 41316 8105 41318
rect 11236 41370 11292 41372
rect 11316 41370 11372 41372
rect 11396 41370 11452 41372
rect 11476 41370 11532 41372
rect 11236 41318 11282 41370
rect 11282 41318 11292 41370
rect 11316 41318 11346 41370
rect 11346 41318 11358 41370
rect 11358 41318 11372 41370
rect 11396 41318 11410 41370
rect 11410 41318 11422 41370
rect 11422 41318 11452 41370
rect 11476 41318 11486 41370
rect 11486 41318 11532 41370
rect 11236 41316 11292 41318
rect 11316 41316 11372 41318
rect 11396 41316 11452 41318
rect 11476 41316 11532 41318
rect 14663 41370 14719 41372
rect 14743 41370 14799 41372
rect 14823 41370 14879 41372
rect 14903 41370 14959 41372
rect 14663 41318 14709 41370
rect 14709 41318 14719 41370
rect 14743 41318 14773 41370
rect 14773 41318 14785 41370
rect 14785 41318 14799 41370
rect 14823 41318 14837 41370
rect 14837 41318 14849 41370
rect 14849 41318 14879 41370
rect 14903 41318 14913 41370
rect 14913 41318 14959 41370
rect 14663 41316 14719 41318
rect 14743 41316 14799 41318
rect 14823 41316 14879 41318
rect 14903 41316 14959 41318
rect 7809 40282 7865 40284
rect 7889 40282 7945 40284
rect 7969 40282 8025 40284
rect 8049 40282 8105 40284
rect 7809 40230 7855 40282
rect 7855 40230 7865 40282
rect 7889 40230 7919 40282
rect 7919 40230 7931 40282
rect 7931 40230 7945 40282
rect 7969 40230 7983 40282
rect 7983 40230 7995 40282
rect 7995 40230 8025 40282
rect 8049 40230 8059 40282
rect 8059 40230 8105 40282
rect 7809 40228 7865 40230
rect 7889 40228 7945 40230
rect 7969 40228 8025 40230
rect 8049 40228 8105 40230
rect 9523 40826 9579 40828
rect 9603 40826 9659 40828
rect 9683 40826 9739 40828
rect 9763 40826 9819 40828
rect 9523 40774 9569 40826
rect 9569 40774 9579 40826
rect 9603 40774 9633 40826
rect 9633 40774 9645 40826
rect 9645 40774 9659 40826
rect 9683 40774 9697 40826
rect 9697 40774 9709 40826
rect 9709 40774 9739 40826
rect 9763 40774 9773 40826
rect 9773 40774 9819 40826
rect 9523 40772 9579 40774
rect 9603 40772 9659 40774
rect 9683 40772 9739 40774
rect 9763 40772 9819 40774
rect 12950 40826 13006 40828
rect 13030 40826 13086 40828
rect 13110 40826 13166 40828
rect 13190 40826 13246 40828
rect 12950 40774 12996 40826
rect 12996 40774 13006 40826
rect 13030 40774 13060 40826
rect 13060 40774 13072 40826
rect 13072 40774 13086 40826
rect 13110 40774 13124 40826
rect 13124 40774 13136 40826
rect 13136 40774 13166 40826
rect 13190 40774 13200 40826
rect 13200 40774 13246 40826
rect 12950 40772 13006 40774
rect 13030 40772 13086 40774
rect 13110 40772 13166 40774
rect 13190 40772 13246 40774
rect 11236 40282 11292 40284
rect 11316 40282 11372 40284
rect 11396 40282 11452 40284
rect 11476 40282 11532 40284
rect 11236 40230 11282 40282
rect 11282 40230 11292 40282
rect 11316 40230 11346 40282
rect 11346 40230 11358 40282
rect 11358 40230 11372 40282
rect 11396 40230 11410 40282
rect 11410 40230 11422 40282
rect 11422 40230 11452 40282
rect 11476 40230 11486 40282
rect 11486 40230 11532 40282
rect 11236 40228 11292 40230
rect 11316 40228 11372 40230
rect 11396 40228 11452 40230
rect 11476 40228 11532 40230
rect 14663 40282 14719 40284
rect 14743 40282 14799 40284
rect 14823 40282 14879 40284
rect 14903 40282 14959 40284
rect 14663 40230 14709 40282
rect 14709 40230 14719 40282
rect 14743 40230 14773 40282
rect 14773 40230 14785 40282
rect 14785 40230 14799 40282
rect 14823 40230 14837 40282
rect 14837 40230 14849 40282
rect 14849 40230 14879 40282
rect 14903 40230 14913 40282
rect 14913 40230 14959 40282
rect 14663 40228 14719 40230
rect 14743 40228 14799 40230
rect 14823 40228 14879 40230
rect 14903 40228 14959 40230
rect 9523 39738 9579 39740
rect 9603 39738 9659 39740
rect 9683 39738 9739 39740
rect 9763 39738 9819 39740
rect 9523 39686 9569 39738
rect 9569 39686 9579 39738
rect 9603 39686 9633 39738
rect 9633 39686 9645 39738
rect 9645 39686 9659 39738
rect 9683 39686 9697 39738
rect 9697 39686 9709 39738
rect 9709 39686 9739 39738
rect 9763 39686 9773 39738
rect 9773 39686 9819 39738
rect 9523 39684 9579 39686
rect 9603 39684 9659 39686
rect 9683 39684 9739 39686
rect 9763 39684 9819 39686
rect 12950 39738 13006 39740
rect 13030 39738 13086 39740
rect 13110 39738 13166 39740
rect 13190 39738 13246 39740
rect 12950 39686 12996 39738
rect 12996 39686 13006 39738
rect 13030 39686 13060 39738
rect 13060 39686 13072 39738
rect 13072 39686 13086 39738
rect 13110 39686 13124 39738
rect 13124 39686 13136 39738
rect 13136 39686 13166 39738
rect 13190 39686 13200 39738
rect 13200 39686 13246 39738
rect 12950 39684 13006 39686
rect 13030 39684 13086 39686
rect 13110 39684 13166 39686
rect 13190 39684 13246 39686
rect 14002 39480 14058 39536
rect 14186 39480 14242 39536
rect 7286 37168 7342 37224
rect 6096 26682 6152 26684
rect 6176 26682 6232 26684
rect 6256 26682 6312 26684
rect 6336 26682 6392 26684
rect 6096 26630 6142 26682
rect 6142 26630 6152 26682
rect 6176 26630 6206 26682
rect 6206 26630 6218 26682
rect 6218 26630 6232 26682
rect 6256 26630 6270 26682
rect 6270 26630 6282 26682
rect 6282 26630 6312 26682
rect 6336 26630 6346 26682
rect 6346 26630 6392 26682
rect 6096 26628 6152 26630
rect 6176 26628 6232 26630
rect 6256 26628 6312 26630
rect 6336 26628 6392 26630
rect 6096 25594 6152 25596
rect 6176 25594 6232 25596
rect 6256 25594 6312 25596
rect 6336 25594 6392 25596
rect 6096 25542 6142 25594
rect 6142 25542 6152 25594
rect 6176 25542 6206 25594
rect 6206 25542 6218 25594
rect 6218 25542 6232 25594
rect 6256 25542 6270 25594
rect 6270 25542 6282 25594
rect 6282 25542 6312 25594
rect 6336 25542 6346 25594
rect 6346 25542 6392 25594
rect 6096 25540 6152 25542
rect 6176 25540 6232 25542
rect 6256 25540 6312 25542
rect 6336 25540 6392 25542
rect 6096 24506 6152 24508
rect 6176 24506 6232 24508
rect 6256 24506 6312 24508
rect 6336 24506 6392 24508
rect 6096 24454 6142 24506
rect 6142 24454 6152 24506
rect 6176 24454 6206 24506
rect 6206 24454 6218 24506
rect 6218 24454 6232 24506
rect 6256 24454 6270 24506
rect 6270 24454 6282 24506
rect 6282 24454 6312 24506
rect 6336 24454 6346 24506
rect 6346 24454 6392 24506
rect 6096 24452 6152 24454
rect 6176 24452 6232 24454
rect 6256 24452 6312 24454
rect 6336 24452 6392 24454
rect 6096 23418 6152 23420
rect 6176 23418 6232 23420
rect 6256 23418 6312 23420
rect 6336 23418 6392 23420
rect 6096 23366 6142 23418
rect 6142 23366 6152 23418
rect 6176 23366 6206 23418
rect 6206 23366 6218 23418
rect 6218 23366 6232 23418
rect 6256 23366 6270 23418
rect 6270 23366 6282 23418
rect 6282 23366 6312 23418
rect 6336 23366 6346 23418
rect 6346 23366 6392 23418
rect 6096 23364 6152 23366
rect 6176 23364 6232 23366
rect 6256 23364 6312 23366
rect 6336 23364 6392 23366
rect 6096 22330 6152 22332
rect 6176 22330 6232 22332
rect 6256 22330 6312 22332
rect 6336 22330 6392 22332
rect 6096 22278 6142 22330
rect 6142 22278 6152 22330
rect 6176 22278 6206 22330
rect 6206 22278 6218 22330
rect 6218 22278 6232 22330
rect 6256 22278 6270 22330
rect 6270 22278 6282 22330
rect 6282 22278 6312 22330
rect 6336 22278 6346 22330
rect 6346 22278 6392 22330
rect 6096 22276 6152 22278
rect 6176 22276 6232 22278
rect 6256 22276 6312 22278
rect 6336 22276 6392 22278
rect 6096 21242 6152 21244
rect 6176 21242 6232 21244
rect 6256 21242 6312 21244
rect 6336 21242 6392 21244
rect 6096 21190 6142 21242
rect 6142 21190 6152 21242
rect 6176 21190 6206 21242
rect 6206 21190 6218 21242
rect 6218 21190 6232 21242
rect 6256 21190 6270 21242
rect 6270 21190 6282 21242
rect 6282 21190 6312 21242
rect 6336 21190 6346 21242
rect 6346 21190 6392 21242
rect 6096 21188 6152 21190
rect 6176 21188 6232 21190
rect 6256 21188 6312 21190
rect 6336 21188 6392 21190
rect 6096 20154 6152 20156
rect 6176 20154 6232 20156
rect 6256 20154 6312 20156
rect 6336 20154 6392 20156
rect 6096 20102 6142 20154
rect 6142 20102 6152 20154
rect 6176 20102 6206 20154
rect 6206 20102 6218 20154
rect 6218 20102 6232 20154
rect 6256 20102 6270 20154
rect 6270 20102 6282 20154
rect 6282 20102 6312 20154
rect 6336 20102 6346 20154
rect 6346 20102 6392 20154
rect 6096 20100 6152 20102
rect 6176 20100 6232 20102
rect 6256 20100 6312 20102
rect 6336 20100 6392 20102
rect 6096 19066 6152 19068
rect 6176 19066 6232 19068
rect 6256 19066 6312 19068
rect 6336 19066 6392 19068
rect 6096 19014 6142 19066
rect 6142 19014 6152 19066
rect 6176 19014 6206 19066
rect 6206 19014 6218 19066
rect 6218 19014 6232 19066
rect 6256 19014 6270 19066
rect 6270 19014 6282 19066
rect 6282 19014 6312 19066
rect 6336 19014 6346 19066
rect 6346 19014 6392 19066
rect 6096 19012 6152 19014
rect 6176 19012 6232 19014
rect 6256 19012 6312 19014
rect 6336 19012 6392 19014
rect 6090 18672 6146 18728
rect 6096 17978 6152 17980
rect 6176 17978 6232 17980
rect 6256 17978 6312 17980
rect 6336 17978 6392 17980
rect 6096 17926 6142 17978
rect 6142 17926 6152 17978
rect 6176 17926 6206 17978
rect 6206 17926 6218 17978
rect 6218 17926 6232 17978
rect 6256 17926 6270 17978
rect 6270 17926 6282 17978
rect 6282 17926 6312 17978
rect 6336 17926 6346 17978
rect 6346 17926 6392 17978
rect 6096 17924 6152 17926
rect 6176 17924 6232 17926
rect 6256 17924 6312 17926
rect 6336 17924 6392 17926
rect 5906 12144 5962 12200
rect 4986 9696 5042 9752
rect 5722 9696 5778 9752
rect 4382 7642 4438 7644
rect 4462 7642 4518 7644
rect 4542 7642 4598 7644
rect 4622 7642 4678 7644
rect 4382 7590 4428 7642
rect 4428 7590 4438 7642
rect 4462 7590 4492 7642
rect 4492 7590 4504 7642
rect 4504 7590 4518 7642
rect 4542 7590 4556 7642
rect 4556 7590 4568 7642
rect 4568 7590 4598 7642
rect 4622 7590 4632 7642
rect 4632 7590 4678 7642
rect 4382 7588 4438 7590
rect 4462 7588 4518 7590
rect 4542 7588 4598 7590
rect 4622 7588 4678 7590
rect 4382 6554 4438 6556
rect 4462 6554 4518 6556
rect 4542 6554 4598 6556
rect 4622 6554 4678 6556
rect 4382 6502 4428 6554
rect 4428 6502 4438 6554
rect 4462 6502 4492 6554
rect 4492 6502 4504 6554
rect 4504 6502 4518 6554
rect 4542 6502 4556 6554
rect 4556 6502 4568 6554
rect 4568 6502 4598 6554
rect 4622 6502 4632 6554
rect 4632 6502 4678 6554
rect 4382 6500 4438 6502
rect 4462 6500 4518 6502
rect 4542 6500 4598 6502
rect 4622 6500 4678 6502
rect 6096 16890 6152 16892
rect 6176 16890 6232 16892
rect 6256 16890 6312 16892
rect 6336 16890 6392 16892
rect 6096 16838 6142 16890
rect 6142 16838 6152 16890
rect 6176 16838 6206 16890
rect 6206 16838 6218 16890
rect 6218 16838 6232 16890
rect 6256 16838 6270 16890
rect 6270 16838 6282 16890
rect 6282 16838 6312 16890
rect 6336 16838 6346 16890
rect 6346 16838 6392 16890
rect 6096 16836 6152 16838
rect 6176 16836 6232 16838
rect 6256 16836 6312 16838
rect 6336 16836 6392 16838
rect 6096 15802 6152 15804
rect 6176 15802 6232 15804
rect 6256 15802 6312 15804
rect 6336 15802 6392 15804
rect 6096 15750 6142 15802
rect 6142 15750 6152 15802
rect 6176 15750 6206 15802
rect 6206 15750 6218 15802
rect 6218 15750 6232 15802
rect 6256 15750 6270 15802
rect 6270 15750 6282 15802
rect 6282 15750 6312 15802
rect 6336 15750 6346 15802
rect 6346 15750 6392 15802
rect 6096 15748 6152 15750
rect 6176 15748 6232 15750
rect 6256 15748 6312 15750
rect 6336 15748 6392 15750
rect 6096 14714 6152 14716
rect 6176 14714 6232 14716
rect 6256 14714 6312 14716
rect 6336 14714 6392 14716
rect 6096 14662 6142 14714
rect 6142 14662 6152 14714
rect 6176 14662 6206 14714
rect 6206 14662 6218 14714
rect 6218 14662 6232 14714
rect 6256 14662 6270 14714
rect 6270 14662 6282 14714
rect 6282 14662 6312 14714
rect 6336 14662 6346 14714
rect 6346 14662 6392 14714
rect 6096 14660 6152 14662
rect 6176 14660 6232 14662
rect 6256 14660 6312 14662
rect 6336 14660 6392 14662
rect 7809 39194 7865 39196
rect 7889 39194 7945 39196
rect 7969 39194 8025 39196
rect 8049 39194 8105 39196
rect 7809 39142 7855 39194
rect 7855 39142 7865 39194
rect 7889 39142 7919 39194
rect 7919 39142 7931 39194
rect 7931 39142 7945 39194
rect 7969 39142 7983 39194
rect 7983 39142 7995 39194
rect 7995 39142 8025 39194
rect 8049 39142 8059 39194
rect 8059 39142 8105 39194
rect 7809 39140 7865 39142
rect 7889 39140 7945 39142
rect 7969 39140 8025 39142
rect 8049 39140 8105 39142
rect 7809 38106 7865 38108
rect 7889 38106 7945 38108
rect 7969 38106 8025 38108
rect 8049 38106 8105 38108
rect 7809 38054 7855 38106
rect 7855 38054 7865 38106
rect 7889 38054 7919 38106
rect 7919 38054 7931 38106
rect 7931 38054 7945 38106
rect 7969 38054 7983 38106
rect 7983 38054 7995 38106
rect 7995 38054 8025 38106
rect 8049 38054 8059 38106
rect 8059 38054 8105 38106
rect 7809 38052 7865 38054
rect 7889 38052 7945 38054
rect 7969 38052 8025 38054
rect 8049 38052 8105 38054
rect 7809 37018 7865 37020
rect 7889 37018 7945 37020
rect 7969 37018 8025 37020
rect 8049 37018 8105 37020
rect 7809 36966 7855 37018
rect 7855 36966 7865 37018
rect 7889 36966 7919 37018
rect 7919 36966 7931 37018
rect 7931 36966 7945 37018
rect 7969 36966 7983 37018
rect 7983 36966 7995 37018
rect 7995 36966 8025 37018
rect 8049 36966 8059 37018
rect 8059 36966 8105 37018
rect 7809 36964 7865 36966
rect 7889 36964 7945 36966
rect 7969 36964 8025 36966
rect 8049 36964 8105 36966
rect 7809 35930 7865 35932
rect 7889 35930 7945 35932
rect 7969 35930 8025 35932
rect 8049 35930 8105 35932
rect 7809 35878 7855 35930
rect 7855 35878 7865 35930
rect 7889 35878 7919 35930
rect 7919 35878 7931 35930
rect 7931 35878 7945 35930
rect 7969 35878 7983 35930
rect 7983 35878 7995 35930
rect 7995 35878 8025 35930
rect 8049 35878 8059 35930
rect 8059 35878 8105 35930
rect 7809 35876 7865 35878
rect 7889 35876 7945 35878
rect 7969 35876 8025 35878
rect 8049 35876 8105 35878
rect 7809 34842 7865 34844
rect 7889 34842 7945 34844
rect 7969 34842 8025 34844
rect 8049 34842 8105 34844
rect 7809 34790 7855 34842
rect 7855 34790 7865 34842
rect 7889 34790 7919 34842
rect 7919 34790 7931 34842
rect 7931 34790 7945 34842
rect 7969 34790 7983 34842
rect 7983 34790 7995 34842
rect 7995 34790 8025 34842
rect 8049 34790 8059 34842
rect 8059 34790 8105 34842
rect 7809 34788 7865 34790
rect 7889 34788 7945 34790
rect 7969 34788 8025 34790
rect 8049 34788 8105 34790
rect 7809 33754 7865 33756
rect 7889 33754 7945 33756
rect 7969 33754 8025 33756
rect 8049 33754 8105 33756
rect 7809 33702 7855 33754
rect 7855 33702 7865 33754
rect 7889 33702 7919 33754
rect 7919 33702 7931 33754
rect 7931 33702 7945 33754
rect 7969 33702 7983 33754
rect 7983 33702 7995 33754
rect 7995 33702 8025 33754
rect 8049 33702 8059 33754
rect 8059 33702 8105 33754
rect 7809 33700 7865 33702
rect 7889 33700 7945 33702
rect 7969 33700 8025 33702
rect 8049 33700 8105 33702
rect 7809 32666 7865 32668
rect 7889 32666 7945 32668
rect 7969 32666 8025 32668
rect 8049 32666 8105 32668
rect 7809 32614 7855 32666
rect 7855 32614 7865 32666
rect 7889 32614 7919 32666
rect 7919 32614 7931 32666
rect 7931 32614 7945 32666
rect 7969 32614 7983 32666
rect 7983 32614 7995 32666
rect 7995 32614 8025 32666
rect 8049 32614 8059 32666
rect 8059 32614 8105 32666
rect 7809 32612 7865 32614
rect 7889 32612 7945 32614
rect 7969 32612 8025 32614
rect 8049 32612 8105 32614
rect 11236 39194 11292 39196
rect 11316 39194 11372 39196
rect 11396 39194 11452 39196
rect 11476 39194 11532 39196
rect 11236 39142 11282 39194
rect 11282 39142 11292 39194
rect 11316 39142 11346 39194
rect 11346 39142 11358 39194
rect 11358 39142 11372 39194
rect 11396 39142 11410 39194
rect 11410 39142 11422 39194
rect 11422 39142 11452 39194
rect 11476 39142 11486 39194
rect 11486 39142 11532 39194
rect 11236 39140 11292 39142
rect 11316 39140 11372 39142
rect 11396 39140 11452 39142
rect 11476 39140 11532 39142
rect 9523 38650 9579 38652
rect 9603 38650 9659 38652
rect 9683 38650 9739 38652
rect 9763 38650 9819 38652
rect 9523 38598 9569 38650
rect 9569 38598 9579 38650
rect 9603 38598 9633 38650
rect 9633 38598 9645 38650
rect 9645 38598 9659 38650
rect 9683 38598 9697 38650
rect 9697 38598 9709 38650
rect 9709 38598 9739 38650
rect 9763 38598 9773 38650
rect 9773 38598 9819 38650
rect 9523 38596 9579 38598
rect 9603 38596 9659 38598
rect 9683 38596 9739 38598
rect 9763 38596 9819 38598
rect 7286 21664 7342 21720
rect 7102 19896 7158 19952
rect 7010 19760 7066 19816
rect 6096 13626 6152 13628
rect 6176 13626 6232 13628
rect 6256 13626 6312 13628
rect 6336 13626 6392 13628
rect 6096 13574 6142 13626
rect 6142 13574 6152 13626
rect 6176 13574 6206 13626
rect 6206 13574 6218 13626
rect 6218 13574 6232 13626
rect 6256 13574 6270 13626
rect 6270 13574 6282 13626
rect 6282 13574 6312 13626
rect 6336 13574 6346 13626
rect 6346 13574 6392 13626
rect 6096 13572 6152 13574
rect 6176 13572 6232 13574
rect 6256 13572 6312 13574
rect 6336 13572 6392 13574
rect 6096 12538 6152 12540
rect 6176 12538 6232 12540
rect 6256 12538 6312 12540
rect 6336 12538 6392 12540
rect 6096 12486 6142 12538
rect 6142 12486 6152 12538
rect 6176 12486 6206 12538
rect 6206 12486 6218 12538
rect 6218 12486 6232 12538
rect 6256 12486 6270 12538
rect 6270 12486 6282 12538
rect 6282 12486 6312 12538
rect 6336 12486 6346 12538
rect 6346 12486 6392 12538
rect 6096 12484 6152 12486
rect 6176 12484 6232 12486
rect 6256 12484 6312 12486
rect 6336 12484 6392 12486
rect 6096 11450 6152 11452
rect 6176 11450 6232 11452
rect 6256 11450 6312 11452
rect 6336 11450 6392 11452
rect 6096 11398 6142 11450
rect 6142 11398 6152 11450
rect 6176 11398 6206 11450
rect 6206 11398 6218 11450
rect 6218 11398 6232 11450
rect 6256 11398 6270 11450
rect 6270 11398 6282 11450
rect 6282 11398 6312 11450
rect 6336 11398 6346 11450
rect 6346 11398 6392 11450
rect 6096 11396 6152 11398
rect 6176 11396 6232 11398
rect 6256 11396 6312 11398
rect 6336 11396 6392 11398
rect 6096 10362 6152 10364
rect 6176 10362 6232 10364
rect 6256 10362 6312 10364
rect 6336 10362 6392 10364
rect 6096 10310 6142 10362
rect 6142 10310 6152 10362
rect 6176 10310 6206 10362
rect 6206 10310 6218 10362
rect 6218 10310 6232 10362
rect 6256 10310 6270 10362
rect 6270 10310 6282 10362
rect 6282 10310 6312 10362
rect 6336 10310 6346 10362
rect 6346 10310 6392 10362
rect 6096 10308 6152 10310
rect 6176 10308 6232 10310
rect 6256 10308 6312 10310
rect 6336 10308 6392 10310
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6336 9274 6392 9276
rect 6096 9222 6142 9274
rect 6142 9222 6152 9274
rect 6176 9222 6206 9274
rect 6206 9222 6218 9274
rect 6218 9222 6232 9274
rect 6256 9222 6270 9274
rect 6270 9222 6282 9274
rect 6282 9222 6312 9274
rect 6336 9222 6346 9274
rect 6346 9222 6392 9274
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 6336 9220 6392 9222
rect 7286 21528 7342 21584
rect 7809 31578 7865 31580
rect 7889 31578 7945 31580
rect 7969 31578 8025 31580
rect 8049 31578 8105 31580
rect 7809 31526 7855 31578
rect 7855 31526 7865 31578
rect 7889 31526 7919 31578
rect 7919 31526 7931 31578
rect 7931 31526 7945 31578
rect 7969 31526 7983 31578
rect 7983 31526 7995 31578
rect 7995 31526 8025 31578
rect 8049 31526 8059 31578
rect 8059 31526 8105 31578
rect 7809 31524 7865 31526
rect 7889 31524 7945 31526
rect 7969 31524 8025 31526
rect 8049 31524 8105 31526
rect 7809 30490 7865 30492
rect 7889 30490 7945 30492
rect 7969 30490 8025 30492
rect 8049 30490 8105 30492
rect 7809 30438 7855 30490
rect 7855 30438 7865 30490
rect 7889 30438 7919 30490
rect 7919 30438 7931 30490
rect 7931 30438 7945 30490
rect 7969 30438 7983 30490
rect 7983 30438 7995 30490
rect 7995 30438 8025 30490
rect 8049 30438 8059 30490
rect 8059 30438 8105 30490
rect 7809 30436 7865 30438
rect 7889 30436 7945 30438
rect 7969 30436 8025 30438
rect 8049 30436 8105 30438
rect 7809 29402 7865 29404
rect 7889 29402 7945 29404
rect 7969 29402 8025 29404
rect 8049 29402 8105 29404
rect 7809 29350 7855 29402
rect 7855 29350 7865 29402
rect 7889 29350 7919 29402
rect 7919 29350 7931 29402
rect 7931 29350 7945 29402
rect 7969 29350 7983 29402
rect 7983 29350 7995 29402
rect 7995 29350 8025 29402
rect 8049 29350 8059 29402
rect 8059 29350 8105 29402
rect 7809 29348 7865 29350
rect 7889 29348 7945 29350
rect 7969 29348 8025 29350
rect 8049 29348 8105 29350
rect 7809 28314 7865 28316
rect 7889 28314 7945 28316
rect 7969 28314 8025 28316
rect 8049 28314 8105 28316
rect 7809 28262 7855 28314
rect 7855 28262 7865 28314
rect 7889 28262 7919 28314
rect 7919 28262 7931 28314
rect 7931 28262 7945 28314
rect 7969 28262 7983 28314
rect 7983 28262 7995 28314
rect 7995 28262 8025 28314
rect 8049 28262 8059 28314
rect 8059 28262 8105 28314
rect 7809 28260 7865 28262
rect 7889 28260 7945 28262
rect 7969 28260 8025 28262
rect 8049 28260 8105 28262
rect 7809 27226 7865 27228
rect 7889 27226 7945 27228
rect 7969 27226 8025 27228
rect 8049 27226 8105 27228
rect 7809 27174 7855 27226
rect 7855 27174 7865 27226
rect 7889 27174 7919 27226
rect 7919 27174 7931 27226
rect 7931 27174 7945 27226
rect 7969 27174 7983 27226
rect 7983 27174 7995 27226
rect 7995 27174 8025 27226
rect 8049 27174 8059 27226
rect 8059 27174 8105 27226
rect 7809 27172 7865 27174
rect 7889 27172 7945 27174
rect 7969 27172 8025 27174
rect 8049 27172 8105 27174
rect 7286 20304 7342 20360
rect 7194 16088 7250 16144
rect 7102 12824 7158 12880
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6336 8186 6392 8188
rect 6096 8134 6142 8186
rect 6142 8134 6152 8186
rect 6176 8134 6206 8186
rect 6206 8134 6218 8186
rect 6218 8134 6232 8186
rect 6256 8134 6270 8186
rect 6270 8134 6282 8186
rect 6282 8134 6312 8186
rect 6336 8134 6346 8186
rect 6346 8134 6392 8186
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6336 8132 6392 8134
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6336 7098 6392 7100
rect 6096 7046 6142 7098
rect 6142 7046 6152 7098
rect 6176 7046 6206 7098
rect 6206 7046 6218 7098
rect 6218 7046 6232 7098
rect 6256 7046 6270 7098
rect 6270 7046 6282 7098
rect 6282 7046 6312 7098
rect 6336 7046 6346 7098
rect 6346 7046 6392 7098
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6336 7044 6392 7046
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6336 6010 6392 6012
rect 6096 5958 6142 6010
rect 6142 5958 6152 6010
rect 6176 5958 6206 6010
rect 6206 5958 6218 6010
rect 6218 5958 6232 6010
rect 6256 5958 6270 6010
rect 6270 5958 6282 6010
rect 6282 5958 6312 6010
rect 6336 5958 6346 6010
rect 6346 5958 6392 6010
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6336 5956 6392 5958
rect 7010 7948 7066 7984
rect 7010 7928 7012 7948
rect 7012 7928 7064 7948
rect 7064 7928 7066 7948
rect 4382 5466 4438 5468
rect 4462 5466 4518 5468
rect 4542 5466 4598 5468
rect 4622 5466 4678 5468
rect 4382 5414 4428 5466
rect 4428 5414 4438 5466
rect 4462 5414 4492 5466
rect 4492 5414 4504 5466
rect 4504 5414 4518 5466
rect 4542 5414 4556 5466
rect 4556 5414 4568 5466
rect 4568 5414 4598 5466
rect 4622 5414 4632 5466
rect 4632 5414 4678 5466
rect 4382 5412 4438 5414
rect 4462 5412 4518 5414
rect 4542 5412 4598 5414
rect 4622 5412 4678 5414
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6336 4922 6392 4924
rect 6096 4870 6142 4922
rect 6142 4870 6152 4922
rect 6176 4870 6206 4922
rect 6206 4870 6218 4922
rect 6218 4870 6232 4922
rect 6256 4870 6270 4922
rect 6270 4870 6282 4922
rect 6282 4870 6312 4922
rect 6336 4870 6346 4922
rect 6346 4870 6392 4922
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6336 4868 6392 4870
rect 4382 4378 4438 4380
rect 4462 4378 4518 4380
rect 4542 4378 4598 4380
rect 4622 4378 4678 4380
rect 4382 4326 4428 4378
rect 4428 4326 4438 4378
rect 4462 4326 4492 4378
rect 4492 4326 4504 4378
rect 4504 4326 4518 4378
rect 4542 4326 4556 4378
rect 4556 4326 4568 4378
rect 4568 4326 4598 4378
rect 4622 4326 4632 4378
rect 4632 4326 4678 4378
rect 4382 4324 4438 4326
rect 4462 4324 4518 4326
rect 4542 4324 4598 4326
rect 4622 4324 4678 4326
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6336 3834 6392 3836
rect 6096 3782 6142 3834
rect 6142 3782 6152 3834
rect 6176 3782 6206 3834
rect 6206 3782 6218 3834
rect 6218 3782 6232 3834
rect 6256 3782 6270 3834
rect 6270 3782 6282 3834
rect 6282 3782 6312 3834
rect 6336 3782 6346 3834
rect 6346 3782 6392 3834
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6336 3780 6392 3782
rect 4382 3290 4438 3292
rect 4462 3290 4518 3292
rect 4542 3290 4598 3292
rect 4622 3290 4678 3292
rect 4382 3238 4428 3290
rect 4428 3238 4438 3290
rect 4462 3238 4492 3290
rect 4492 3238 4504 3290
rect 4504 3238 4518 3290
rect 4542 3238 4556 3290
rect 4556 3238 4568 3290
rect 4568 3238 4598 3290
rect 4622 3238 4632 3290
rect 4632 3238 4678 3290
rect 4382 3236 4438 3238
rect 4462 3236 4518 3238
rect 4542 3236 4598 3238
rect 4622 3236 4678 3238
rect 7809 26138 7865 26140
rect 7889 26138 7945 26140
rect 7969 26138 8025 26140
rect 8049 26138 8105 26140
rect 7809 26086 7855 26138
rect 7855 26086 7865 26138
rect 7889 26086 7919 26138
rect 7919 26086 7931 26138
rect 7931 26086 7945 26138
rect 7969 26086 7983 26138
rect 7983 26086 7995 26138
rect 7995 26086 8025 26138
rect 8049 26086 8059 26138
rect 8059 26086 8105 26138
rect 7809 26084 7865 26086
rect 7889 26084 7945 26086
rect 7969 26084 8025 26086
rect 8049 26084 8105 26086
rect 8758 31184 8814 31240
rect 11236 38106 11292 38108
rect 11316 38106 11372 38108
rect 11396 38106 11452 38108
rect 11476 38106 11532 38108
rect 11236 38054 11282 38106
rect 11282 38054 11292 38106
rect 11316 38054 11346 38106
rect 11346 38054 11358 38106
rect 11358 38054 11372 38106
rect 11396 38054 11410 38106
rect 11410 38054 11422 38106
rect 11422 38054 11452 38106
rect 11476 38054 11486 38106
rect 11486 38054 11532 38106
rect 11236 38052 11292 38054
rect 11316 38052 11372 38054
rect 11396 38052 11452 38054
rect 11476 38052 11532 38054
rect 9523 37562 9579 37564
rect 9603 37562 9659 37564
rect 9683 37562 9739 37564
rect 9763 37562 9819 37564
rect 9523 37510 9569 37562
rect 9569 37510 9579 37562
rect 9603 37510 9633 37562
rect 9633 37510 9645 37562
rect 9645 37510 9659 37562
rect 9683 37510 9697 37562
rect 9697 37510 9709 37562
rect 9709 37510 9739 37562
rect 9763 37510 9773 37562
rect 9773 37510 9819 37562
rect 9523 37508 9579 37510
rect 9603 37508 9659 37510
rect 9683 37508 9739 37510
rect 9763 37508 9819 37510
rect 11236 37018 11292 37020
rect 11316 37018 11372 37020
rect 11396 37018 11452 37020
rect 11476 37018 11532 37020
rect 11236 36966 11282 37018
rect 11282 36966 11292 37018
rect 11316 36966 11346 37018
rect 11346 36966 11358 37018
rect 11358 36966 11372 37018
rect 11396 36966 11410 37018
rect 11410 36966 11422 37018
rect 11422 36966 11452 37018
rect 11476 36966 11486 37018
rect 11486 36966 11532 37018
rect 11236 36964 11292 36966
rect 11316 36964 11372 36966
rect 11396 36964 11452 36966
rect 11476 36964 11532 36966
rect 11794 38120 11850 38176
rect 12950 38650 13006 38652
rect 13030 38650 13086 38652
rect 13110 38650 13166 38652
rect 13190 38650 13246 38652
rect 12950 38598 12996 38650
rect 12996 38598 13006 38650
rect 13030 38598 13060 38650
rect 13060 38598 13072 38650
rect 13072 38598 13086 38650
rect 13110 38598 13124 38650
rect 13124 38598 13136 38650
rect 13136 38598 13166 38650
rect 13190 38598 13200 38650
rect 13200 38598 13246 38650
rect 12950 38596 13006 38598
rect 13030 38596 13086 38598
rect 13110 38596 13166 38598
rect 13190 38596 13246 38598
rect 13910 38936 13966 38992
rect 12950 37562 13006 37564
rect 13030 37562 13086 37564
rect 13110 37562 13166 37564
rect 13190 37562 13246 37564
rect 12950 37510 12996 37562
rect 12996 37510 13006 37562
rect 13030 37510 13060 37562
rect 13060 37510 13072 37562
rect 13072 37510 13086 37562
rect 13110 37510 13124 37562
rect 13124 37510 13136 37562
rect 13136 37510 13166 37562
rect 13190 37510 13200 37562
rect 13200 37510 13246 37562
rect 12950 37508 13006 37510
rect 13030 37508 13086 37510
rect 13110 37508 13166 37510
rect 13190 37508 13246 37510
rect 12806 37204 12808 37224
rect 12808 37204 12860 37224
rect 12860 37204 12862 37224
rect 11334 36644 11390 36680
rect 11334 36624 11336 36644
rect 11336 36624 11388 36644
rect 11388 36624 11390 36644
rect 9523 36474 9579 36476
rect 9603 36474 9659 36476
rect 9683 36474 9739 36476
rect 9763 36474 9819 36476
rect 9523 36422 9569 36474
rect 9569 36422 9579 36474
rect 9603 36422 9633 36474
rect 9633 36422 9645 36474
rect 9645 36422 9659 36474
rect 9683 36422 9697 36474
rect 9697 36422 9709 36474
rect 9709 36422 9739 36474
rect 9763 36422 9773 36474
rect 9773 36422 9819 36474
rect 9523 36420 9579 36422
rect 9603 36420 9659 36422
rect 9683 36420 9739 36422
rect 9763 36420 9819 36422
rect 9523 35386 9579 35388
rect 9603 35386 9659 35388
rect 9683 35386 9739 35388
rect 9763 35386 9819 35388
rect 9523 35334 9569 35386
rect 9569 35334 9579 35386
rect 9603 35334 9633 35386
rect 9633 35334 9645 35386
rect 9645 35334 9659 35386
rect 9683 35334 9697 35386
rect 9697 35334 9709 35386
rect 9709 35334 9739 35386
rect 9763 35334 9773 35386
rect 9773 35334 9819 35386
rect 9523 35332 9579 35334
rect 9603 35332 9659 35334
rect 9683 35332 9739 35334
rect 9763 35332 9819 35334
rect 11236 35930 11292 35932
rect 11316 35930 11372 35932
rect 11396 35930 11452 35932
rect 11476 35930 11532 35932
rect 11236 35878 11282 35930
rect 11282 35878 11292 35930
rect 11316 35878 11346 35930
rect 11346 35878 11358 35930
rect 11358 35878 11372 35930
rect 11396 35878 11410 35930
rect 11410 35878 11422 35930
rect 11422 35878 11452 35930
rect 11476 35878 11486 35930
rect 11486 35878 11532 35930
rect 11236 35876 11292 35878
rect 11316 35876 11372 35878
rect 11396 35876 11452 35878
rect 11476 35876 11532 35878
rect 10966 34992 11022 35048
rect 9523 34298 9579 34300
rect 9603 34298 9659 34300
rect 9683 34298 9739 34300
rect 9763 34298 9819 34300
rect 9523 34246 9569 34298
rect 9569 34246 9579 34298
rect 9603 34246 9633 34298
rect 9633 34246 9645 34298
rect 9645 34246 9659 34298
rect 9683 34246 9697 34298
rect 9697 34246 9709 34298
rect 9709 34246 9739 34298
rect 9763 34246 9773 34298
rect 9773 34246 9819 34298
rect 9523 34244 9579 34246
rect 9603 34244 9659 34246
rect 9683 34244 9739 34246
rect 9763 34244 9819 34246
rect 9523 33210 9579 33212
rect 9603 33210 9659 33212
rect 9683 33210 9739 33212
rect 9763 33210 9819 33212
rect 9523 33158 9569 33210
rect 9569 33158 9579 33210
rect 9603 33158 9633 33210
rect 9633 33158 9645 33210
rect 9645 33158 9659 33210
rect 9683 33158 9697 33210
rect 9697 33158 9709 33210
rect 9709 33158 9739 33210
rect 9763 33158 9773 33210
rect 9773 33158 9819 33210
rect 9523 33156 9579 33158
rect 9603 33156 9659 33158
rect 9683 33156 9739 33158
rect 9763 33156 9819 33158
rect 9523 32122 9579 32124
rect 9603 32122 9659 32124
rect 9683 32122 9739 32124
rect 9763 32122 9819 32124
rect 9523 32070 9569 32122
rect 9569 32070 9579 32122
rect 9603 32070 9633 32122
rect 9633 32070 9645 32122
rect 9645 32070 9659 32122
rect 9683 32070 9697 32122
rect 9697 32070 9709 32122
rect 9709 32070 9739 32122
rect 9763 32070 9773 32122
rect 9773 32070 9819 32122
rect 9523 32068 9579 32070
rect 9603 32068 9659 32070
rect 9683 32068 9739 32070
rect 9763 32068 9819 32070
rect 7809 25050 7865 25052
rect 7889 25050 7945 25052
rect 7969 25050 8025 25052
rect 8049 25050 8105 25052
rect 7809 24998 7855 25050
rect 7855 24998 7865 25050
rect 7889 24998 7919 25050
rect 7919 24998 7931 25050
rect 7931 24998 7945 25050
rect 7969 24998 7983 25050
rect 7983 24998 7995 25050
rect 7995 24998 8025 25050
rect 8049 24998 8059 25050
rect 8059 24998 8105 25050
rect 7809 24996 7865 24998
rect 7889 24996 7945 24998
rect 7969 24996 8025 24998
rect 8049 24996 8105 24998
rect 7809 23962 7865 23964
rect 7889 23962 7945 23964
rect 7969 23962 8025 23964
rect 8049 23962 8105 23964
rect 7809 23910 7855 23962
rect 7855 23910 7865 23962
rect 7889 23910 7919 23962
rect 7919 23910 7931 23962
rect 7931 23910 7945 23962
rect 7969 23910 7983 23962
rect 7983 23910 7995 23962
rect 7995 23910 8025 23962
rect 8049 23910 8059 23962
rect 8059 23910 8105 23962
rect 7809 23908 7865 23910
rect 7889 23908 7945 23910
rect 7969 23908 8025 23910
rect 8049 23908 8105 23910
rect 7809 22874 7865 22876
rect 7889 22874 7945 22876
rect 7969 22874 8025 22876
rect 8049 22874 8105 22876
rect 7809 22822 7855 22874
rect 7855 22822 7865 22874
rect 7889 22822 7919 22874
rect 7919 22822 7931 22874
rect 7931 22822 7945 22874
rect 7969 22822 7983 22874
rect 7983 22822 7995 22874
rect 7995 22822 8025 22874
rect 8049 22822 8059 22874
rect 8059 22822 8105 22874
rect 7809 22820 7865 22822
rect 7889 22820 7945 22822
rect 7969 22820 8025 22822
rect 8049 22820 8105 22822
rect 7809 21786 7865 21788
rect 7889 21786 7945 21788
rect 7969 21786 8025 21788
rect 8049 21786 8105 21788
rect 7809 21734 7855 21786
rect 7855 21734 7865 21786
rect 7889 21734 7919 21786
rect 7919 21734 7931 21786
rect 7931 21734 7945 21786
rect 7969 21734 7983 21786
rect 7983 21734 7995 21786
rect 7995 21734 8025 21786
rect 8049 21734 8059 21786
rect 8059 21734 8105 21786
rect 7809 21732 7865 21734
rect 7889 21732 7945 21734
rect 7969 21732 8025 21734
rect 8049 21732 8105 21734
rect 7809 20698 7865 20700
rect 7889 20698 7945 20700
rect 7969 20698 8025 20700
rect 8049 20698 8105 20700
rect 7809 20646 7855 20698
rect 7855 20646 7865 20698
rect 7889 20646 7919 20698
rect 7919 20646 7931 20698
rect 7931 20646 7945 20698
rect 7969 20646 7983 20698
rect 7983 20646 7995 20698
rect 7995 20646 8025 20698
rect 8049 20646 8059 20698
rect 8059 20646 8105 20698
rect 7809 20644 7865 20646
rect 7889 20644 7945 20646
rect 7969 20644 8025 20646
rect 8049 20644 8105 20646
rect 8206 20576 8262 20632
rect 8206 19760 8262 19816
rect 7809 19610 7865 19612
rect 7889 19610 7945 19612
rect 7969 19610 8025 19612
rect 8049 19610 8105 19612
rect 7809 19558 7855 19610
rect 7855 19558 7865 19610
rect 7889 19558 7919 19610
rect 7919 19558 7931 19610
rect 7931 19558 7945 19610
rect 7969 19558 7983 19610
rect 7983 19558 7995 19610
rect 7995 19558 8025 19610
rect 8049 19558 8059 19610
rect 8059 19558 8105 19610
rect 7809 19556 7865 19558
rect 7889 19556 7945 19558
rect 7969 19556 8025 19558
rect 8049 19556 8105 19558
rect 7809 18522 7865 18524
rect 7889 18522 7945 18524
rect 7969 18522 8025 18524
rect 8049 18522 8105 18524
rect 7809 18470 7855 18522
rect 7855 18470 7865 18522
rect 7889 18470 7919 18522
rect 7919 18470 7931 18522
rect 7931 18470 7945 18522
rect 7969 18470 7983 18522
rect 7983 18470 7995 18522
rect 7995 18470 8025 18522
rect 8049 18470 8059 18522
rect 8059 18470 8105 18522
rect 7809 18468 7865 18470
rect 7889 18468 7945 18470
rect 7969 18468 8025 18470
rect 8049 18468 8105 18470
rect 7809 17434 7865 17436
rect 7889 17434 7945 17436
rect 7969 17434 8025 17436
rect 8049 17434 8105 17436
rect 7809 17382 7855 17434
rect 7855 17382 7865 17434
rect 7889 17382 7919 17434
rect 7919 17382 7931 17434
rect 7931 17382 7945 17434
rect 7969 17382 7983 17434
rect 7983 17382 7995 17434
rect 7995 17382 8025 17434
rect 8049 17382 8059 17434
rect 8059 17382 8105 17434
rect 7809 17380 7865 17382
rect 7889 17380 7945 17382
rect 7969 17380 8025 17382
rect 8049 17380 8105 17382
rect 8206 17312 8262 17368
rect 8942 29008 8998 29064
rect 9218 29008 9274 29064
rect 8758 26288 8814 26344
rect 8482 23196 8484 23216
rect 8484 23196 8536 23216
rect 8536 23196 8538 23216
rect 8482 23160 8538 23196
rect 8482 23044 8538 23080
rect 8482 23024 8484 23044
rect 8484 23024 8536 23044
rect 8536 23024 8538 23044
rect 8482 21800 8538 21856
rect 8850 21800 8906 21856
rect 7809 16346 7865 16348
rect 7889 16346 7945 16348
rect 7969 16346 8025 16348
rect 8049 16346 8105 16348
rect 7809 16294 7855 16346
rect 7855 16294 7865 16346
rect 7889 16294 7919 16346
rect 7919 16294 7931 16346
rect 7931 16294 7945 16346
rect 7969 16294 7983 16346
rect 7983 16294 7995 16346
rect 7995 16294 8025 16346
rect 8049 16294 8059 16346
rect 8059 16294 8105 16346
rect 7809 16292 7865 16294
rect 7889 16292 7945 16294
rect 7969 16292 8025 16294
rect 8049 16292 8105 16294
rect 7809 15258 7865 15260
rect 7889 15258 7945 15260
rect 7969 15258 8025 15260
rect 8049 15258 8105 15260
rect 7809 15206 7855 15258
rect 7855 15206 7865 15258
rect 7889 15206 7919 15258
rect 7919 15206 7931 15258
rect 7931 15206 7945 15258
rect 7969 15206 7983 15258
rect 7983 15206 7995 15258
rect 7995 15206 8025 15258
rect 8049 15206 8059 15258
rect 8059 15206 8105 15258
rect 7809 15204 7865 15206
rect 7889 15204 7945 15206
rect 7969 15204 8025 15206
rect 8049 15204 8105 15206
rect 8206 14320 8262 14376
rect 7809 14170 7865 14172
rect 7889 14170 7945 14172
rect 7969 14170 8025 14172
rect 8049 14170 8105 14172
rect 7809 14118 7855 14170
rect 7855 14118 7865 14170
rect 7889 14118 7919 14170
rect 7919 14118 7931 14170
rect 7931 14118 7945 14170
rect 7969 14118 7983 14170
rect 7983 14118 7995 14170
rect 7995 14118 8025 14170
rect 8049 14118 8059 14170
rect 8059 14118 8105 14170
rect 7809 14116 7865 14118
rect 7889 14116 7945 14118
rect 7969 14116 8025 14118
rect 8049 14116 8105 14118
rect 8298 13912 8354 13968
rect 8298 13640 8354 13696
rect 7809 13082 7865 13084
rect 7889 13082 7945 13084
rect 7969 13082 8025 13084
rect 8049 13082 8105 13084
rect 7809 13030 7855 13082
rect 7855 13030 7865 13082
rect 7889 13030 7919 13082
rect 7919 13030 7931 13082
rect 7931 13030 7945 13082
rect 7969 13030 7983 13082
rect 7983 13030 7995 13082
rect 7995 13030 8025 13082
rect 8049 13030 8059 13082
rect 8059 13030 8105 13082
rect 7809 13028 7865 13030
rect 7889 13028 7945 13030
rect 7969 13028 8025 13030
rect 8049 13028 8105 13030
rect 7654 12724 7656 12744
rect 7656 12724 7708 12744
rect 7708 12724 7710 12744
rect 7654 12688 7710 12724
rect 7809 11994 7865 11996
rect 7889 11994 7945 11996
rect 7969 11994 8025 11996
rect 8049 11994 8105 11996
rect 7809 11942 7855 11994
rect 7855 11942 7865 11994
rect 7889 11942 7919 11994
rect 7919 11942 7931 11994
rect 7931 11942 7945 11994
rect 7969 11942 7983 11994
rect 7983 11942 7995 11994
rect 7995 11942 8025 11994
rect 8049 11942 8059 11994
rect 8059 11942 8105 11994
rect 7809 11940 7865 11942
rect 7889 11940 7945 11942
rect 7969 11940 8025 11942
rect 8049 11940 8105 11942
rect 7809 10906 7865 10908
rect 7889 10906 7945 10908
rect 7969 10906 8025 10908
rect 8049 10906 8105 10908
rect 7809 10854 7855 10906
rect 7855 10854 7865 10906
rect 7889 10854 7919 10906
rect 7919 10854 7931 10906
rect 7931 10854 7945 10906
rect 7969 10854 7983 10906
rect 7983 10854 7995 10906
rect 7995 10854 8025 10906
rect 8049 10854 8059 10906
rect 8059 10854 8105 10906
rect 7809 10852 7865 10854
rect 7889 10852 7945 10854
rect 7969 10852 8025 10854
rect 8049 10852 8105 10854
rect 9126 19624 9182 19680
rect 8482 14184 8538 14240
rect 7809 9818 7865 9820
rect 7889 9818 7945 9820
rect 7969 9818 8025 9820
rect 8049 9818 8105 9820
rect 7809 9766 7855 9818
rect 7855 9766 7865 9818
rect 7889 9766 7919 9818
rect 7919 9766 7931 9818
rect 7931 9766 7945 9818
rect 7969 9766 7983 9818
rect 7983 9766 7995 9818
rect 7995 9766 8025 9818
rect 8049 9766 8059 9818
rect 8059 9766 8105 9818
rect 7809 9764 7865 9766
rect 7889 9764 7945 9766
rect 7969 9764 8025 9766
rect 8049 9764 8105 9766
rect 7809 8730 7865 8732
rect 7889 8730 7945 8732
rect 7969 8730 8025 8732
rect 8049 8730 8105 8732
rect 7809 8678 7855 8730
rect 7855 8678 7865 8730
rect 7889 8678 7919 8730
rect 7919 8678 7931 8730
rect 7931 8678 7945 8730
rect 7969 8678 7983 8730
rect 7983 8678 7995 8730
rect 7995 8678 8025 8730
rect 8049 8678 8059 8730
rect 8059 8678 8105 8730
rect 7809 8676 7865 8678
rect 7889 8676 7945 8678
rect 7969 8676 8025 8678
rect 8049 8676 8105 8678
rect 7809 7642 7865 7644
rect 7889 7642 7945 7644
rect 7969 7642 8025 7644
rect 8049 7642 8105 7644
rect 7809 7590 7855 7642
rect 7855 7590 7865 7642
rect 7889 7590 7919 7642
rect 7919 7590 7931 7642
rect 7931 7590 7945 7642
rect 7969 7590 7983 7642
rect 7983 7590 7995 7642
rect 7995 7590 8025 7642
rect 8049 7590 8059 7642
rect 8059 7590 8105 7642
rect 7809 7588 7865 7590
rect 7889 7588 7945 7590
rect 7969 7588 8025 7590
rect 8049 7588 8105 7590
rect 7809 6554 7865 6556
rect 7889 6554 7945 6556
rect 7969 6554 8025 6556
rect 8049 6554 8105 6556
rect 7809 6502 7855 6554
rect 7855 6502 7865 6554
rect 7889 6502 7919 6554
rect 7919 6502 7931 6554
rect 7931 6502 7945 6554
rect 7969 6502 7983 6554
rect 7983 6502 7995 6554
rect 7995 6502 8025 6554
rect 8049 6502 8059 6554
rect 8059 6502 8105 6554
rect 7809 6500 7865 6502
rect 7889 6500 7945 6502
rect 7969 6500 8025 6502
rect 8049 6500 8105 6502
rect 8298 6332 8300 6352
rect 8300 6332 8352 6352
rect 8352 6332 8354 6352
rect 8298 6296 8354 6332
rect 8206 5652 8208 5672
rect 8208 5652 8260 5672
rect 8260 5652 8262 5672
rect 8206 5616 8262 5652
rect 7809 5466 7865 5468
rect 7889 5466 7945 5468
rect 7969 5466 8025 5468
rect 8049 5466 8105 5468
rect 7809 5414 7855 5466
rect 7855 5414 7865 5466
rect 7889 5414 7919 5466
rect 7919 5414 7931 5466
rect 7931 5414 7945 5466
rect 7969 5414 7983 5466
rect 7983 5414 7995 5466
rect 7995 5414 8025 5466
rect 8049 5414 8059 5466
rect 8059 5414 8105 5466
rect 7809 5412 7865 5414
rect 7889 5412 7945 5414
rect 7969 5412 8025 5414
rect 8049 5412 8105 5414
rect 7809 4378 7865 4380
rect 7889 4378 7945 4380
rect 7969 4378 8025 4380
rect 8049 4378 8105 4380
rect 7809 4326 7855 4378
rect 7855 4326 7865 4378
rect 7889 4326 7919 4378
rect 7919 4326 7931 4378
rect 7931 4326 7945 4378
rect 7969 4326 7983 4378
rect 7983 4326 7995 4378
rect 7995 4326 8025 4378
rect 8049 4326 8059 4378
rect 8059 4326 8105 4378
rect 7809 4324 7865 4326
rect 7889 4324 7945 4326
rect 7969 4324 8025 4326
rect 8049 4324 8105 4326
rect 7809 3290 7865 3292
rect 7889 3290 7945 3292
rect 7969 3290 8025 3292
rect 8049 3290 8105 3292
rect 7809 3238 7855 3290
rect 7855 3238 7865 3290
rect 7889 3238 7919 3290
rect 7919 3238 7931 3290
rect 7931 3238 7945 3290
rect 7969 3238 7983 3290
rect 7983 3238 7995 3290
rect 7995 3238 8025 3290
rect 8049 3238 8059 3290
rect 8059 3238 8105 3290
rect 7809 3236 7865 3238
rect 7889 3236 7945 3238
rect 7969 3236 8025 3238
rect 8049 3236 8105 3238
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6336 2746 6392 2748
rect 6096 2694 6142 2746
rect 6142 2694 6152 2746
rect 6176 2694 6206 2746
rect 6206 2694 6218 2746
rect 6218 2694 6232 2746
rect 6256 2694 6270 2746
rect 6270 2694 6282 2746
rect 6282 2694 6312 2746
rect 6336 2694 6346 2746
rect 6346 2694 6392 2746
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 6336 2692 6392 2694
rect 5814 2624 5870 2680
rect 6642 2624 6698 2680
rect 4382 2202 4438 2204
rect 4462 2202 4518 2204
rect 4542 2202 4598 2204
rect 4622 2202 4678 2204
rect 4382 2150 4428 2202
rect 4428 2150 4438 2202
rect 4462 2150 4492 2202
rect 4492 2150 4504 2202
rect 4504 2150 4518 2202
rect 4542 2150 4556 2202
rect 4556 2150 4568 2202
rect 4568 2150 4598 2202
rect 4622 2150 4632 2202
rect 4632 2150 4678 2202
rect 4382 2148 4438 2150
rect 4462 2148 4518 2150
rect 4542 2148 4598 2150
rect 4622 2148 4678 2150
rect 7654 2624 7710 2680
rect 7809 2202 7865 2204
rect 7889 2202 7945 2204
rect 7969 2202 8025 2204
rect 8049 2202 8105 2204
rect 7809 2150 7855 2202
rect 7855 2150 7865 2202
rect 7889 2150 7919 2202
rect 7919 2150 7931 2202
rect 7931 2150 7945 2202
rect 7969 2150 7983 2202
rect 7983 2150 7995 2202
rect 7995 2150 8025 2202
rect 8049 2150 8059 2202
rect 8059 2150 8105 2202
rect 7809 2148 7865 2150
rect 7889 2148 7945 2150
rect 7969 2148 8025 2150
rect 8049 2148 8105 2150
rect 2669 1658 2725 1660
rect 2749 1658 2805 1660
rect 2829 1658 2885 1660
rect 2909 1658 2965 1660
rect 2669 1606 2715 1658
rect 2715 1606 2725 1658
rect 2749 1606 2779 1658
rect 2779 1606 2791 1658
rect 2791 1606 2805 1658
rect 2829 1606 2843 1658
rect 2843 1606 2855 1658
rect 2855 1606 2885 1658
rect 2909 1606 2919 1658
rect 2919 1606 2965 1658
rect 2669 1604 2725 1606
rect 2749 1604 2805 1606
rect 2829 1604 2885 1606
rect 2909 1604 2965 1606
rect 6096 1658 6152 1660
rect 6176 1658 6232 1660
rect 6256 1658 6312 1660
rect 6336 1658 6392 1660
rect 6096 1606 6142 1658
rect 6142 1606 6152 1658
rect 6176 1606 6206 1658
rect 6206 1606 6218 1658
rect 6218 1606 6232 1658
rect 6256 1606 6270 1658
rect 6270 1606 6282 1658
rect 6282 1606 6312 1658
rect 6336 1606 6346 1658
rect 6346 1606 6392 1658
rect 6096 1604 6152 1606
rect 6176 1604 6232 1606
rect 6256 1604 6312 1606
rect 6336 1604 6392 1606
rect 4382 1114 4438 1116
rect 4462 1114 4518 1116
rect 4542 1114 4598 1116
rect 4622 1114 4678 1116
rect 4382 1062 4428 1114
rect 4428 1062 4438 1114
rect 4462 1062 4492 1114
rect 4492 1062 4504 1114
rect 4504 1062 4518 1114
rect 4542 1062 4556 1114
rect 4556 1062 4568 1114
rect 4568 1062 4598 1114
rect 4622 1062 4632 1114
rect 4632 1062 4678 1114
rect 4382 1060 4438 1062
rect 4462 1060 4518 1062
rect 4542 1060 4598 1062
rect 4622 1060 4678 1062
rect 7809 1114 7865 1116
rect 7889 1114 7945 1116
rect 7969 1114 8025 1116
rect 8049 1114 8105 1116
rect 7809 1062 7855 1114
rect 7855 1062 7865 1114
rect 7889 1062 7919 1114
rect 7919 1062 7931 1114
rect 7931 1062 7945 1114
rect 7969 1062 7983 1114
rect 7983 1062 7995 1114
rect 7995 1062 8025 1114
rect 8049 1062 8059 1114
rect 8059 1062 8105 1114
rect 7809 1060 7865 1062
rect 7889 1060 7945 1062
rect 7969 1060 8025 1062
rect 8049 1060 8105 1062
rect 9523 31034 9579 31036
rect 9603 31034 9659 31036
rect 9683 31034 9739 31036
rect 9763 31034 9819 31036
rect 9523 30982 9569 31034
rect 9569 30982 9579 31034
rect 9603 30982 9633 31034
rect 9633 30982 9645 31034
rect 9645 30982 9659 31034
rect 9683 30982 9697 31034
rect 9697 30982 9709 31034
rect 9709 30982 9739 31034
rect 9763 30982 9773 31034
rect 9773 30982 9819 31034
rect 9523 30980 9579 30982
rect 9603 30980 9659 30982
rect 9683 30980 9739 30982
rect 9763 30980 9819 30982
rect 11236 34842 11292 34844
rect 11316 34842 11372 34844
rect 11396 34842 11452 34844
rect 11476 34842 11532 34844
rect 11236 34790 11282 34842
rect 11282 34790 11292 34842
rect 11316 34790 11346 34842
rect 11346 34790 11358 34842
rect 11358 34790 11372 34842
rect 11396 34790 11410 34842
rect 11410 34790 11422 34842
rect 11422 34790 11452 34842
rect 11476 34790 11486 34842
rect 11486 34790 11532 34842
rect 11236 34788 11292 34790
rect 11316 34788 11372 34790
rect 11396 34788 11452 34790
rect 11476 34788 11532 34790
rect 12806 37168 12862 37204
rect 12990 36624 13046 36680
rect 12950 36474 13006 36476
rect 13030 36474 13086 36476
rect 13110 36474 13166 36476
rect 13190 36474 13246 36476
rect 12950 36422 12996 36474
rect 12996 36422 13006 36474
rect 13030 36422 13060 36474
rect 13060 36422 13072 36474
rect 13072 36422 13086 36474
rect 13110 36422 13124 36474
rect 13124 36422 13136 36474
rect 13136 36422 13166 36474
rect 13190 36422 13200 36474
rect 13200 36422 13246 36474
rect 12950 36420 13006 36422
rect 13030 36420 13086 36422
rect 13110 36420 13166 36422
rect 13190 36420 13246 36422
rect 11236 33754 11292 33756
rect 11316 33754 11372 33756
rect 11396 33754 11452 33756
rect 11476 33754 11532 33756
rect 11236 33702 11282 33754
rect 11282 33702 11292 33754
rect 11316 33702 11346 33754
rect 11346 33702 11358 33754
rect 11358 33702 11372 33754
rect 11396 33702 11410 33754
rect 11410 33702 11422 33754
rect 11422 33702 11452 33754
rect 11476 33702 11486 33754
rect 11486 33702 11532 33754
rect 11236 33700 11292 33702
rect 11316 33700 11372 33702
rect 11396 33700 11452 33702
rect 11476 33700 11532 33702
rect 11426 33088 11482 33144
rect 9523 29946 9579 29948
rect 9603 29946 9659 29948
rect 9683 29946 9739 29948
rect 9763 29946 9819 29948
rect 9523 29894 9569 29946
rect 9569 29894 9579 29946
rect 9603 29894 9633 29946
rect 9633 29894 9645 29946
rect 9645 29894 9659 29946
rect 9683 29894 9697 29946
rect 9697 29894 9709 29946
rect 9709 29894 9739 29946
rect 9763 29894 9773 29946
rect 9773 29894 9819 29946
rect 9523 29892 9579 29894
rect 9603 29892 9659 29894
rect 9683 29892 9739 29894
rect 9763 29892 9819 29894
rect 9523 28858 9579 28860
rect 9603 28858 9659 28860
rect 9683 28858 9739 28860
rect 9763 28858 9819 28860
rect 9523 28806 9569 28858
rect 9569 28806 9579 28858
rect 9603 28806 9633 28858
rect 9633 28806 9645 28858
rect 9645 28806 9659 28858
rect 9683 28806 9697 28858
rect 9697 28806 9709 28858
rect 9709 28806 9739 28858
rect 9763 28806 9773 28858
rect 9773 28806 9819 28858
rect 9523 28804 9579 28806
rect 9603 28804 9659 28806
rect 9683 28804 9739 28806
rect 9763 28804 9819 28806
rect 9523 27770 9579 27772
rect 9603 27770 9659 27772
rect 9683 27770 9739 27772
rect 9763 27770 9819 27772
rect 9523 27718 9569 27770
rect 9569 27718 9579 27770
rect 9603 27718 9633 27770
rect 9633 27718 9645 27770
rect 9645 27718 9659 27770
rect 9683 27718 9697 27770
rect 9697 27718 9709 27770
rect 9709 27718 9739 27770
rect 9763 27718 9773 27770
rect 9773 27718 9819 27770
rect 9523 27716 9579 27718
rect 9603 27716 9659 27718
rect 9683 27716 9739 27718
rect 9763 27716 9819 27718
rect 9523 26682 9579 26684
rect 9603 26682 9659 26684
rect 9683 26682 9739 26684
rect 9763 26682 9819 26684
rect 9523 26630 9569 26682
rect 9569 26630 9579 26682
rect 9603 26630 9633 26682
rect 9633 26630 9645 26682
rect 9645 26630 9659 26682
rect 9683 26630 9697 26682
rect 9697 26630 9709 26682
rect 9709 26630 9739 26682
rect 9763 26630 9773 26682
rect 9773 26630 9819 26682
rect 9523 26628 9579 26630
rect 9603 26628 9659 26630
rect 9683 26628 9739 26630
rect 9763 26628 9819 26630
rect 9954 25880 10010 25936
rect 9523 25594 9579 25596
rect 9603 25594 9659 25596
rect 9683 25594 9739 25596
rect 9763 25594 9819 25596
rect 9523 25542 9569 25594
rect 9569 25542 9579 25594
rect 9603 25542 9633 25594
rect 9633 25542 9645 25594
rect 9645 25542 9659 25594
rect 9683 25542 9697 25594
rect 9697 25542 9709 25594
rect 9709 25542 9739 25594
rect 9763 25542 9773 25594
rect 9773 25542 9819 25594
rect 9523 25540 9579 25542
rect 9603 25540 9659 25542
rect 9683 25540 9739 25542
rect 9763 25540 9819 25542
rect 9770 24792 9826 24848
rect 9862 24656 9918 24712
rect 9523 24506 9579 24508
rect 9603 24506 9659 24508
rect 9683 24506 9739 24508
rect 9763 24506 9819 24508
rect 9523 24454 9569 24506
rect 9569 24454 9579 24506
rect 9603 24454 9633 24506
rect 9633 24454 9645 24506
rect 9645 24454 9659 24506
rect 9683 24454 9697 24506
rect 9697 24454 9709 24506
rect 9709 24454 9739 24506
rect 9763 24454 9773 24506
rect 9773 24454 9819 24506
rect 9523 24452 9579 24454
rect 9603 24452 9659 24454
rect 9683 24452 9739 24454
rect 9763 24452 9819 24454
rect 9523 23418 9579 23420
rect 9603 23418 9659 23420
rect 9683 23418 9739 23420
rect 9763 23418 9819 23420
rect 9523 23366 9569 23418
rect 9569 23366 9579 23418
rect 9603 23366 9633 23418
rect 9633 23366 9645 23418
rect 9645 23366 9659 23418
rect 9683 23366 9697 23418
rect 9697 23366 9709 23418
rect 9709 23366 9739 23418
rect 9763 23366 9773 23418
rect 9773 23366 9819 23418
rect 9523 23364 9579 23366
rect 9603 23364 9659 23366
rect 9683 23364 9739 23366
rect 9763 23364 9819 23366
rect 9523 22330 9579 22332
rect 9603 22330 9659 22332
rect 9683 22330 9739 22332
rect 9763 22330 9819 22332
rect 9523 22278 9569 22330
rect 9569 22278 9579 22330
rect 9603 22278 9633 22330
rect 9633 22278 9645 22330
rect 9645 22278 9659 22330
rect 9683 22278 9697 22330
rect 9697 22278 9709 22330
rect 9709 22278 9739 22330
rect 9763 22278 9773 22330
rect 9773 22278 9819 22330
rect 9523 22276 9579 22278
rect 9603 22276 9659 22278
rect 9683 22276 9739 22278
rect 9763 22276 9819 22278
rect 10322 31320 10378 31376
rect 11058 32408 11114 32464
rect 11236 32666 11292 32668
rect 11316 32666 11372 32668
rect 11396 32666 11452 32668
rect 11476 32666 11532 32668
rect 11236 32614 11282 32666
rect 11282 32614 11292 32666
rect 11316 32614 11346 32666
rect 11346 32614 11358 32666
rect 11358 32614 11372 32666
rect 11396 32614 11410 32666
rect 11410 32614 11422 32666
rect 11422 32614 11452 32666
rect 11476 32614 11486 32666
rect 11486 32614 11532 32666
rect 11236 32612 11292 32614
rect 11316 32612 11372 32614
rect 11396 32612 11452 32614
rect 11476 32612 11532 32614
rect 10966 31864 11022 31920
rect 11236 31578 11292 31580
rect 11316 31578 11372 31580
rect 11396 31578 11452 31580
rect 11476 31578 11532 31580
rect 11236 31526 11282 31578
rect 11282 31526 11292 31578
rect 11316 31526 11346 31578
rect 11346 31526 11358 31578
rect 11358 31526 11372 31578
rect 11396 31526 11410 31578
rect 11410 31526 11422 31578
rect 11422 31526 11452 31578
rect 11476 31526 11486 31578
rect 11486 31526 11532 31578
rect 11236 31524 11292 31526
rect 11316 31524 11372 31526
rect 11396 31524 11452 31526
rect 11476 31524 11532 31526
rect 11794 32272 11850 32328
rect 11518 31048 11574 31104
rect 11236 30490 11292 30492
rect 11316 30490 11372 30492
rect 11396 30490 11452 30492
rect 11476 30490 11532 30492
rect 11236 30438 11282 30490
rect 11282 30438 11292 30490
rect 11316 30438 11346 30490
rect 11346 30438 11358 30490
rect 11358 30438 11372 30490
rect 11396 30438 11410 30490
rect 11410 30438 11422 30490
rect 11422 30438 11452 30490
rect 11476 30438 11486 30490
rect 11486 30438 11532 30490
rect 11236 30436 11292 30438
rect 11316 30436 11372 30438
rect 11396 30436 11452 30438
rect 11476 30436 11532 30438
rect 10414 24792 10470 24848
rect 9494 21392 9550 21448
rect 9954 21972 9956 21992
rect 9956 21972 10008 21992
rect 10008 21972 10010 21992
rect 9954 21936 10010 21972
rect 9862 21392 9918 21448
rect 9523 21242 9579 21244
rect 9603 21242 9659 21244
rect 9683 21242 9739 21244
rect 9763 21242 9819 21244
rect 9523 21190 9569 21242
rect 9569 21190 9579 21242
rect 9603 21190 9633 21242
rect 9633 21190 9645 21242
rect 9645 21190 9659 21242
rect 9683 21190 9697 21242
rect 9697 21190 9709 21242
rect 9709 21190 9739 21242
rect 9763 21190 9773 21242
rect 9773 21190 9819 21242
rect 9523 21188 9579 21190
rect 9603 21188 9659 21190
rect 9683 21188 9739 21190
rect 9763 21188 9819 21190
rect 9126 14864 9182 14920
rect 8942 14184 8998 14240
rect 9034 13776 9090 13832
rect 8758 11736 8814 11792
rect 9523 20154 9579 20156
rect 9603 20154 9659 20156
rect 9683 20154 9739 20156
rect 9763 20154 9819 20156
rect 9523 20102 9569 20154
rect 9569 20102 9579 20154
rect 9603 20102 9633 20154
rect 9633 20102 9645 20154
rect 9645 20102 9659 20154
rect 9683 20102 9697 20154
rect 9697 20102 9709 20154
rect 9709 20102 9739 20154
rect 9763 20102 9773 20154
rect 9773 20102 9819 20154
rect 9523 20100 9579 20102
rect 9603 20100 9659 20102
rect 9683 20100 9739 20102
rect 9763 20100 9819 20102
rect 9678 19236 9734 19272
rect 9678 19216 9680 19236
rect 9680 19216 9732 19236
rect 9732 19216 9734 19236
rect 9523 19066 9579 19068
rect 9603 19066 9659 19068
rect 9683 19066 9739 19068
rect 9763 19066 9819 19068
rect 9523 19014 9569 19066
rect 9569 19014 9579 19066
rect 9603 19014 9633 19066
rect 9633 19014 9645 19066
rect 9645 19014 9659 19066
rect 9683 19014 9697 19066
rect 9697 19014 9709 19066
rect 9709 19014 9739 19066
rect 9763 19014 9773 19066
rect 9773 19014 9819 19066
rect 9523 19012 9579 19014
rect 9603 19012 9659 19014
rect 9683 19012 9739 19014
rect 9763 19012 9819 19014
rect 9678 18808 9734 18864
rect 9523 17978 9579 17980
rect 9603 17978 9659 17980
rect 9683 17978 9739 17980
rect 9763 17978 9819 17980
rect 9523 17926 9569 17978
rect 9569 17926 9579 17978
rect 9603 17926 9633 17978
rect 9633 17926 9645 17978
rect 9645 17926 9659 17978
rect 9683 17926 9697 17978
rect 9697 17926 9709 17978
rect 9709 17926 9739 17978
rect 9763 17926 9773 17978
rect 9773 17926 9819 17978
rect 9523 17924 9579 17926
rect 9603 17924 9659 17926
rect 9683 17924 9739 17926
rect 9763 17924 9819 17926
rect 9523 16890 9579 16892
rect 9603 16890 9659 16892
rect 9683 16890 9739 16892
rect 9763 16890 9819 16892
rect 9523 16838 9569 16890
rect 9569 16838 9579 16890
rect 9603 16838 9633 16890
rect 9633 16838 9645 16890
rect 9645 16838 9659 16890
rect 9683 16838 9697 16890
rect 9697 16838 9709 16890
rect 9709 16838 9739 16890
rect 9763 16838 9773 16890
rect 9773 16838 9819 16890
rect 9523 16836 9579 16838
rect 9603 16836 9659 16838
rect 9683 16836 9739 16838
rect 9763 16836 9819 16838
rect 9523 15802 9579 15804
rect 9603 15802 9659 15804
rect 9683 15802 9739 15804
rect 9763 15802 9819 15804
rect 9523 15750 9569 15802
rect 9569 15750 9579 15802
rect 9603 15750 9633 15802
rect 9633 15750 9645 15802
rect 9645 15750 9659 15802
rect 9683 15750 9697 15802
rect 9697 15750 9709 15802
rect 9709 15750 9739 15802
rect 9763 15750 9773 15802
rect 9773 15750 9819 15802
rect 9523 15748 9579 15750
rect 9603 15748 9659 15750
rect 9683 15748 9739 15750
rect 9763 15748 9819 15750
rect 9523 14714 9579 14716
rect 9603 14714 9659 14716
rect 9683 14714 9739 14716
rect 9763 14714 9819 14716
rect 9523 14662 9569 14714
rect 9569 14662 9579 14714
rect 9603 14662 9633 14714
rect 9633 14662 9645 14714
rect 9645 14662 9659 14714
rect 9683 14662 9697 14714
rect 9697 14662 9709 14714
rect 9709 14662 9739 14714
rect 9763 14662 9773 14714
rect 9773 14662 9819 14714
rect 9523 14660 9579 14662
rect 9603 14660 9659 14662
rect 9683 14660 9739 14662
rect 9763 14660 9819 14662
rect 9523 13626 9579 13628
rect 9603 13626 9659 13628
rect 9683 13626 9739 13628
rect 9763 13626 9819 13628
rect 9523 13574 9569 13626
rect 9569 13574 9579 13626
rect 9603 13574 9633 13626
rect 9633 13574 9645 13626
rect 9645 13574 9659 13626
rect 9683 13574 9697 13626
rect 9697 13574 9709 13626
rect 9709 13574 9739 13626
rect 9763 13574 9773 13626
rect 9773 13574 9819 13626
rect 9523 13572 9579 13574
rect 9603 13572 9659 13574
rect 9683 13572 9739 13574
rect 9763 13572 9819 13574
rect 9770 12844 9826 12880
rect 9770 12824 9772 12844
rect 9772 12824 9824 12844
rect 9824 12824 9826 12844
rect 9523 12538 9579 12540
rect 9603 12538 9659 12540
rect 9683 12538 9739 12540
rect 9763 12538 9819 12540
rect 9523 12486 9569 12538
rect 9569 12486 9579 12538
rect 9603 12486 9633 12538
rect 9633 12486 9645 12538
rect 9645 12486 9659 12538
rect 9683 12486 9697 12538
rect 9697 12486 9709 12538
rect 9709 12486 9739 12538
rect 9763 12486 9773 12538
rect 9773 12486 9819 12538
rect 9523 12484 9579 12486
rect 9603 12484 9659 12486
rect 9683 12484 9739 12486
rect 9763 12484 9819 12486
rect 10138 18944 10194 19000
rect 10046 18672 10102 18728
rect 10230 15000 10286 15056
rect 9954 13368 10010 13424
rect 10230 14456 10286 14512
rect 9678 12280 9734 12336
rect 9954 12144 10010 12200
rect 9523 11450 9579 11452
rect 9603 11450 9659 11452
rect 9683 11450 9739 11452
rect 9763 11450 9819 11452
rect 9523 11398 9569 11450
rect 9569 11398 9579 11450
rect 9603 11398 9633 11450
rect 9633 11398 9645 11450
rect 9645 11398 9659 11450
rect 9683 11398 9697 11450
rect 9697 11398 9709 11450
rect 9709 11398 9739 11450
rect 9763 11398 9773 11450
rect 9773 11398 9819 11450
rect 9523 11396 9579 11398
rect 9603 11396 9659 11398
rect 9683 11396 9739 11398
rect 9763 11396 9819 11398
rect 9523 10362 9579 10364
rect 9603 10362 9659 10364
rect 9683 10362 9739 10364
rect 9763 10362 9819 10364
rect 9523 10310 9569 10362
rect 9569 10310 9579 10362
rect 9603 10310 9633 10362
rect 9633 10310 9645 10362
rect 9645 10310 9659 10362
rect 9683 10310 9697 10362
rect 9697 10310 9709 10362
rect 9709 10310 9739 10362
rect 9763 10310 9773 10362
rect 9773 10310 9819 10362
rect 9523 10308 9579 10310
rect 9603 10308 9659 10310
rect 9683 10308 9739 10310
rect 9763 10308 9819 10310
rect 9402 10104 9458 10160
rect 9310 9968 9366 10024
rect 10506 19252 10508 19272
rect 10508 19252 10560 19272
rect 10560 19252 10562 19272
rect 10506 19216 10562 19252
rect 11610 29824 11666 29880
rect 11236 29402 11292 29404
rect 11316 29402 11372 29404
rect 11396 29402 11452 29404
rect 11476 29402 11532 29404
rect 11236 29350 11282 29402
rect 11282 29350 11292 29402
rect 11316 29350 11346 29402
rect 11346 29350 11358 29402
rect 11358 29350 11372 29402
rect 11396 29350 11410 29402
rect 11410 29350 11422 29402
rect 11422 29350 11452 29402
rect 11476 29350 11486 29402
rect 11486 29350 11532 29402
rect 11236 29348 11292 29350
rect 11316 29348 11372 29350
rect 11396 29348 11452 29350
rect 11476 29348 11532 29350
rect 11236 28314 11292 28316
rect 11316 28314 11372 28316
rect 11396 28314 11452 28316
rect 11476 28314 11532 28316
rect 11236 28262 11282 28314
rect 11282 28262 11292 28314
rect 11316 28262 11346 28314
rect 11346 28262 11358 28314
rect 11358 28262 11372 28314
rect 11396 28262 11410 28314
rect 11410 28262 11422 28314
rect 11422 28262 11452 28314
rect 11476 28262 11486 28314
rect 11486 28262 11532 28314
rect 11236 28260 11292 28262
rect 11316 28260 11372 28262
rect 11396 28260 11452 28262
rect 11476 28260 11532 28262
rect 11236 27226 11292 27228
rect 11316 27226 11372 27228
rect 11396 27226 11452 27228
rect 11476 27226 11532 27228
rect 11236 27174 11282 27226
rect 11282 27174 11292 27226
rect 11316 27174 11346 27226
rect 11346 27174 11358 27226
rect 11358 27174 11372 27226
rect 11396 27174 11410 27226
rect 11410 27174 11422 27226
rect 11422 27174 11452 27226
rect 11476 27174 11486 27226
rect 11486 27174 11532 27226
rect 11236 27172 11292 27174
rect 11316 27172 11372 27174
rect 11396 27172 11452 27174
rect 11476 27172 11532 27174
rect 11236 26138 11292 26140
rect 11316 26138 11372 26140
rect 11396 26138 11452 26140
rect 11476 26138 11532 26140
rect 11236 26086 11282 26138
rect 11282 26086 11292 26138
rect 11316 26086 11346 26138
rect 11346 26086 11358 26138
rect 11358 26086 11372 26138
rect 11396 26086 11410 26138
rect 11410 26086 11422 26138
rect 11422 26086 11452 26138
rect 11476 26086 11486 26138
rect 11486 26086 11532 26138
rect 11236 26084 11292 26086
rect 11316 26084 11372 26086
rect 11396 26084 11452 26086
rect 11476 26084 11532 26086
rect 10506 18128 10562 18184
rect 11236 25050 11292 25052
rect 11316 25050 11372 25052
rect 11396 25050 11452 25052
rect 11476 25050 11532 25052
rect 11236 24998 11282 25050
rect 11282 24998 11292 25050
rect 11316 24998 11346 25050
rect 11346 24998 11358 25050
rect 11358 24998 11372 25050
rect 11396 24998 11410 25050
rect 11410 24998 11422 25050
rect 11422 24998 11452 25050
rect 11476 24998 11486 25050
rect 11486 24998 11532 25050
rect 11236 24996 11292 24998
rect 11316 24996 11372 24998
rect 11396 24996 11452 24998
rect 11476 24996 11532 24998
rect 11236 23962 11292 23964
rect 11316 23962 11372 23964
rect 11396 23962 11452 23964
rect 11476 23962 11532 23964
rect 11236 23910 11282 23962
rect 11282 23910 11292 23962
rect 11316 23910 11346 23962
rect 11346 23910 11358 23962
rect 11358 23910 11372 23962
rect 11396 23910 11410 23962
rect 11410 23910 11422 23962
rect 11422 23910 11452 23962
rect 11476 23910 11486 23962
rect 11486 23910 11532 23962
rect 11236 23908 11292 23910
rect 11316 23908 11372 23910
rect 11396 23908 11452 23910
rect 11476 23908 11532 23910
rect 11150 23160 11206 23216
rect 11236 22874 11292 22876
rect 11316 22874 11372 22876
rect 11396 22874 11452 22876
rect 11476 22874 11532 22876
rect 11236 22822 11282 22874
rect 11282 22822 11292 22874
rect 11316 22822 11346 22874
rect 11346 22822 11358 22874
rect 11358 22822 11372 22874
rect 11396 22822 11410 22874
rect 11410 22822 11422 22874
rect 11422 22822 11452 22874
rect 11476 22822 11486 22874
rect 11486 22822 11532 22874
rect 11236 22820 11292 22822
rect 11316 22820 11372 22822
rect 11396 22820 11452 22822
rect 11476 22820 11532 22822
rect 11058 21392 11114 21448
rect 11236 21786 11292 21788
rect 11316 21786 11372 21788
rect 11396 21786 11452 21788
rect 11476 21786 11532 21788
rect 11236 21734 11282 21786
rect 11282 21734 11292 21786
rect 11316 21734 11346 21786
rect 11346 21734 11358 21786
rect 11358 21734 11372 21786
rect 11396 21734 11410 21786
rect 11410 21734 11422 21786
rect 11422 21734 11452 21786
rect 11476 21734 11486 21786
rect 11486 21734 11532 21786
rect 11236 21732 11292 21734
rect 11316 21732 11372 21734
rect 11396 21732 11452 21734
rect 11476 21732 11532 21734
rect 11236 20698 11292 20700
rect 11316 20698 11372 20700
rect 11396 20698 11452 20700
rect 11476 20698 11532 20700
rect 11236 20646 11282 20698
rect 11282 20646 11292 20698
rect 11316 20646 11346 20698
rect 11346 20646 11358 20698
rect 11358 20646 11372 20698
rect 11396 20646 11410 20698
rect 11410 20646 11422 20698
rect 11422 20646 11452 20698
rect 11476 20646 11486 20698
rect 11486 20646 11532 20698
rect 11236 20644 11292 20646
rect 11316 20644 11372 20646
rect 11396 20644 11452 20646
rect 11476 20644 11532 20646
rect 11242 19760 11298 19816
rect 11518 19760 11574 19816
rect 11236 19610 11292 19612
rect 11316 19610 11372 19612
rect 11396 19610 11452 19612
rect 11476 19610 11532 19612
rect 11236 19558 11282 19610
rect 11282 19558 11292 19610
rect 11316 19558 11346 19610
rect 11346 19558 11358 19610
rect 11358 19558 11372 19610
rect 11396 19558 11410 19610
rect 11410 19558 11422 19610
rect 11422 19558 11452 19610
rect 11476 19558 11486 19610
rect 11486 19558 11532 19610
rect 11236 19556 11292 19558
rect 11316 19556 11372 19558
rect 11396 19556 11452 19558
rect 11476 19556 11532 19558
rect 11518 19352 11574 19408
rect 11242 19080 11298 19136
rect 10414 15408 10470 15464
rect 11058 17856 11114 17912
rect 10874 16768 10930 16824
rect 10782 16632 10838 16688
rect 11236 18522 11292 18524
rect 11316 18522 11372 18524
rect 11396 18522 11452 18524
rect 11476 18522 11532 18524
rect 11236 18470 11282 18522
rect 11282 18470 11292 18522
rect 11316 18470 11346 18522
rect 11346 18470 11358 18522
rect 11358 18470 11372 18522
rect 11396 18470 11410 18522
rect 11410 18470 11422 18522
rect 11422 18470 11452 18522
rect 11476 18470 11486 18522
rect 11486 18470 11532 18522
rect 11236 18468 11292 18470
rect 11316 18468 11372 18470
rect 11396 18468 11452 18470
rect 11476 18468 11532 18470
rect 11242 17720 11298 17776
rect 11426 17720 11482 17776
rect 11236 17434 11292 17436
rect 11316 17434 11372 17436
rect 11396 17434 11452 17436
rect 11476 17434 11532 17436
rect 11236 17382 11282 17434
rect 11282 17382 11292 17434
rect 11316 17382 11346 17434
rect 11346 17382 11358 17434
rect 11358 17382 11372 17434
rect 11396 17382 11410 17434
rect 11410 17382 11422 17434
rect 11422 17382 11452 17434
rect 11476 17382 11486 17434
rect 11486 17382 11532 17434
rect 11236 17380 11292 17382
rect 11316 17380 11372 17382
rect 11396 17380 11452 17382
rect 11476 17380 11532 17382
rect 14663 39194 14719 39196
rect 14743 39194 14799 39196
rect 14823 39194 14879 39196
rect 14903 39194 14959 39196
rect 14663 39142 14709 39194
rect 14709 39142 14719 39194
rect 14743 39142 14773 39194
rect 14773 39142 14785 39194
rect 14785 39142 14799 39194
rect 14823 39142 14837 39194
rect 14837 39142 14849 39194
rect 14849 39142 14879 39194
rect 14903 39142 14913 39194
rect 14913 39142 14959 39194
rect 14663 39140 14719 39142
rect 14743 39140 14799 39142
rect 14823 39140 14879 39142
rect 14903 39140 14959 39142
rect 14370 38664 14426 38720
rect 13634 38392 13690 38448
rect 14186 38392 14242 38448
rect 13450 38120 13506 38176
rect 13818 37848 13874 37904
rect 14370 37576 14426 37632
rect 14186 37304 14242 37360
rect 13634 37168 13690 37224
rect 13634 36760 13690 36816
rect 11794 27784 11850 27840
rect 11978 28872 12034 28928
rect 13266 35536 13322 35592
rect 12950 35386 13006 35388
rect 13030 35386 13086 35388
rect 13110 35386 13166 35388
rect 13190 35386 13246 35388
rect 12950 35334 12996 35386
rect 12996 35334 13006 35386
rect 13030 35334 13060 35386
rect 13060 35334 13072 35386
rect 13072 35334 13086 35386
rect 13110 35334 13124 35386
rect 13124 35334 13136 35386
rect 13136 35334 13166 35386
rect 13190 35334 13200 35386
rect 13200 35334 13246 35386
rect 12950 35332 13006 35334
rect 13030 35332 13086 35334
rect 13110 35332 13166 35334
rect 13190 35332 13246 35334
rect 12950 34298 13006 34300
rect 13030 34298 13086 34300
rect 13110 34298 13166 34300
rect 13190 34298 13246 34300
rect 12950 34246 12996 34298
rect 12996 34246 13006 34298
rect 13030 34246 13060 34298
rect 13060 34246 13072 34298
rect 13072 34246 13086 34298
rect 13110 34246 13124 34298
rect 13124 34246 13136 34298
rect 13136 34246 13166 34298
rect 13190 34246 13200 34298
rect 13200 34246 13246 34298
rect 12950 34244 13006 34246
rect 13030 34244 13086 34246
rect 13110 34244 13166 34246
rect 13190 34244 13246 34246
rect 12622 33088 12678 33144
rect 14370 36488 14426 36544
rect 13818 36216 13874 36272
rect 13726 35672 13782 35728
rect 13818 35128 13874 35184
rect 13542 35012 13598 35048
rect 13542 34992 13544 35012
rect 13544 34992 13596 35012
rect 13596 34992 13598 35012
rect 12622 31764 12624 31784
rect 12624 31764 12676 31784
rect 12676 31764 12678 31784
rect 12622 31728 12678 31764
rect 12438 31048 12494 31104
rect 12950 33210 13006 33212
rect 13030 33210 13086 33212
rect 13110 33210 13166 33212
rect 13190 33210 13246 33212
rect 12950 33158 12996 33210
rect 12996 33158 13006 33210
rect 13030 33158 13060 33210
rect 13060 33158 13072 33210
rect 13072 33158 13086 33210
rect 13110 33158 13124 33210
rect 13124 33158 13136 33210
rect 13136 33158 13166 33210
rect 13190 33158 13200 33210
rect 13200 33158 13246 33210
rect 12950 33156 13006 33158
rect 13030 33156 13086 33158
rect 13110 33156 13166 33158
rect 13190 33156 13246 33158
rect 12950 32122 13006 32124
rect 13030 32122 13086 32124
rect 13110 32122 13166 32124
rect 13190 32122 13246 32124
rect 12950 32070 12996 32122
rect 12996 32070 13006 32122
rect 13030 32070 13060 32122
rect 13060 32070 13072 32122
rect 13072 32070 13086 32122
rect 13110 32070 13124 32122
rect 13124 32070 13136 32122
rect 13136 32070 13166 32122
rect 13190 32070 13200 32122
rect 13200 32070 13246 32122
rect 12950 32068 13006 32070
rect 13030 32068 13086 32070
rect 13110 32068 13166 32070
rect 13190 32068 13246 32070
rect 12990 31320 13046 31376
rect 13910 34584 13966 34640
rect 13634 34040 13690 34096
rect 13634 32952 13690 33008
rect 13542 32272 13598 32328
rect 13450 31184 13506 31240
rect 13726 31864 13782 31920
rect 13358 31048 13414 31104
rect 12950 31034 13006 31036
rect 13030 31034 13086 31036
rect 13110 31034 13166 31036
rect 13190 31034 13246 31036
rect 12950 30982 12996 31034
rect 12996 30982 13006 31034
rect 13030 30982 13060 31034
rect 13060 30982 13072 31034
rect 13072 30982 13086 31034
rect 13110 30982 13124 31034
rect 13124 30982 13136 31034
rect 13136 30982 13166 31034
rect 13190 30982 13200 31034
rect 13200 30982 13246 31034
rect 12950 30980 13006 30982
rect 13030 30980 13086 30982
rect 13110 30980 13166 30982
rect 13190 30980 13246 30982
rect 12898 30232 12954 30288
rect 13358 30232 13414 30288
rect 12950 29946 13006 29948
rect 13030 29946 13086 29948
rect 13110 29946 13166 29948
rect 13190 29946 13246 29948
rect 12950 29894 12996 29946
rect 12996 29894 13006 29946
rect 13030 29894 13060 29946
rect 13060 29894 13072 29946
rect 13072 29894 13086 29946
rect 13110 29894 13124 29946
rect 13124 29894 13136 29946
rect 13136 29894 13166 29946
rect 13190 29894 13200 29946
rect 13200 29894 13246 29946
rect 12950 29892 13006 29894
rect 13030 29892 13086 29894
rect 13110 29892 13166 29894
rect 13190 29892 13246 29894
rect 12898 29164 12954 29200
rect 12898 29144 12900 29164
rect 12900 29144 12952 29164
rect 12952 29144 12954 29164
rect 12162 26424 12218 26480
rect 12530 26968 12586 27024
rect 12346 25880 12402 25936
rect 12950 28858 13006 28860
rect 13030 28858 13086 28860
rect 13110 28858 13166 28860
rect 13190 28858 13246 28860
rect 12950 28806 12996 28858
rect 12996 28806 13006 28858
rect 13030 28806 13060 28858
rect 13060 28806 13072 28858
rect 13072 28806 13086 28858
rect 13110 28806 13124 28858
rect 13124 28806 13136 28858
rect 13136 28806 13166 28858
rect 13190 28806 13200 28858
rect 13200 28806 13246 28858
rect 12950 28804 13006 28806
rect 13030 28804 13086 28806
rect 13110 28804 13166 28806
rect 13190 28804 13246 28806
rect 12950 27770 13006 27772
rect 13030 27770 13086 27772
rect 13110 27770 13166 27772
rect 13190 27770 13246 27772
rect 12950 27718 12996 27770
rect 12996 27718 13006 27770
rect 13030 27718 13060 27770
rect 13060 27718 13072 27770
rect 13072 27718 13086 27770
rect 13110 27718 13124 27770
rect 13124 27718 13136 27770
rect 13136 27718 13166 27770
rect 13190 27718 13200 27770
rect 13200 27718 13246 27770
rect 12950 27716 13006 27718
rect 13030 27716 13086 27718
rect 13110 27716 13166 27718
rect 13190 27716 13246 27718
rect 12990 27240 13046 27296
rect 13910 33496 13966 33552
rect 14370 34312 14426 34368
rect 14186 34040 14242 34096
rect 14186 32952 14242 33008
rect 14370 33224 14426 33280
rect 14278 32408 14334 32464
rect 13910 31864 13966 31920
rect 14002 31320 14058 31376
rect 13910 30776 13966 30832
rect 13634 29688 13690 29744
rect 13910 29552 13966 29608
rect 13634 28600 13690 28656
rect 13818 28056 13874 28112
rect 13358 26968 13414 27024
rect 12950 26682 13006 26684
rect 13030 26682 13086 26684
rect 13110 26682 13166 26684
rect 13190 26682 13246 26684
rect 12950 26630 12996 26682
rect 12996 26630 13006 26682
rect 13030 26630 13060 26682
rect 13060 26630 13072 26682
rect 13072 26630 13086 26682
rect 13110 26630 13124 26682
rect 13124 26630 13136 26682
rect 13136 26630 13166 26682
rect 13190 26630 13200 26682
rect 13200 26630 13246 26682
rect 12950 26628 13006 26630
rect 13030 26628 13086 26630
rect 13110 26628 13166 26630
rect 13190 26628 13246 26630
rect 13266 26152 13322 26208
rect 12806 26016 12862 26072
rect 13634 27512 13690 27568
rect 13910 26968 13966 27024
rect 14370 32172 14372 32192
rect 14372 32172 14424 32192
rect 14424 32172 14426 32192
rect 14370 32136 14426 32172
rect 14278 29144 14334 29200
rect 14186 28600 14242 28656
rect 14186 27512 14242 27568
rect 14370 27784 14426 27840
rect 13818 26732 13820 26752
rect 13820 26732 13872 26752
rect 13872 26732 13874 26752
rect 13818 26696 13874 26732
rect 12950 25594 13006 25596
rect 13030 25594 13086 25596
rect 13110 25594 13166 25596
rect 13190 25594 13246 25596
rect 12950 25542 12996 25594
rect 12996 25542 13006 25594
rect 13030 25542 13060 25594
rect 13060 25542 13072 25594
rect 13072 25542 13086 25594
rect 13110 25542 13124 25594
rect 13124 25542 13136 25594
rect 13136 25542 13166 25594
rect 13190 25542 13200 25594
rect 13200 25542 13246 25594
rect 12950 25540 13006 25542
rect 13030 25540 13086 25542
rect 13110 25540 13166 25542
rect 13190 25540 13246 25542
rect 12070 23840 12126 23896
rect 11794 20712 11850 20768
rect 11236 16346 11292 16348
rect 11316 16346 11372 16348
rect 11396 16346 11452 16348
rect 11476 16346 11532 16348
rect 11236 16294 11282 16346
rect 11282 16294 11292 16346
rect 11316 16294 11346 16346
rect 11346 16294 11358 16346
rect 11358 16294 11372 16346
rect 11396 16294 11410 16346
rect 11410 16294 11422 16346
rect 11422 16294 11452 16346
rect 11476 16294 11486 16346
rect 11486 16294 11532 16346
rect 11236 16292 11292 16294
rect 11316 16292 11372 16294
rect 11396 16292 11452 16294
rect 11476 16292 11532 16294
rect 11518 15544 11574 15600
rect 11236 15258 11292 15260
rect 11316 15258 11372 15260
rect 11396 15258 11452 15260
rect 11476 15258 11532 15260
rect 11236 15206 11282 15258
rect 11282 15206 11292 15258
rect 11316 15206 11346 15258
rect 11346 15206 11358 15258
rect 11358 15206 11372 15258
rect 11396 15206 11410 15258
rect 11410 15206 11422 15258
rect 11422 15206 11452 15258
rect 11476 15206 11486 15258
rect 11486 15206 11532 15258
rect 11236 15204 11292 15206
rect 11316 15204 11372 15206
rect 11396 15204 11452 15206
rect 11476 15204 11532 15206
rect 11150 14864 11206 14920
rect 11236 14170 11292 14172
rect 11316 14170 11372 14172
rect 11396 14170 11452 14172
rect 11476 14170 11532 14172
rect 11236 14118 11282 14170
rect 11282 14118 11292 14170
rect 11316 14118 11346 14170
rect 11346 14118 11358 14170
rect 11358 14118 11372 14170
rect 11396 14118 11410 14170
rect 11410 14118 11422 14170
rect 11422 14118 11452 14170
rect 11476 14118 11486 14170
rect 11486 14118 11532 14170
rect 11236 14116 11292 14118
rect 11316 14116 11372 14118
rect 11396 14116 11452 14118
rect 11476 14116 11532 14118
rect 9954 10512 10010 10568
rect 10782 12280 10838 12336
rect 10230 10240 10286 10296
rect 9523 9274 9579 9276
rect 9603 9274 9659 9276
rect 9683 9274 9739 9276
rect 9763 9274 9819 9276
rect 9523 9222 9569 9274
rect 9569 9222 9579 9274
rect 9603 9222 9633 9274
rect 9633 9222 9645 9274
rect 9645 9222 9659 9274
rect 9683 9222 9697 9274
rect 9697 9222 9709 9274
rect 9709 9222 9739 9274
rect 9763 9222 9773 9274
rect 9773 9222 9819 9274
rect 9523 9220 9579 9222
rect 9603 9220 9659 9222
rect 9683 9220 9739 9222
rect 9763 9220 9819 9222
rect 10230 9560 10286 9616
rect 9678 8880 9734 8936
rect 9494 8744 9550 8800
rect 9523 8186 9579 8188
rect 9603 8186 9659 8188
rect 9683 8186 9739 8188
rect 9763 8186 9819 8188
rect 9523 8134 9569 8186
rect 9569 8134 9579 8186
rect 9603 8134 9633 8186
rect 9633 8134 9645 8186
rect 9645 8134 9659 8186
rect 9683 8134 9697 8186
rect 9697 8134 9709 8186
rect 9709 8134 9739 8186
rect 9763 8134 9773 8186
rect 9773 8134 9819 8186
rect 9523 8132 9579 8134
rect 9603 8132 9659 8134
rect 9683 8132 9739 8134
rect 9763 8132 9819 8134
rect 9770 7948 9826 7984
rect 9770 7928 9772 7948
rect 9772 7928 9824 7948
rect 9824 7928 9826 7948
rect 9586 7792 9642 7848
rect 9523 7098 9579 7100
rect 9603 7098 9659 7100
rect 9683 7098 9739 7100
rect 9763 7098 9819 7100
rect 9523 7046 9569 7098
rect 9569 7046 9579 7098
rect 9603 7046 9633 7098
rect 9633 7046 9645 7098
rect 9645 7046 9659 7098
rect 9683 7046 9697 7098
rect 9697 7046 9709 7098
rect 9709 7046 9739 7098
rect 9763 7046 9773 7098
rect 9773 7046 9819 7098
rect 9523 7044 9579 7046
rect 9603 7044 9659 7046
rect 9683 7044 9739 7046
rect 9763 7044 9819 7046
rect 10506 9832 10562 9888
rect 10414 9288 10470 9344
rect 10322 9152 10378 9208
rect 10138 8472 10194 8528
rect 10690 8744 10746 8800
rect 11426 13232 11482 13288
rect 11236 13082 11292 13084
rect 11316 13082 11372 13084
rect 11396 13082 11452 13084
rect 11476 13082 11532 13084
rect 11236 13030 11282 13082
rect 11282 13030 11292 13082
rect 11316 13030 11346 13082
rect 11346 13030 11358 13082
rect 11358 13030 11372 13082
rect 11396 13030 11410 13082
rect 11410 13030 11422 13082
rect 11422 13030 11452 13082
rect 11476 13030 11486 13082
rect 11486 13030 11532 13082
rect 11236 13028 11292 13030
rect 11316 13028 11372 13030
rect 11396 13028 11452 13030
rect 11476 13028 11532 13030
rect 12070 21936 12126 21992
rect 11794 19080 11850 19136
rect 12950 24506 13006 24508
rect 13030 24506 13086 24508
rect 13110 24506 13166 24508
rect 13190 24506 13246 24508
rect 12950 24454 12996 24506
rect 12996 24454 13006 24506
rect 13030 24454 13060 24506
rect 13060 24454 13072 24506
rect 13072 24454 13086 24506
rect 13110 24454 13124 24506
rect 13124 24454 13136 24506
rect 13136 24454 13166 24506
rect 13190 24454 13200 24506
rect 13200 24454 13246 24506
rect 12950 24452 13006 24454
rect 13030 24452 13086 24454
rect 13110 24452 13166 24454
rect 13190 24452 13246 24454
rect 12950 23418 13006 23420
rect 13030 23418 13086 23420
rect 13110 23418 13166 23420
rect 13190 23418 13246 23420
rect 12950 23366 12996 23418
rect 12996 23366 13006 23418
rect 13030 23366 13060 23418
rect 13060 23366 13072 23418
rect 13072 23366 13086 23418
rect 13110 23366 13124 23418
rect 13124 23366 13136 23418
rect 13136 23366 13166 23418
rect 13190 23366 13200 23418
rect 13200 23366 13246 23418
rect 12950 23364 13006 23366
rect 13030 23364 13086 23366
rect 13110 23364 13166 23366
rect 13190 23364 13246 23366
rect 12438 20340 12440 20360
rect 12440 20340 12492 20360
rect 12492 20340 12494 20360
rect 12438 20304 12494 20340
rect 12254 19352 12310 19408
rect 11794 15816 11850 15872
rect 11610 12300 11666 12336
rect 11610 12280 11612 12300
rect 11612 12280 11664 12300
rect 11664 12280 11666 12300
rect 11236 11994 11292 11996
rect 11316 11994 11372 11996
rect 11396 11994 11452 11996
rect 11476 11994 11532 11996
rect 11236 11942 11282 11994
rect 11282 11942 11292 11994
rect 11316 11942 11346 11994
rect 11346 11942 11358 11994
rect 11358 11942 11372 11994
rect 11396 11942 11410 11994
rect 11410 11942 11422 11994
rect 11422 11942 11452 11994
rect 11476 11942 11486 11994
rect 11486 11942 11532 11994
rect 11236 11940 11292 11942
rect 11316 11940 11372 11942
rect 11396 11940 11452 11942
rect 11476 11940 11532 11942
rect 10966 9560 11022 9616
rect 11794 12280 11850 12336
rect 11236 10906 11292 10908
rect 11316 10906 11372 10908
rect 11396 10906 11452 10908
rect 11476 10906 11532 10908
rect 11236 10854 11282 10906
rect 11282 10854 11292 10906
rect 11316 10854 11346 10906
rect 11346 10854 11358 10906
rect 11358 10854 11372 10906
rect 11396 10854 11410 10906
rect 11410 10854 11422 10906
rect 11422 10854 11452 10906
rect 11476 10854 11486 10906
rect 11486 10854 11532 10906
rect 11236 10852 11292 10854
rect 11316 10852 11372 10854
rect 11396 10852 11452 10854
rect 11476 10852 11532 10854
rect 11236 9818 11292 9820
rect 11316 9818 11372 9820
rect 11396 9818 11452 9820
rect 11476 9818 11532 9820
rect 11236 9766 11282 9818
rect 11282 9766 11292 9818
rect 11316 9766 11346 9818
rect 11346 9766 11358 9818
rect 11358 9766 11372 9818
rect 11396 9766 11410 9818
rect 11410 9766 11422 9818
rect 11422 9766 11452 9818
rect 11476 9766 11486 9818
rect 11486 9766 11532 9818
rect 11236 9764 11292 9766
rect 11316 9764 11372 9766
rect 11396 9764 11452 9766
rect 11476 9764 11532 9766
rect 11334 9580 11390 9616
rect 11334 9560 11336 9580
rect 11336 9560 11388 9580
rect 11388 9560 11390 9580
rect 11058 9288 11114 9344
rect 10138 8200 10194 8256
rect 10322 8200 10378 8256
rect 9523 6010 9579 6012
rect 9603 6010 9659 6012
rect 9683 6010 9739 6012
rect 9763 6010 9819 6012
rect 9523 5958 9569 6010
rect 9569 5958 9579 6010
rect 9603 5958 9633 6010
rect 9633 5958 9645 6010
rect 9645 5958 9659 6010
rect 9683 5958 9697 6010
rect 9697 5958 9709 6010
rect 9709 5958 9739 6010
rect 9763 5958 9773 6010
rect 9773 5958 9819 6010
rect 9523 5956 9579 5958
rect 9603 5956 9659 5958
rect 9683 5956 9739 5958
rect 9763 5956 9819 5958
rect 11334 9288 11390 9344
rect 11518 9288 11574 9344
rect 11242 8916 11244 8936
rect 11244 8916 11296 8936
rect 11296 8916 11298 8936
rect 11242 8880 11298 8916
rect 11236 8730 11292 8732
rect 11316 8730 11372 8732
rect 11396 8730 11452 8732
rect 11476 8730 11532 8732
rect 11236 8678 11282 8730
rect 11282 8678 11292 8730
rect 11316 8678 11346 8730
rect 11346 8678 11358 8730
rect 11358 8678 11372 8730
rect 11396 8678 11410 8730
rect 11410 8678 11422 8730
rect 11422 8678 11452 8730
rect 11476 8678 11486 8730
rect 11486 8678 11532 8730
rect 11236 8676 11292 8678
rect 11316 8676 11372 8678
rect 11396 8676 11452 8678
rect 11476 8676 11532 8678
rect 11702 9832 11758 9888
rect 11794 9696 11850 9752
rect 12070 16496 12126 16552
rect 12254 16496 12310 16552
rect 12622 20884 12624 20904
rect 12624 20884 12676 20904
rect 12676 20884 12678 20904
rect 12622 20848 12678 20884
rect 12346 15544 12402 15600
rect 12438 15136 12494 15192
rect 12714 18944 12770 19000
rect 12950 22330 13006 22332
rect 13030 22330 13086 22332
rect 13110 22330 13166 22332
rect 13190 22330 13246 22332
rect 12950 22278 12996 22330
rect 12996 22278 13006 22330
rect 13030 22278 13060 22330
rect 13060 22278 13072 22330
rect 13072 22278 13086 22330
rect 13110 22278 13124 22330
rect 13124 22278 13136 22330
rect 13136 22278 13166 22330
rect 13190 22278 13200 22330
rect 13200 22278 13246 22330
rect 12950 22276 13006 22278
rect 13030 22276 13086 22278
rect 13110 22276 13166 22278
rect 13190 22276 13246 22278
rect 13450 23060 13452 23080
rect 13452 23060 13504 23080
rect 13504 23060 13506 23080
rect 13450 23024 13506 23060
rect 12950 21242 13006 21244
rect 13030 21242 13086 21244
rect 13110 21242 13166 21244
rect 13190 21242 13246 21244
rect 12950 21190 12996 21242
rect 12996 21190 13006 21242
rect 13030 21190 13060 21242
rect 13060 21190 13072 21242
rect 13072 21190 13086 21242
rect 13110 21190 13124 21242
rect 13124 21190 13136 21242
rect 13136 21190 13166 21242
rect 13190 21190 13200 21242
rect 13200 21190 13246 21242
rect 12950 21188 13006 21190
rect 13030 21188 13086 21190
rect 13110 21188 13166 21190
rect 13190 21188 13246 21190
rect 13450 22208 13506 22264
rect 13818 25336 13874 25392
rect 13726 24656 13782 24712
rect 13726 22344 13782 22400
rect 14663 38106 14719 38108
rect 14743 38106 14799 38108
rect 14823 38106 14879 38108
rect 14903 38106 14959 38108
rect 14663 38054 14709 38106
rect 14709 38054 14719 38106
rect 14743 38054 14773 38106
rect 14773 38054 14785 38106
rect 14785 38054 14799 38106
rect 14823 38054 14837 38106
rect 14837 38054 14849 38106
rect 14849 38054 14879 38106
rect 14903 38054 14913 38106
rect 14913 38054 14959 38106
rect 14663 38052 14719 38054
rect 14743 38052 14799 38054
rect 14823 38052 14879 38054
rect 14903 38052 14959 38054
rect 14663 37018 14719 37020
rect 14743 37018 14799 37020
rect 14823 37018 14879 37020
rect 14903 37018 14959 37020
rect 14663 36966 14709 37018
rect 14709 36966 14719 37018
rect 14743 36966 14773 37018
rect 14773 36966 14785 37018
rect 14785 36966 14799 37018
rect 14823 36966 14837 37018
rect 14837 36966 14849 37018
rect 14849 36966 14879 37018
rect 14903 36966 14913 37018
rect 14913 36966 14959 37018
rect 14663 36964 14719 36966
rect 14743 36964 14799 36966
rect 14823 36964 14879 36966
rect 14903 36964 14959 36966
rect 14663 35930 14719 35932
rect 14743 35930 14799 35932
rect 14823 35930 14879 35932
rect 14903 35930 14959 35932
rect 14663 35878 14709 35930
rect 14709 35878 14719 35930
rect 14743 35878 14773 35930
rect 14773 35878 14785 35930
rect 14785 35878 14799 35930
rect 14823 35878 14837 35930
rect 14837 35878 14849 35930
rect 14849 35878 14879 35930
rect 14903 35878 14913 35930
rect 14913 35878 14959 35930
rect 14663 35876 14719 35878
rect 14743 35876 14799 35878
rect 14823 35876 14879 35878
rect 14903 35876 14959 35878
rect 14663 34842 14719 34844
rect 14743 34842 14799 34844
rect 14823 34842 14879 34844
rect 14903 34842 14959 34844
rect 14663 34790 14709 34842
rect 14709 34790 14719 34842
rect 14743 34790 14773 34842
rect 14773 34790 14785 34842
rect 14785 34790 14799 34842
rect 14823 34790 14837 34842
rect 14837 34790 14849 34842
rect 14849 34790 14879 34842
rect 14903 34790 14913 34842
rect 14913 34790 14959 34842
rect 14663 34788 14719 34790
rect 14743 34788 14799 34790
rect 14823 34788 14879 34790
rect 14903 34788 14959 34790
rect 14663 33754 14719 33756
rect 14743 33754 14799 33756
rect 14823 33754 14879 33756
rect 14903 33754 14959 33756
rect 14663 33702 14709 33754
rect 14709 33702 14719 33754
rect 14743 33702 14773 33754
rect 14773 33702 14785 33754
rect 14785 33702 14799 33754
rect 14823 33702 14837 33754
rect 14837 33702 14849 33754
rect 14849 33702 14879 33754
rect 14903 33702 14913 33754
rect 14913 33702 14959 33754
rect 14663 33700 14719 33702
rect 14743 33700 14799 33702
rect 14823 33700 14879 33702
rect 14903 33700 14959 33702
rect 14663 32666 14719 32668
rect 14743 32666 14799 32668
rect 14823 32666 14879 32668
rect 14903 32666 14959 32668
rect 14663 32614 14709 32666
rect 14709 32614 14719 32666
rect 14743 32614 14773 32666
rect 14773 32614 14785 32666
rect 14785 32614 14799 32666
rect 14823 32614 14837 32666
rect 14837 32614 14849 32666
rect 14849 32614 14879 32666
rect 14903 32614 14913 32666
rect 14913 32614 14959 32666
rect 14663 32612 14719 32614
rect 14743 32612 14799 32614
rect 14823 32612 14879 32614
rect 14903 32612 14959 32614
rect 14663 31578 14719 31580
rect 14743 31578 14799 31580
rect 14823 31578 14879 31580
rect 14903 31578 14959 31580
rect 14663 31526 14709 31578
rect 14709 31526 14719 31578
rect 14743 31526 14773 31578
rect 14773 31526 14785 31578
rect 14785 31526 14799 31578
rect 14823 31526 14837 31578
rect 14837 31526 14849 31578
rect 14849 31526 14879 31578
rect 14903 31526 14913 31578
rect 14913 31526 14959 31578
rect 14663 31524 14719 31526
rect 14743 31524 14799 31526
rect 14823 31524 14879 31526
rect 14903 31524 14959 31526
rect 14663 30490 14719 30492
rect 14743 30490 14799 30492
rect 14823 30490 14879 30492
rect 14903 30490 14959 30492
rect 14663 30438 14709 30490
rect 14709 30438 14719 30490
rect 14743 30438 14773 30490
rect 14773 30438 14785 30490
rect 14785 30438 14799 30490
rect 14823 30438 14837 30490
rect 14837 30438 14849 30490
rect 14849 30438 14879 30490
rect 14903 30438 14913 30490
rect 14913 30438 14959 30490
rect 14663 30436 14719 30438
rect 14743 30436 14799 30438
rect 14823 30436 14879 30438
rect 14903 30436 14959 30438
rect 14663 29402 14719 29404
rect 14743 29402 14799 29404
rect 14823 29402 14879 29404
rect 14903 29402 14959 29404
rect 14663 29350 14709 29402
rect 14709 29350 14719 29402
rect 14743 29350 14773 29402
rect 14773 29350 14785 29402
rect 14785 29350 14799 29402
rect 14823 29350 14837 29402
rect 14837 29350 14849 29402
rect 14849 29350 14879 29402
rect 14903 29350 14913 29402
rect 14913 29350 14959 29402
rect 14663 29348 14719 29350
rect 14743 29348 14799 29350
rect 14823 29348 14879 29350
rect 14903 29348 14959 29350
rect 14554 28872 14610 28928
rect 14370 25200 14426 25256
rect 14186 24556 14188 24576
rect 14188 24556 14240 24576
rect 14240 24556 14242 24576
rect 14186 24520 14242 24556
rect 14370 24248 14426 24304
rect 14370 23704 14426 23760
rect 14370 23468 14372 23488
rect 14372 23468 14424 23488
rect 14424 23468 14426 23488
rect 14370 23432 14426 23468
rect 14370 23196 14372 23216
rect 14372 23196 14424 23216
rect 14424 23196 14426 23216
rect 14370 23160 14426 23196
rect 12950 20154 13006 20156
rect 13030 20154 13086 20156
rect 13110 20154 13166 20156
rect 13190 20154 13246 20156
rect 12950 20102 12996 20154
rect 12996 20102 13006 20154
rect 13030 20102 13060 20154
rect 13060 20102 13072 20154
rect 13072 20102 13086 20154
rect 13110 20102 13124 20154
rect 13124 20102 13136 20154
rect 13136 20102 13166 20154
rect 13190 20102 13200 20154
rect 13200 20102 13246 20154
rect 12950 20100 13006 20102
rect 13030 20100 13086 20102
rect 13110 20100 13166 20102
rect 13190 20100 13246 20102
rect 12950 19066 13006 19068
rect 13030 19066 13086 19068
rect 13110 19066 13166 19068
rect 13190 19066 13246 19068
rect 12950 19014 12996 19066
rect 12996 19014 13006 19066
rect 13030 19014 13060 19066
rect 13060 19014 13072 19066
rect 13072 19014 13086 19066
rect 13110 19014 13124 19066
rect 13124 19014 13136 19066
rect 13136 19014 13166 19066
rect 13190 19014 13200 19066
rect 13200 19014 13246 19066
rect 12950 19012 13006 19014
rect 13030 19012 13086 19014
rect 13110 19012 13166 19014
rect 13190 19012 13246 19014
rect 12806 18808 12862 18864
rect 13174 18672 13230 18728
rect 13174 18128 13230 18184
rect 12950 17978 13006 17980
rect 13030 17978 13086 17980
rect 13110 17978 13166 17980
rect 13190 17978 13246 17980
rect 12950 17926 12996 17978
rect 12996 17926 13006 17978
rect 13030 17926 13060 17978
rect 13060 17926 13072 17978
rect 13072 17926 13086 17978
rect 13110 17926 13124 17978
rect 13124 17926 13136 17978
rect 13136 17926 13166 17978
rect 13190 17926 13200 17978
rect 13200 17926 13246 17978
rect 12950 17924 13006 17926
rect 13030 17924 13086 17926
rect 13110 17924 13166 17926
rect 13190 17924 13246 17926
rect 12950 16890 13006 16892
rect 13030 16890 13086 16892
rect 13110 16890 13166 16892
rect 13190 16890 13246 16892
rect 12950 16838 12996 16890
rect 12996 16838 13006 16890
rect 13030 16838 13060 16890
rect 13060 16838 13072 16890
rect 13072 16838 13086 16890
rect 13110 16838 13124 16890
rect 13124 16838 13136 16890
rect 13136 16838 13166 16890
rect 13190 16838 13200 16890
rect 13200 16838 13246 16890
rect 12950 16836 13006 16838
rect 13030 16836 13086 16838
rect 13110 16836 13166 16838
rect 13190 16836 13246 16838
rect 12714 16788 12770 16824
rect 12714 16768 12716 16788
rect 12716 16768 12768 16788
rect 12768 16768 12770 16788
rect 12990 16632 13046 16688
rect 13726 21256 13782 21312
rect 13542 21120 13598 21176
rect 13358 17992 13414 18048
rect 12714 16108 12770 16144
rect 12714 16088 12716 16108
rect 12716 16088 12768 16108
rect 12768 16088 12770 16108
rect 11978 10376 12034 10432
rect 11978 10104 12034 10160
rect 12346 13232 12402 13288
rect 12530 13812 12532 13832
rect 12532 13812 12584 13832
rect 12584 13812 12586 13832
rect 12530 13776 12586 13812
rect 12254 12552 12310 12608
rect 13082 16224 13138 16280
rect 12714 14864 12770 14920
rect 12622 12416 12678 12472
rect 12622 11736 12678 11792
rect 12346 11192 12402 11248
rect 12950 15802 13006 15804
rect 13030 15802 13086 15804
rect 13110 15802 13166 15804
rect 13190 15802 13246 15804
rect 12950 15750 12996 15802
rect 12996 15750 13006 15802
rect 13030 15750 13060 15802
rect 13060 15750 13072 15802
rect 13072 15750 13086 15802
rect 13110 15750 13124 15802
rect 13124 15750 13136 15802
rect 13136 15750 13166 15802
rect 13190 15750 13200 15802
rect 13200 15750 13246 15802
rect 12950 15748 13006 15750
rect 13030 15748 13086 15750
rect 13110 15748 13166 15750
rect 13190 15748 13246 15750
rect 12898 15000 12954 15056
rect 13634 20168 13690 20224
rect 13818 20984 13874 21040
rect 14462 22344 14518 22400
rect 14462 22072 14518 22128
rect 14278 21528 14334 21584
rect 14094 20440 14150 20496
rect 12950 14714 13006 14716
rect 13030 14714 13086 14716
rect 13110 14714 13166 14716
rect 13190 14714 13246 14716
rect 12950 14662 12996 14714
rect 12996 14662 13006 14714
rect 13030 14662 13060 14714
rect 13060 14662 13072 14714
rect 13072 14662 13086 14714
rect 13110 14662 13124 14714
rect 13124 14662 13136 14714
rect 13136 14662 13166 14714
rect 13190 14662 13200 14714
rect 13200 14662 13246 14714
rect 12950 14660 13006 14662
rect 13030 14660 13086 14662
rect 13110 14660 13166 14662
rect 13190 14660 13246 14662
rect 12950 13626 13006 13628
rect 13030 13626 13086 13628
rect 13110 13626 13166 13628
rect 13190 13626 13246 13628
rect 12950 13574 12996 13626
rect 12996 13574 13006 13626
rect 13030 13574 13060 13626
rect 13060 13574 13072 13626
rect 13072 13574 13086 13626
rect 13110 13574 13124 13626
rect 13124 13574 13136 13626
rect 13136 13574 13166 13626
rect 13190 13574 13200 13626
rect 13200 13574 13246 13626
rect 12950 13572 13006 13574
rect 13030 13572 13086 13574
rect 13110 13572 13166 13574
rect 13190 13572 13246 13574
rect 13634 17040 13690 17096
rect 13542 16088 13598 16144
rect 13818 16904 13874 16960
rect 13818 16224 13874 16280
rect 13542 15272 13598 15328
rect 13726 15816 13782 15872
rect 13634 14592 13690 14648
rect 13082 13388 13138 13424
rect 13082 13368 13084 13388
rect 13084 13368 13136 13388
rect 13136 13368 13138 13388
rect 13082 13232 13138 13288
rect 13266 13096 13322 13152
rect 13082 12824 13138 12880
rect 12950 12538 13006 12540
rect 13030 12538 13086 12540
rect 13110 12538 13166 12540
rect 13190 12538 13246 12540
rect 12950 12486 12996 12538
rect 12996 12486 13006 12538
rect 13030 12486 13060 12538
rect 13060 12486 13072 12538
rect 13072 12486 13086 12538
rect 13110 12486 13124 12538
rect 13124 12486 13136 12538
rect 13136 12486 13166 12538
rect 13190 12486 13200 12538
rect 13200 12486 13246 12538
rect 12950 12484 13006 12486
rect 13030 12484 13086 12486
rect 13110 12484 13166 12486
rect 13190 12484 13246 12486
rect 13726 13812 13728 13832
rect 13728 13812 13780 13832
rect 13780 13812 13782 13832
rect 13726 13776 13782 13812
rect 13634 13640 13690 13696
rect 12950 11450 13006 11452
rect 13030 11450 13086 11452
rect 13110 11450 13166 11452
rect 13190 11450 13246 11452
rect 12950 11398 12996 11450
rect 12996 11398 13006 11450
rect 13030 11398 13060 11450
rect 13060 11398 13072 11450
rect 13072 11398 13086 11450
rect 13110 11398 13124 11450
rect 13124 11398 13136 11450
rect 13136 11398 13166 11450
rect 13190 11398 13200 11450
rect 13200 11398 13246 11450
rect 12950 11396 13006 11398
rect 13030 11396 13086 11398
rect 13110 11396 13166 11398
rect 13190 11396 13246 11398
rect 11978 9152 12034 9208
rect 11702 9016 11758 9072
rect 10598 7792 10654 7848
rect 9770 5616 9826 5672
rect 9523 4922 9579 4924
rect 9603 4922 9659 4924
rect 9683 4922 9739 4924
rect 9763 4922 9819 4924
rect 9523 4870 9569 4922
rect 9569 4870 9579 4922
rect 9603 4870 9633 4922
rect 9633 4870 9645 4922
rect 9645 4870 9659 4922
rect 9683 4870 9697 4922
rect 9697 4870 9709 4922
rect 9709 4870 9739 4922
rect 9763 4870 9773 4922
rect 9773 4870 9819 4922
rect 9523 4868 9579 4870
rect 9603 4868 9659 4870
rect 9683 4868 9739 4870
rect 9763 4868 9819 4870
rect 10966 5208 11022 5264
rect 11242 7964 11244 7984
rect 11244 7964 11296 7984
rect 11296 7964 11298 7984
rect 11242 7928 11298 7964
rect 11236 7642 11292 7644
rect 11316 7642 11372 7644
rect 11396 7642 11452 7644
rect 11476 7642 11532 7644
rect 11236 7590 11282 7642
rect 11282 7590 11292 7642
rect 11316 7590 11346 7642
rect 11346 7590 11358 7642
rect 11358 7590 11372 7642
rect 11396 7590 11410 7642
rect 11410 7590 11422 7642
rect 11422 7590 11452 7642
rect 11476 7590 11486 7642
rect 11486 7590 11532 7642
rect 11236 7588 11292 7590
rect 11316 7588 11372 7590
rect 11396 7588 11452 7590
rect 11476 7588 11532 7590
rect 11236 6554 11292 6556
rect 11316 6554 11372 6556
rect 11396 6554 11452 6556
rect 11476 6554 11532 6556
rect 11236 6502 11282 6554
rect 11282 6502 11292 6554
rect 11316 6502 11346 6554
rect 11346 6502 11358 6554
rect 11358 6502 11372 6554
rect 11396 6502 11410 6554
rect 11410 6502 11422 6554
rect 11422 6502 11452 6554
rect 11476 6502 11486 6554
rect 11486 6502 11532 6554
rect 11236 6500 11292 6502
rect 11316 6500 11372 6502
rect 11396 6500 11452 6502
rect 11476 6500 11532 6502
rect 11978 8200 12034 8256
rect 11886 6024 11942 6080
rect 11886 5888 11942 5944
rect 11236 5466 11292 5468
rect 11316 5466 11372 5468
rect 11396 5466 11452 5468
rect 11476 5466 11532 5468
rect 11236 5414 11282 5466
rect 11282 5414 11292 5466
rect 11316 5414 11346 5466
rect 11346 5414 11358 5466
rect 11358 5414 11372 5466
rect 11396 5414 11410 5466
rect 11410 5414 11422 5466
rect 11422 5414 11452 5466
rect 11476 5414 11486 5466
rect 11486 5414 11532 5466
rect 11236 5412 11292 5414
rect 11316 5412 11372 5414
rect 11396 5412 11452 5414
rect 11476 5412 11532 5414
rect 11236 4378 11292 4380
rect 11316 4378 11372 4380
rect 11396 4378 11452 4380
rect 11476 4378 11532 4380
rect 11236 4326 11282 4378
rect 11282 4326 11292 4378
rect 11316 4326 11346 4378
rect 11346 4326 11358 4378
rect 11358 4326 11372 4378
rect 11396 4326 11410 4378
rect 11410 4326 11422 4378
rect 11422 4326 11452 4378
rect 11476 4326 11486 4378
rect 11486 4326 11532 4378
rect 11236 4324 11292 4326
rect 11316 4324 11372 4326
rect 11396 4324 11452 4326
rect 11476 4324 11532 4326
rect 12254 9424 12310 9480
rect 12438 10240 12494 10296
rect 12530 9696 12586 9752
rect 12950 10362 13006 10364
rect 13030 10362 13086 10364
rect 13110 10362 13166 10364
rect 13190 10362 13246 10364
rect 12950 10310 12996 10362
rect 12996 10310 13006 10362
rect 13030 10310 13060 10362
rect 13060 10310 13072 10362
rect 13072 10310 13086 10362
rect 13110 10310 13124 10362
rect 13124 10310 13136 10362
rect 13136 10310 13166 10362
rect 13190 10310 13200 10362
rect 13200 10310 13246 10362
rect 12950 10308 13006 10310
rect 13030 10308 13086 10310
rect 13110 10308 13166 10310
rect 13190 10308 13246 10310
rect 14370 20168 14426 20224
rect 14370 19080 14426 19136
rect 14462 18808 14518 18864
rect 14094 17176 14150 17232
rect 14002 13640 14058 13696
rect 13910 13368 13966 13424
rect 13910 12688 13966 12744
rect 12714 10104 12770 10160
rect 12714 9596 12716 9616
rect 12716 9596 12768 9616
rect 12768 9596 12770 9616
rect 12714 9560 12770 9596
rect 12622 9152 12678 9208
rect 12438 8744 12494 8800
rect 12162 6432 12218 6488
rect 12070 5092 12126 5128
rect 12070 5072 12072 5092
rect 12072 5072 12124 5092
rect 12124 5072 12126 5092
rect 9523 3834 9579 3836
rect 9603 3834 9659 3836
rect 9683 3834 9739 3836
rect 9763 3834 9819 3836
rect 9523 3782 9569 3834
rect 9569 3782 9579 3834
rect 9603 3782 9633 3834
rect 9633 3782 9645 3834
rect 9645 3782 9659 3834
rect 9683 3782 9697 3834
rect 9697 3782 9709 3834
rect 9709 3782 9739 3834
rect 9763 3782 9773 3834
rect 9773 3782 9819 3834
rect 9523 3780 9579 3782
rect 9603 3780 9659 3782
rect 9683 3780 9739 3782
rect 9763 3780 9819 3782
rect 11236 3290 11292 3292
rect 11316 3290 11372 3292
rect 11396 3290 11452 3292
rect 11476 3290 11532 3292
rect 11236 3238 11282 3290
rect 11282 3238 11292 3290
rect 11316 3238 11346 3290
rect 11346 3238 11358 3290
rect 11358 3238 11372 3290
rect 11396 3238 11410 3290
rect 11410 3238 11422 3290
rect 11422 3238 11452 3290
rect 11476 3238 11486 3290
rect 11486 3238 11532 3290
rect 11236 3236 11292 3238
rect 11316 3236 11372 3238
rect 11396 3236 11452 3238
rect 11476 3236 11532 3238
rect 9523 2746 9579 2748
rect 9603 2746 9659 2748
rect 9683 2746 9739 2748
rect 9763 2746 9819 2748
rect 9523 2694 9569 2746
rect 9569 2694 9579 2746
rect 9603 2694 9633 2746
rect 9633 2694 9645 2746
rect 9645 2694 9659 2746
rect 9683 2694 9697 2746
rect 9697 2694 9709 2746
rect 9709 2694 9739 2746
rect 9763 2694 9773 2746
rect 9773 2694 9819 2746
rect 9523 2692 9579 2694
rect 9603 2692 9659 2694
rect 9683 2692 9739 2694
rect 9763 2692 9819 2694
rect 10874 2624 10930 2680
rect 11236 2202 11292 2204
rect 11316 2202 11372 2204
rect 11396 2202 11452 2204
rect 11476 2202 11532 2204
rect 11236 2150 11282 2202
rect 11282 2150 11292 2202
rect 11316 2150 11346 2202
rect 11346 2150 11358 2202
rect 11358 2150 11372 2202
rect 11396 2150 11410 2202
rect 11410 2150 11422 2202
rect 11422 2150 11452 2202
rect 11476 2150 11486 2202
rect 11486 2150 11532 2202
rect 11236 2148 11292 2150
rect 11316 2148 11372 2150
rect 11396 2148 11452 2150
rect 11476 2148 11532 2150
rect 12530 8608 12586 8664
rect 13266 9424 13322 9480
rect 12950 9274 13006 9276
rect 13030 9274 13086 9276
rect 13110 9274 13166 9276
rect 13190 9274 13246 9276
rect 12950 9222 12996 9274
rect 12996 9222 13006 9274
rect 13030 9222 13060 9274
rect 13060 9222 13072 9274
rect 13072 9222 13086 9274
rect 13110 9222 13124 9274
rect 13124 9222 13136 9274
rect 13136 9222 13166 9274
rect 13190 9222 13200 9274
rect 13200 9222 13246 9274
rect 12950 9220 13006 9222
rect 13030 9220 13086 9222
rect 13110 9220 13166 9222
rect 13190 9220 13246 9222
rect 13450 9968 13506 10024
rect 12990 8472 13046 8528
rect 12950 8186 13006 8188
rect 13030 8186 13086 8188
rect 13110 8186 13166 8188
rect 13190 8186 13246 8188
rect 12950 8134 12996 8186
rect 12996 8134 13006 8186
rect 13030 8134 13060 8186
rect 13060 8134 13072 8186
rect 13072 8134 13086 8186
rect 13110 8134 13124 8186
rect 13124 8134 13136 8186
rect 13136 8134 13166 8186
rect 13190 8134 13200 8186
rect 13200 8134 13246 8186
rect 12950 8132 13006 8134
rect 13030 8132 13086 8134
rect 13110 8132 13166 8134
rect 13190 8132 13246 8134
rect 12898 7792 12954 7848
rect 13358 8916 13360 8936
rect 13360 8916 13412 8936
rect 13412 8916 13414 8936
rect 13358 8880 13414 8916
rect 13358 7928 13414 7984
rect 12950 7098 13006 7100
rect 13030 7098 13086 7100
rect 13110 7098 13166 7100
rect 13190 7098 13246 7100
rect 12950 7046 12996 7098
rect 12996 7046 13006 7098
rect 13030 7046 13060 7098
rect 13060 7046 13072 7098
rect 13072 7046 13086 7098
rect 13110 7046 13124 7098
rect 13124 7046 13136 7098
rect 13136 7046 13166 7098
rect 13190 7046 13200 7098
rect 13200 7046 13246 7098
rect 12950 7044 13006 7046
rect 13030 7044 13086 7046
rect 13110 7044 13166 7046
rect 13190 7044 13246 7046
rect 12898 6840 12954 6896
rect 12990 6432 13046 6488
rect 12714 6024 12770 6080
rect 12950 6010 13006 6012
rect 13030 6010 13086 6012
rect 13110 6010 13166 6012
rect 13190 6010 13246 6012
rect 12950 5958 12996 6010
rect 12996 5958 13006 6010
rect 13030 5958 13060 6010
rect 13060 5958 13072 6010
rect 13072 5958 13086 6010
rect 13110 5958 13124 6010
rect 13124 5958 13136 6010
rect 13136 5958 13166 6010
rect 13190 5958 13200 6010
rect 13200 5958 13246 6010
rect 12950 5956 13006 5958
rect 13030 5956 13086 5958
rect 13110 5956 13166 5958
rect 13190 5956 13246 5958
rect 12622 5616 12678 5672
rect 12950 4922 13006 4924
rect 13030 4922 13086 4924
rect 13110 4922 13166 4924
rect 13190 4922 13246 4924
rect 12950 4870 12996 4922
rect 12996 4870 13006 4922
rect 13030 4870 13060 4922
rect 13060 4870 13072 4922
rect 13072 4870 13086 4922
rect 13110 4870 13124 4922
rect 13124 4870 13136 4922
rect 13136 4870 13166 4922
rect 13190 4870 13200 4922
rect 13200 4870 13246 4922
rect 12950 4868 13006 4870
rect 13030 4868 13086 4870
rect 13110 4868 13166 4870
rect 13190 4868 13246 4870
rect 9523 1658 9579 1660
rect 9603 1658 9659 1660
rect 9683 1658 9739 1660
rect 9763 1658 9819 1660
rect 9523 1606 9569 1658
rect 9569 1606 9579 1658
rect 9603 1606 9633 1658
rect 9633 1606 9645 1658
rect 9645 1606 9659 1658
rect 9683 1606 9697 1658
rect 9697 1606 9709 1658
rect 9709 1606 9739 1658
rect 9763 1606 9773 1658
rect 9773 1606 9819 1658
rect 9523 1604 9579 1606
rect 9603 1604 9659 1606
rect 9683 1604 9739 1606
rect 9763 1604 9819 1606
rect 11702 1808 11758 1864
rect 11236 1114 11292 1116
rect 11316 1114 11372 1116
rect 11396 1114 11452 1116
rect 11476 1114 11532 1116
rect 11236 1062 11282 1114
rect 11282 1062 11292 1114
rect 11316 1062 11346 1114
rect 11346 1062 11358 1114
rect 11358 1062 11372 1114
rect 11396 1062 11410 1114
rect 11410 1062 11422 1114
rect 11422 1062 11452 1114
rect 11476 1062 11486 1114
rect 11486 1062 11532 1114
rect 11236 1060 11292 1062
rect 11316 1060 11372 1062
rect 11396 1060 11452 1062
rect 11476 1060 11532 1062
rect 12950 3834 13006 3836
rect 13030 3834 13086 3836
rect 13110 3834 13166 3836
rect 13190 3834 13246 3836
rect 12950 3782 12996 3834
rect 12996 3782 13006 3834
rect 13030 3782 13060 3834
rect 13060 3782 13072 3834
rect 13072 3782 13086 3834
rect 13110 3782 13124 3834
rect 13124 3782 13136 3834
rect 13136 3782 13166 3834
rect 13190 3782 13200 3834
rect 13200 3782 13246 3834
rect 12950 3780 13006 3782
rect 13030 3780 13086 3782
rect 13110 3780 13166 3782
rect 13190 3780 13246 3782
rect 14002 12416 14058 12472
rect 14278 17176 14334 17232
rect 14278 16632 14334 16688
rect 14278 15000 14334 15056
rect 14186 14456 14242 14512
rect 14278 13776 14334 13832
rect 14186 13504 14242 13560
rect 14186 12960 14242 13016
rect 13726 10104 13782 10160
rect 13910 9832 13966 9888
rect 13818 9424 13874 9480
rect 13910 8472 13966 8528
rect 13726 8200 13782 8256
rect 13634 6840 13690 6896
rect 13542 6296 13598 6352
rect 13726 6296 13782 6352
rect 14094 11736 14150 11792
rect 14278 11464 14334 11520
rect 14186 10684 14188 10704
rect 14188 10684 14240 10704
rect 14240 10684 14242 10704
rect 14186 10648 14242 10684
rect 14094 10512 14150 10568
rect 14462 9288 14518 9344
rect 14370 9036 14426 9072
rect 14370 9016 14372 9036
rect 14372 9016 14424 9036
rect 14424 9016 14426 9036
rect 14278 8200 14334 8256
rect 14278 7928 14334 7984
rect 14663 28314 14719 28316
rect 14743 28314 14799 28316
rect 14823 28314 14879 28316
rect 14903 28314 14959 28316
rect 14663 28262 14709 28314
rect 14709 28262 14719 28314
rect 14743 28262 14773 28314
rect 14773 28262 14785 28314
rect 14785 28262 14799 28314
rect 14823 28262 14837 28314
rect 14837 28262 14849 28314
rect 14849 28262 14879 28314
rect 14903 28262 14913 28314
rect 14913 28262 14959 28314
rect 14663 28260 14719 28262
rect 14743 28260 14799 28262
rect 14823 28260 14879 28262
rect 14903 28260 14959 28262
rect 14663 27226 14719 27228
rect 14743 27226 14799 27228
rect 14823 27226 14879 27228
rect 14903 27226 14959 27228
rect 14663 27174 14709 27226
rect 14709 27174 14719 27226
rect 14743 27174 14773 27226
rect 14773 27174 14785 27226
rect 14785 27174 14799 27226
rect 14823 27174 14837 27226
rect 14837 27174 14849 27226
rect 14849 27174 14879 27226
rect 14903 27174 14913 27226
rect 14913 27174 14959 27226
rect 14663 27172 14719 27174
rect 14743 27172 14799 27174
rect 14823 27172 14879 27174
rect 14903 27172 14959 27174
rect 14922 26424 14978 26480
rect 14663 26138 14719 26140
rect 14743 26138 14799 26140
rect 14823 26138 14879 26140
rect 14903 26138 14959 26140
rect 14663 26086 14709 26138
rect 14709 26086 14719 26138
rect 14743 26086 14773 26138
rect 14773 26086 14785 26138
rect 14785 26086 14799 26138
rect 14823 26086 14837 26138
rect 14837 26086 14849 26138
rect 14849 26086 14879 26138
rect 14903 26086 14913 26138
rect 14913 26086 14959 26138
rect 14663 26084 14719 26086
rect 14743 26084 14799 26086
rect 14823 26084 14879 26086
rect 14903 26084 14959 26086
rect 14663 25050 14719 25052
rect 14743 25050 14799 25052
rect 14823 25050 14879 25052
rect 14903 25050 14959 25052
rect 14663 24998 14709 25050
rect 14709 24998 14719 25050
rect 14743 24998 14773 25050
rect 14773 24998 14785 25050
rect 14785 24998 14799 25050
rect 14823 24998 14837 25050
rect 14837 24998 14849 25050
rect 14849 24998 14879 25050
rect 14903 24998 14913 25050
rect 14913 24998 14959 25050
rect 14663 24996 14719 24998
rect 14743 24996 14799 24998
rect 14823 24996 14879 24998
rect 14903 24996 14959 24998
rect 14663 23962 14719 23964
rect 14743 23962 14799 23964
rect 14823 23962 14879 23964
rect 14903 23962 14959 23964
rect 14663 23910 14709 23962
rect 14709 23910 14719 23962
rect 14743 23910 14773 23962
rect 14773 23910 14785 23962
rect 14785 23910 14799 23962
rect 14823 23910 14837 23962
rect 14837 23910 14849 23962
rect 14849 23910 14879 23962
rect 14903 23910 14913 23962
rect 14913 23910 14959 23962
rect 14663 23908 14719 23910
rect 14743 23908 14799 23910
rect 14823 23908 14879 23910
rect 14903 23908 14959 23910
rect 14663 22874 14719 22876
rect 14743 22874 14799 22876
rect 14823 22874 14879 22876
rect 14903 22874 14959 22876
rect 14663 22822 14709 22874
rect 14709 22822 14719 22874
rect 14743 22822 14773 22874
rect 14773 22822 14785 22874
rect 14785 22822 14799 22874
rect 14823 22822 14837 22874
rect 14837 22822 14849 22874
rect 14849 22822 14879 22874
rect 14903 22822 14913 22874
rect 14913 22822 14959 22874
rect 14663 22820 14719 22822
rect 14743 22820 14799 22822
rect 14823 22820 14879 22822
rect 14903 22820 14959 22822
rect 14922 22380 14924 22400
rect 14924 22380 14976 22400
rect 14976 22380 14978 22400
rect 14922 22344 14978 22380
rect 14663 21786 14719 21788
rect 14743 21786 14799 21788
rect 14823 21786 14879 21788
rect 14903 21786 14959 21788
rect 14663 21734 14709 21786
rect 14709 21734 14719 21786
rect 14743 21734 14773 21786
rect 14773 21734 14785 21786
rect 14785 21734 14799 21786
rect 14823 21734 14837 21786
rect 14837 21734 14849 21786
rect 14849 21734 14879 21786
rect 14903 21734 14913 21786
rect 14913 21734 14959 21786
rect 14663 21732 14719 21734
rect 14743 21732 14799 21734
rect 14823 21732 14879 21734
rect 14903 21732 14959 21734
rect 14663 20698 14719 20700
rect 14743 20698 14799 20700
rect 14823 20698 14879 20700
rect 14903 20698 14959 20700
rect 14663 20646 14709 20698
rect 14709 20646 14719 20698
rect 14743 20646 14773 20698
rect 14773 20646 14785 20698
rect 14785 20646 14799 20698
rect 14823 20646 14837 20698
rect 14837 20646 14849 20698
rect 14849 20646 14879 20698
rect 14903 20646 14913 20698
rect 14913 20646 14959 20698
rect 14663 20644 14719 20646
rect 14743 20644 14799 20646
rect 14823 20644 14879 20646
rect 14903 20644 14959 20646
rect 14646 19780 14702 19816
rect 14646 19760 14648 19780
rect 14648 19760 14700 19780
rect 14700 19760 14702 19780
rect 14663 19610 14719 19612
rect 14743 19610 14799 19612
rect 14823 19610 14879 19612
rect 14903 19610 14959 19612
rect 14663 19558 14709 19610
rect 14709 19558 14719 19610
rect 14743 19558 14773 19610
rect 14773 19558 14785 19610
rect 14785 19558 14799 19610
rect 14823 19558 14837 19610
rect 14837 19558 14849 19610
rect 14849 19558 14879 19610
rect 14903 19558 14913 19610
rect 14913 19558 14959 19610
rect 14663 19556 14719 19558
rect 14743 19556 14799 19558
rect 14823 19556 14879 19558
rect 14903 19556 14959 19558
rect 14663 18522 14719 18524
rect 14743 18522 14799 18524
rect 14823 18522 14879 18524
rect 14903 18522 14959 18524
rect 14663 18470 14709 18522
rect 14709 18470 14719 18522
rect 14743 18470 14773 18522
rect 14773 18470 14785 18522
rect 14785 18470 14799 18522
rect 14823 18470 14837 18522
rect 14837 18470 14849 18522
rect 14849 18470 14879 18522
rect 14903 18470 14913 18522
rect 14913 18470 14959 18522
rect 14663 18468 14719 18470
rect 14743 18468 14799 18470
rect 14823 18468 14879 18470
rect 14903 18468 14959 18470
rect 14663 17434 14719 17436
rect 14743 17434 14799 17436
rect 14823 17434 14879 17436
rect 14903 17434 14959 17436
rect 14663 17382 14709 17434
rect 14709 17382 14719 17434
rect 14743 17382 14773 17434
rect 14773 17382 14785 17434
rect 14785 17382 14799 17434
rect 14823 17382 14837 17434
rect 14837 17382 14849 17434
rect 14849 17382 14879 17434
rect 14903 17382 14913 17434
rect 14913 17382 14959 17434
rect 14663 17380 14719 17382
rect 14743 17380 14799 17382
rect 14823 17380 14879 17382
rect 14903 17380 14959 17382
rect 14663 16346 14719 16348
rect 14743 16346 14799 16348
rect 14823 16346 14879 16348
rect 14903 16346 14959 16348
rect 14663 16294 14709 16346
rect 14709 16294 14719 16346
rect 14743 16294 14773 16346
rect 14773 16294 14785 16346
rect 14785 16294 14799 16346
rect 14823 16294 14837 16346
rect 14837 16294 14849 16346
rect 14849 16294 14879 16346
rect 14903 16294 14913 16346
rect 14913 16294 14959 16346
rect 14663 16292 14719 16294
rect 14743 16292 14799 16294
rect 14823 16292 14879 16294
rect 14903 16292 14959 16294
rect 14830 15544 14886 15600
rect 14663 15258 14719 15260
rect 14743 15258 14799 15260
rect 14823 15258 14879 15260
rect 14903 15258 14959 15260
rect 14663 15206 14709 15258
rect 14709 15206 14719 15258
rect 14743 15206 14773 15258
rect 14773 15206 14785 15258
rect 14785 15206 14799 15258
rect 14823 15206 14837 15258
rect 14837 15206 14849 15258
rect 14849 15206 14879 15258
rect 14903 15206 14913 15258
rect 14913 15206 14959 15258
rect 14663 15204 14719 15206
rect 14743 15204 14799 15206
rect 14823 15204 14879 15206
rect 14903 15204 14959 15206
rect 14830 14728 14886 14784
rect 14663 14170 14719 14172
rect 14743 14170 14799 14172
rect 14823 14170 14879 14172
rect 14903 14170 14959 14172
rect 14663 14118 14709 14170
rect 14709 14118 14719 14170
rect 14743 14118 14773 14170
rect 14773 14118 14785 14170
rect 14785 14118 14799 14170
rect 14823 14118 14837 14170
rect 14837 14118 14849 14170
rect 14849 14118 14879 14170
rect 14903 14118 14913 14170
rect 14913 14118 14959 14170
rect 14663 14116 14719 14118
rect 14743 14116 14799 14118
rect 14823 14116 14879 14118
rect 14903 14116 14959 14118
rect 14663 13082 14719 13084
rect 14743 13082 14799 13084
rect 14823 13082 14879 13084
rect 14903 13082 14959 13084
rect 14663 13030 14709 13082
rect 14709 13030 14719 13082
rect 14743 13030 14773 13082
rect 14773 13030 14785 13082
rect 14785 13030 14799 13082
rect 14823 13030 14837 13082
rect 14837 13030 14849 13082
rect 14849 13030 14879 13082
rect 14903 13030 14913 13082
rect 14913 13030 14959 13082
rect 14663 13028 14719 13030
rect 14743 13028 14799 13030
rect 14823 13028 14879 13030
rect 14903 13028 14959 13030
rect 14663 11994 14719 11996
rect 14743 11994 14799 11996
rect 14823 11994 14879 11996
rect 14903 11994 14959 11996
rect 14663 11942 14709 11994
rect 14709 11942 14719 11994
rect 14743 11942 14773 11994
rect 14773 11942 14785 11994
rect 14785 11942 14799 11994
rect 14823 11942 14837 11994
rect 14837 11942 14849 11994
rect 14849 11942 14879 11994
rect 14903 11942 14913 11994
rect 14913 11942 14959 11994
rect 14663 11940 14719 11942
rect 14743 11940 14799 11942
rect 14823 11940 14879 11942
rect 14903 11940 14959 11942
rect 14663 10906 14719 10908
rect 14743 10906 14799 10908
rect 14823 10906 14879 10908
rect 14903 10906 14959 10908
rect 14663 10854 14709 10906
rect 14709 10854 14719 10906
rect 14743 10854 14773 10906
rect 14773 10854 14785 10906
rect 14785 10854 14799 10906
rect 14823 10854 14837 10906
rect 14837 10854 14849 10906
rect 14849 10854 14879 10906
rect 14903 10854 14913 10906
rect 14913 10854 14959 10906
rect 14663 10852 14719 10854
rect 14743 10852 14799 10854
rect 14823 10852 14879 10854
rect 14903 10852 14959 10854
rect 14646 10376 14702 10432
rect 14663 9818 14719 9820
rect 14743 9818 14799 9820
rect 14823 9818 14879 9820
rect 14903 9818 14959 9820
rect 14663 9766 14709 9818
rect 14709 9766 14719 9818
rect 14743 9766 14773 9818
rect 14773 9766 14785 9818
rect 14785 9766 14799 9818
rect 14823 9766 14837 9818
rect 14837 9766 14849 9818
rect 14849 9766 14879 9818
rect 14903 9766 14913 9818
rect 14913 9766 14959 9818
rect 14663 9764 14719 9766
rect 14743 9764 14799 9766
rect 14823 9764 14879 9766
rect 14903 9764 14959 9766
rect 14663 8730 14719 8732
rect 14743 8730 14799 8732
rect 14823 8730 14879 8732
rect 14903 8730 14959 8732
rect 14663 8678 14709 8730
rect 14709 8678 14719 8730
rect 14743 8678 14773 8730
rect 14773 8678 14785 8730
rect 14785 8678 14799 8730
rect 14823 8678 14837 8730
rect 14837 8678 14849 8730
rect 14849 8678 14879 8730
rect 14903 8678 14913 8730
rect 14913 8678 14959 8730
rect 14663 8676 14719 8678
rect 14743 8676 14799 8678
rect 14823 8676 14879 8678
rect 14903 8676 14959 8678
rect 14186 7828 14188 7848
rect 14188 7828 14240 7848
rect 14240 7828 14242 7848
rect 14186 7792 14242 7828
rect 14278 7112 14334 7168
rect 13910 6704 13966 6760
rect 13910 5480 13966 5536
rect 14663 7642 14719 7644
rect 14743 7642 14799 7644
rect 14823 7642 14879 7644
rect 14903 7642 14959 7644
rect 14663 7590 14709 7642
rect 14709 7590 14719 7642
rect 14743 7590 14773 7642
rect 14773 7590 14785 7642
rect 14785 7590 14799 7642
rect 14823 7590 14837 7642
rect 14837 7590 14849 7642
rect 14849 7590 14879 7642
rect 14903 7590 14913 7642
rect 14913 7590 14959 7642
rect 14663 7588 14719 7590
rect 14743 7588 14799 7590
rect 14823 7588 14879 7590
rect 14903 7588 14959 7590
rect 14554 7384 14610 7440
rect 14663 6554 14719 6556
rect 14743 6554 14799 6556
rect 14823 6554 14879 6556
rect 14903 6554 14959 6556
rect 14663 6502 14709 6554
rect 14709 6502 14719 6554
rect 14743 6502 14773 6554
rect 14773 6502 14785 6554
rect 14785 6502 14799 6554
rect 14823 6502 14837 6554
rect 14837 6502 14849 6554
rect 14849 6502 14879 6554
rect 14903 6502 14913 6554
rect 14913 6502 14959 6554
rect 14663 6500 14719 6502
rect 14743 6500 14799 6502
rect 14823 6500 14879 6502
rect 14903 6500 14959 6502
rect 14370 6160 14426 6216
rect 14830 5752 14886 5808
rect 14278 5480 14334 5536
rect 14663 5466 14719 5468
rect 14743 5466 14799 5468
rect 14823 5466 14879 5468
rect 14903 5466 14959 5468
rect 14663 5414 14709 5466
rect 14709 5414 14719 5466
rect 14743 5414 14773 5466
rect 14773 5414 14785 5466
rect 14785 5414 14799 5466
rect 14823 5414 14837 5466
rect 14837 5414 14849 5466
rect 14849 5414 14879 5466
rect 14903 5414 14913 5466
rect 14913 5414 14959 5466
rect 14663 5412 14719 5414
rect 14743 5412 14799 5414
rect 14823 5412 14879 5414
rect 14903 5412 14959 5414
rect 14002 5228 14058 5264
rect 14002 5208 14004 5228
rect 14004 5208 14056 5228
rect 14056 5208 14058 5228
rect 14278 4936 14334 4992
rect 14663 4378 14719 4380
rect 14743 4378 14799 4380
rect 14823 4378 14879 4380
rect 14903 4378 14959 4380
rect 14663 4326 14709 4378
rect 14709 4326 14719 4378
rect 14743 4326 14773 4378
rect 14773 4326 14785 4378
rect 14785 4326 14799 4378
rect 14823 4326 14837 4378
rect 14837 4326 14849 4378
rect 14849 4326 14879 4378
rect 14903 4326 14913 4378
rect 14913 4326 14959 4378
rect 14663 4324 14719 4326
rect 14743 4324 14799 4326
rect 14823 4324 14879 4326
rect 14903 4324 14959 4326
rect 14370 3984 14426 4040
rect 14663 3290 14719 3292
rect 14743 3290 14799 3292
rect 14823 3290 14879 3292
rect 14903 3290 14959 3292
rect 14663 3238 14709 3290
rect 14709 3238 14719 3290
rect 14743 3238 14773 3290
rect 14773 3238 14785 3290
rect 14785 3238 14799 3290
rect 14823 3238 14837 3290
rect 14837 3238 14849 3290
rect 14849 3238 14879 3290
rect 14903 3238 14913 3290
rect 14913 3238 14959 3290
rect 14663 3236 14719 3238
rect 14743 3236 14799 3238
rect 14823 3236 14879 3238
rect 14903 3236 14959 3238
rect 12950 2746 13006 2748
rect 13030 2746 13086 2748
rect 13110 2746 13166 2748
rect 13190 2746 13246 2748
rect 12950 2694 12996 2746
rect 12996 2694 13006 2746
rect 13030 2694 13060 2746
rect 13060 2694 13072 2746
rect 13072 2694 13086 2746
rect 13110 2694 13124 2746
rect 13124 2694 13136 2746
rect 13136 2694 13166 2746
rect 13190 2694 13200 2746
rect 13200 2694 13246 2746
rect 12950 2692 13006 2694
rect 13030 2692 13086 2694
rect 13110 2692 13166 2694
rect 13190 2692 13246 2694
rect 14663 2202 14719 2204
rect 14743 2202 14799 2204
rect 14823 2202 14879 2204
rect 14903 2202 14959 2204
rect 14663 2150 14709 2202
rect 14709 2150 14719 2202
rect 14743 2150 14773 2202
rect 14773 2150 14785 2202
rect 14785 2150 14799 2202
rect 14823 2150 14837 2202
rect 14837 2150 14849 2202
rect 14849 2150 14879 2202
rect 14903 2150 14913 2202
rect 14913 2150 14959 2202
rect 14663 2148 14719 2150
rect 14743 2148 14799 2150
rect 14823 2148 14879 2150
rect 14903 2148 14959 2150
rect 15106 35980 15108 36000
rect 15108 35980 15160 36000
rect 15160 35980 15162 36000
rect 15106 35944 15162 35980
rect 15106 34856 15162 34912
rect 15106 31592 15162 31648
rect 15106 30540 15108 30560
rect 15108 30540 15160 30560
rect 15160 30540 15162 30560
rect 15106 30504 15162 30540
rect 15106 24792 15162 24848
rect 15106 23976 15162 24032
rect 15106 22924 15108 22944
rect 15108 22924 15160 22944
rect 15160 22924 15162 22944
rect 15106 22888 15162 22924
rect 15290 35536 15346 35592
rect 15290 29688 15346 29744
rect 15290 25608 15346 25664
rect 15106 21800 15162 21856
rect 15106 18536 15162 18592
rect 15382 21936 15438 21992
rect 15290 20712 15346 20768
rect 15198 18128 15254 18184
rect 15198 16496 15254 16552
rect 15106 16360 15162 16416
rect 15106 14184 15162 14240
rect 15290 14320 15346 14376
rect 15198 13096 15254 13152
rect 15106 11872 15162 11928
rect 15198 10920 15254 10976
rect 15106 9832 15162 9888
rect 15106 8744 15162 8800
rect 15106 6840 15162 6896
rect 15198 6160 15254 6216
rect 15106 5480 15162 5536
rect 12950 1658 13006 1660
rect 13030 1658 13086 1660
rect 13110 1658 13166 1660
rect 13190 1658 13246 1660
rect 12950 1606 12996 1658
rect 12996 1606 13006 1658
rect 13030 1606 13060 1658
rect 13060 1606 13072 1658
rect 13072 1606 13086 1658
rect 13110 1606 13124 1658
rect 13124 1606 13136 1658
rect 13136 1606 13166 1658
rect 13190 1606 13200 1658
rect 13200 1606 13246 1658
rect 12950 1604 13006 1606
rect 13030 1604 13086 1606
rect 13110 1604 13166 1606
rect 13190 1604 13246 1606
rect 15658 22208 15714 22264
rect 15566 19896 15622 19952
rect 14663 1114 14719 1116
rect 14743 1114 14799 1116
rect 14823 1114 14879 1116
rect 14903 1114 14959 1116
rect 14663 1062 14709 1114
rect 14709 1062 14719 1114
rect 14743 1062 14773 1114
rect 14773 1062 14785 1114
rect 14785 1062 14799 1114
rect 14823 1062 14837 1114
rect 14837 1062 14849 1114
rect 14849 1062 14879 1114
rect 14903 1062 14913 1114
rect 14913 1062 14959 1114
rect 14663 1060 14719 1062
rect 14743 1060 14799 1062
rect 14823 1060 14879 1062
rect 14903 1060 14959 1062
<< metal3 >>
rect 4372 43552 4688 43553
rect 4372 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4688 43552
rect 4372 43487 4688 43488
rect 7799 43552 8115 43553
rect 7799 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8115 43552
rect 7799 43487 8115 43488
rect 11226 43552 11542 43553
rect 11226 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11542 43552
rect 11226 43487 11542 43488
rect 14653 43552 14969 43553
rect 14653 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14969 43552
rect 14653 43487 14969 43488
rect 2659 43008 2975 43009
rect 2659 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2975 43008
rect 2659 42943 2975 42944
rect 6086 43008 6402 43009
rect 6086 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6402 43008
rect 6086 42943 6402 42944
rect 9513 43008 9829 43009
rect 9513 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9829 43008
rect 9513 42943 9829 42944
rect 12940 43008 13256 43009
rect 12940 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13256 43008
rect 12940 42943 13256 42944
rect 4372 42464 4688 42465
rect 4372 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4688 42464
rect 4372 42399 4688 42400
rect 7799 42464 8115 42465
rect 7799 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8115 42464
rect 7799 42399 8115 42400
rect 11226 42464 11542 42465
rect 11226 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11542 42464
rect 11226 42399 11542 42400
rect 14653 42464 14969 42465
rect 14653 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14969 42464
rect 14653 42399 14969 42400
rect 5390 42060 5396 42124
rect 5460 42122 5466 42124
rect 11697 42122 11763 42125
rect 5460 42120 11763 42122
rect 5460 42064 11702 42120
rect 11758 42064 11763 42120
rect 5460 42062 11763 42064
rect 5460 42060 5466 42062
rect 11697 42059 11763 42062
rect 2659 41920 2975 41921
rect 2659 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2975 41920
rect 2659 41855 2975 41856
rect 6086 41920 6402 41921
rect 6086 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6402 41920
rect 6086 41855 6402 41856
rect 9513 41920 9829 41921
rect 9513 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9829 41920
rect 9513 41855 9829 41856
rect 12940 41920 13256 41921
rect 12940 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13256 41920
rect 12940 41855 13256 41856
rect 5717 41852 5783 41853
rect 5717 41848 5764 41852
rect 5828 41850 5834 41852
rect 6545 41850 6611 41853
rect 6678 41850 6684 41852
rect 5717 41792 5722 41848
rect 5717 41788 5764 41792
rect 5828 41790 5874 41850
rect 6545 41848 6684 41850
rect 6545 41792 6550 41848
rect 6606 41792 6684 41848
rect 6545 41790 6684 41792
rect 5828 41788 5834 41790
rect 5717 41787 5783 41788
rect 6545 41787 6611 41790
rect 6678 41788 6684 41790
rect 6748 41788 6754 41852
rect 7414 41788 7420 41852
rect 7484 41850 7490 41852
rect 8109 41850 8175 41853
rect 10961 41852 11027 41853
rect 10910 41850 10916 41852
rect 7484 41848 8175 41850
rect 7484 41792 8114 41848
rect 8170 41792 8175 41848
rect 7484 41790 8175 41792
rect 10870 41790 10916 41850
rect 10980 41848 11027 41852
rect 11022 41792 11027 41848
rect 7484 41788 7490 41790
rect 8109 41787 8175 41790
rect 10910 41788 10916 41790
rect 10980 41788 11027 41792
rect 10961 41787 11027 41788
rect 3918 41516 3924 41580
rect 3988 41578 3994 41580
rect 7281 41578 7347 41581
rect 3988 41576 7347 41578
rect 3988 41520 7286 41576
rect 7342 41520 7347 41576
rect 3988 41518 7347 41520
rect 3988 41516 3994 41518
rect 7281 41515 7347 41518
rect 10726 41516 10732 41580
rect 10796 41578 10802 41580
rect 12433 41578 12499 41581
rect 10796 41576 12499 41578
rect 10796 41520 12438 41576
rect 12494 41520 12499 41576
rect 10796 41518 12499 41520
rect 10796 41516 10802 41518
rect 12433 41515 12499 41518
rect 4372 41376 4688 41377
rect 4372 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4688 41376
rect 4372 41311 4688 41312
rect 7799 41376 8115 41377
rect 7799 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8115 41376
rect 7799 41311 8115 41312
rect 11226 41376 11542 41377
rect 11226 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11542 41376
rect 11226 41311 11542 41312
rect 14653 41376 14969 41377
rect 14653 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14969 41376
rect 14653 41311 14969 41312
rect 2659 40832 2975 40833
rect 2659 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2975 40832
rect 2659 40767 2975 40768
rect 6086 40832 6402 40833
rect 6086 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6402 40832
rect 6086 40767 6402 40768
rect 9513 40832 9829 40833
rect 9513 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9829 40832
rect 9513 40767 9829 40768
rect 12940 40832 13256 40833
rect 12940 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13256 40832
rect 12940 40767 13256 40768
rect 0 40626 160 40656
rect 749 40626 815 40629
rect 0 40624 815 40626
rect 0 40568 754 40624
rect 810 40568 815 40624
rect 0 40566 815 40568
rect 0 40536 160 40566
rect 749 40563 815 40566
rect 4372 40288 4688 40289
rect 4372 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4688 40288
rect 4372 40223 4688 40224
rect 7799 40288 8115 40289
rect 7799 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8115 40288
rect 7799 40223 8115 40224
rect 11226 40288 11542 40289
rect 11226 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11542 40288
rect 11226 40223 11542 40224
rect 14653 40288 14969 40289
rect 14653 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14969 40288
rect 14653 40223 14969 40224
rect 1393 39944 1459 39949
rect 1393 39888 1398 39944
rect 1454 39888 1459 39944
rect 1393 39883 1459 39888
rect 0 39810 160 39840
rect 1396 39810 1456 39883
rect 0 39750 1456 39810
rect 0 39720 160 39750
rect 2659 39744 2975 39745
rect 2659 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2975 39744
rect 2659 39679 2975 39680
rect 6086 39744 6402 39745
rect 6086 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6402 39744
rect 6086 39679 6402 39680
rect 9513 39744 9829 39745
rect 9513 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9829 39744
rect 9513 39679 9829 39680
rect 12940 39744 13256 39745
rect 12940 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13256 39744
rect 12940 39679 13256 39680
rect 13997 39536 14063 39541
rect 13997 39480 14002 39536
rect 14058 39480 14063 39536
rect 13997 39475 14063 39480
rect 14181 39538 14247 39541
rect 15840 39538 16000 39568
rect 14181 39536 16000 39538
rect 14181 39480 14186 39536
rect 14242 39480 16000 39536
rect 14181 39478 16000 39480
rect 14181 39475 14247 39478
rect 14000 39402 14060 39475
rect 15840 39448 16000 39478
rect 14000 39342 15164 39402
rect 15104 39266 15164 39342
rect 15840 39266 16000 39296
rect 15104 39206 16000 39266
rect 4372 39200 4688 39201
rect 4372 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4688 39200
rect 4372 39135 4688 39136
rect 7799 39200 8115 39201
rect 7799 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8115 39200
rect 7799 39135 8115 39136
rect 11226 39200 11542 39201
rect 11226 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11542 39200
rect 11226 39135 11542 39136
rect 14653 39200 14969 39201
rect 14653 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14969 39200
rect 15840 39176 16000 39206
rect 14653 39135 14969 39136
rect 0 38994 160 39024
rect 749 38994 815 38997
rect 0 38992 815 38994
rect 0 38936 754 38992
rect 810 38936 815 38992
rect 0 38934 815 38936
rect 0 38904 160 38934
rect 749 38931 815 38934
rect 13905 38994 13971 38997
rect 15840 38994 16000 39024
rect 13905 38992 16000 38994
rect 13905 38936 13910 38992
rect 13966 38936 16000 38992
rect 13905 38934 16000 38936
rect 13905 38931 13971 38934
rect 15840 38904 16000 38934
rect 14365 38722 14431 38725
rect 15840 38722 16000 38752
rect 14365 38720 16000 38722
rect 14365 38664 14370 38720
rect 14426 38664 16000 38720
rect 14365 38662 16000 38664
rect 14365 38659 14431 38662
rect 2659 38656 2975 38657
rect 2659 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2975 38656
rect 2659 38591 2975 38592
rect 6086 38656 6402 38657
rect 6086 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6402 38656
rect 6086 38591 6402 38592
rect 9513 38656 9829 38657
rect 9513 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9829 38656
rect 9513 38591 9829 38592
rect 12940 38656 13256 38657
rect 12940 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13256 38656
rect 15840 38632 16000 38662
rect 12940 38591 13256 38592
rect 13629 38450 13695 38453
rect 14181 38450 14247 38453
rect 15840 38450 16000 38480
rect 13629 38448 14106 38450
rect 13629 38392 13634 38448
rect 13690 38392 14106 38448
rect 13629 38390 14106 38392
rect 13629 38387 13695 38390
rect 14046 38314 14106 38390
rect 14181 38448 16000 38450
rect 14181 38392 14186 38448
rect 14242 38392 16000 38448
rect 14181 38390 16000 38392
rect 14181 38387 14247 38390
rect 15840 38360 16000 38390
rect 14046 38254 15164 38314
rect 0 38178 160 38208
rect 749 38178 815 38181
rect 0 38176 815 38178
rect 0 38120 754 38176
rect 810 38120 815 38176
rect 0 38118 815 38120
rect 0 38088 160 38118
rect 749 38115 815 38118
rect 11789 38178 11855 38181
rect 13445 38178 13511 38181
rect 11789 38176 13511 38178
rect 11789 38120 11794 38176
rect 11850 38120 13450 38176
rect 13506 38120 13511 38176
rect 11789 38118 13511 38120
rect 15104 38178 15164 38254
rect 15840 38178 16000 38208
rect 15104 38118 16000 38178
rect 11789 38115 11855 38118
rect 13445 38115 13511 38118
rect 4372 38112 4688 38113
rect 4372 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4688 38112
rect 4372 38047 4688 38048
rect 7799 38112 8115 38113
rect 7799 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8115 38112
rect 7799 38047 8115 38048
rect 11226 38112 11542 38113
rect 11226 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11542 38112
rect 11226 38047 11542 38048
rect 14653 38112 14969 38113
rect 14653 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14969 38112
rect 15840 38088 16000 38118
rect 14653 38047 14969 38048
rect 13813 37906 13879 37909
rect 15840 37906 16000 37936
rect 13813 37904 16000 37906
rect 13813 37848 13818 37904
rect 13874 37848 16000 37904
rect 13813 37846 16000 37848
rect 13813 37843 13879 37846
rect 15840 37816 16000 37846
rect 14365 37634 14431 37637
rect 15840 37634 16000 37664
rect 14365 37632 16000 37634
rect 14365 37576 14370 37632
rect 14426 37576 16000 37632
rect 14365 37574 16000 37576
rect 14365 37571 14431 37574
rect 2659 37568 2975 37569
rect 2659 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2975 37568
rect 2659 37503 2975 37504
rect 6086 37568 6402 37569
rect 6086 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6402 37568
rect 6086 37503 6402 37504
rect 9513 37568 9829 37569
rect 9513 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9829 37568
rect 9513 37503 9829 37504
rect 12940 37568 13256 37569
rect 12940 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13256 37568
rect 15840 37544 16000 37574
rect 12940 37503 13256 37504
rect 0 37362 160 37392
rect 749 37362 815 37365
rect 0 37360 815 37362
rect 0 37304 754 37360
rect 810 37304 815 37360
rect 0 37302 815 37304
rect 0 37272 160 37302
rect 749 37299 815 37302
rect 14181 37362 14247 37365
rect 15840 37362 16000 37392
rect 14181 37360 16000 37362
rect 14181 37304 14186 37360
rect 14242 37304 16000 37360
rect 14181 37302 16000 37304
rect 14181 37299 14247 37302
rect 15840 37272 16000 37302
rect 7281 37226 7347 37229
rect 12801 37226 12867 37229
rect 7281 37224 12867 37226
rect 7281 37168 7286 37224
rect 7342 37168 12806 37224
rect 12862 37168 12867 37224
rect 7281 37166 12867 37168
rect 7281 37163 7347 37166
rect 12801 37163 12867 37166
rect 13629 37226 13695 37229
rect 13629 37224 15164 37226
rect 13629 37168 13634 37224
rect 13690 37168 15164 37224
rect 13629 37166 15164 37168
rect 13629 37163 13695 37166
rect 15104 37090 15164 37166
rect 15840 37090 16000 37120
rect 15104 37030 16000 37090
rect 4372 37024 4688 37025
rect 4372 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4688 37024
rect 4372 36959 4688 36960
rect 7799 37024 8115 37025
rect 7799 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8115 37024
rect 7799 36959 8115 36960
rect 11226 37024 11542 37025
rect 11226 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11542 37024
rect 11226 36959 11542 36960
rect 14653 37024 14969 37025
rect 14653 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14969 37024
rect 15840 37000 16000 37030
rect 14653 36959 14969 36960
rect 13629 36818 13695 36821
rect 15840 36818 16000 36848
rect 13629 36816 16000 36818
rect 13629 36760 13634 36816
rect 13690 36760 16000 36816
rect 13629 36758 16000 36760
rect 13629 36755 13695 36758
rect 15840 36728 16000 36758
rect 11329 36682 11395 36685
rect 12985 36682 13051 36685
rect 11329 36680 13051 36682
rect 11329 36624 11334 36680
rect 11390 36624 12990 36680
rect 13046 36624 13051 36680
rect 11329 36622 13051 36624
rect 11329 36619 11395 36622
rect 12985 36619 13051 36622
rect 0 36546 160 36576
rect 749 36546 815 36549
rect 0 36544 815 36546
rect 0 36488 754 36544
rect 810 36488 815 36544
rect 0 36486 815 36488
rect 0 36456 160 36486
rect 749 36483 815 36486
rect 14365 36546 14431 36549
rect 15840 36546 16000 36576
rect 14365 36544 16000 36546
rect 14365 36488 14370 36544
rect 14426 36488 16000 36544
rect 14365 36486 16000 36488
rect 14365 36483 14431 36486
rect 2659 36480 2975 36481
rect 2659 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2975 36480
rect 2659 36415 2975 36416
rect 6086 36480 6402 36481
rect 6086 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6402 36480
rect 6086 36415 6402 36416
rect 9513 36480 9829 36481
rect 9513 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9829 36480
rect 9513 36415 9829 36416
rect 12940 36480 13256 36481
rect 12940 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13256 36480
rect 15840 36456 16000 36486
rect 12940 36415 13256 36416
rect 13813 36274 13879 36277
rect 15840 36274 16000 36304
rect 13813 36272 16000 36274
rect 13813 36216 13818 36272
rect 13874 36216 16000 36272
rect 13813 36214 16000 36216
rect 13813 36211 13879 36214
rect 15840 36184 16000 36214
rect 15101 36002 15167 36005
rect 15840 36002 16000 36032
rect 15101 36000 16000 36002
rect 15101 35944 15106 36000
rect 15162 35944 16000 36000
rect 15101 35942 16000 35944
rect 15101 35939 15167 35942
rect 4372 35936 4688 35937
rect 4372 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4688 35936
rect 4372 35871 4688 35872
rect 7799 35936 8115 35937
rect 7799 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8115 35936
rect 7799 35871 8115 35872
rect 11226 35936 11542 35937
rect 11226 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11542 35936
rect 11226 35871 11542 35872
rect 14653 35936 14969 35937
rect 14653 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14969 35936
rect 15840 35912 16000 35942
rect 14653 35871 14969 35872
rect 1393 35866 1459 35869
rect 798 35864 1459 35866
rect 798 35808 1398 35864
rect 1454 35808 1459 35864
rect 798 35806 1459 35808
rect 0 35730 160 35760
rect 798 35730 858 35806
rect 1393 35803 1459 35806
rect 0 35670 858 35730
rect 13721 35730 13787 35733
rect 15840 35730 16000 35760
rect 13721 35728 16000 35730
rect 13721 35672 13726 35728
rect 13782 35672 16000 35728
rect 13721 35670 16000 35672
rect 0 35640 160 35670
rect 13721 35667 13787 35670
rect 15840 35640 16000 35670
rect 5441 35594 5507 35597
rect 13261 35594 13327 35597
rect 5441 35592 13327 35594
rect 5441 35536 5446 35592
rect 5502 35536 13266 35592
rect 13322 35536 13327 35592
rect 5441 35534 13327 35536
rect 5441 35531 5507 35534
rect 13261 35531 13327 35534
rect 15285 35594 15351 35597
rect 15285 35592 15394 35594
rect 15285 35536 15290 35592
rect 15346 35536 15394 35592
rect 15285 35531 15394 35536
rect 15334 35458 15394 35531
rect 15840 35458 16000 35488
rect 15334 35398 16000 35458
rect 2659 35392 2975 35393
rect 2659 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2975 35392
rect 2659 35327 2975 35328
rect 6086 35392 6402 35393
rect 6086 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6402 35392
rect 6086 35327 6402 35328
rect 9513 35392 9829 35393
rect 9513 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9829 35392
rect 9513 35327 9829 35328
rect 12940 35392 13256 35393
rect 12940 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13256 35392
rect 15840 35368 16000 35398
rect 12940 35327 13256 35328
rect 13813 35186 13879 35189
rect 15840 35186 16000 35216
rect 13813 35184 16000 35186
rect 13813 35128 13818 35184
rect 13874 35128 16000 35184
rect 13813 35126 16000 35128
rect 13813 35123 13879 35126
rect 15840 35096 16000 35126
rect 10961 35050 11027 35053
rect 13537 35050 13603 35053
rect 10961 35048 13603 35050
rect 10961 34992 10966 35048
rect 11022 34992 13542 35048
rect 13598 34992 13603 35048
rect 10961 34990 13603 34992
rect 10961 34987 11027 34990
rect 13537 34987 13603 34990
rect 0 34914 160 34944
rect 749 34914 815 34917
rect 0 34912 815 34914
rect 0 34856 754 34912
rect 810 34856 815 34912
rect 0 34854 815 34856
rect 0 34824 160 34854
rect 749 34851 815 34854
rect 15101 34914 15167 34917
rect 15840 34914 16000 34944
rect 15101 34912 16000 34914
rect 15101 34856 15106 34912
rect 15162 34856 16000 34912
rect 15101 34854 16000 34856
rect 15101 34851 15167 34854
rect 4372 34848 4688 34849
rect 4372 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4688 34848
rect 4372 34783 4688 34784
rect 7799 34848 8115 34849
rect 7799 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8115 34848
rect 7799 34783 8115 34784
rect 11226 34848 11542 34849
rect 11226 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11542 34848
rect 11226 34783 11542 34784
rect 14653 34848 14969 34849
rect 14653 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14969 34848
rect 15840 34824 16000 34854
rect 14653 34783 14969 34784
rect 13905 34642 13971 34645
rect 15840 34642 16000 34672
rect 13905 34640 16000 34642
rect 13905 34584 13910 34640
rect 13966 34584 16000 34640
rect 13905 34582 16000 34584
rect 13905 34579 13971 34582
rect 15840 34552 16000 34582
rect 1393 34506 1459 34509
rect 798 34504 1459 34506
rect 798 34448 1398 34504
rect 1454 34448 1459 34504
rect 798 34446 1459 34448
rect 0 34098 160 34128
rect 798 34098 858 34446
rect 1393 34443 1459 34446
rect 14365 34370 14431 34373
rect 15840 34370 16000 34400
rect 14365 34368 16000 34370
rect 14365 34312 14370 34368
rect 14426 34312 16000 34368
rect 14365 34310 16000 34312
rect 14365 34307 14431 34310
rect 2659 34304 2975 34305
rect 2659 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2975 34304
rect 2659 34239 2975 34240
rect 6086 34304 6402 34305
rect 6086 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6402 34304
rect 6086 34239 6402 34240
rect 9513 34304 9829 34305
rect 9513 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9829 34304
rect 9513 34239 9829 34240
rect 12940 34304 13256 34305
rect 12940 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13256 34304
rect 15840 34280 16000 34310
rect 12940 34239 13256 34240
rect 0 34038 858 34098
rect 13629 34098 13695 34101
rect 14181 34098 14247 34101
rect 15840 34098 16000 34128
rect 13629 34096 14106 34098
rect 13629 34040 13634 34096
rect 13690 34040 14106 34096
rect 13629 34038 14106 34040
rect 0 34008 160 34038
rect 13629 34035 13695 34038
rect 14046 33962 14106 34038
rect 14181 34096 16000 34098
rect 14181 34040 14186 34096
rect 14242 34040 16000 34096
rect 14181 34038 16000 34040
rect 14181 34035 14247 34038
rect 15840 34008 16000 34038
rect 14046 33902 15164 33962
rect 15104 33826 15164 33902
rect 15840 33826 16000 33856
rect 15104 33766 16000 33826
rect 4372 33760 4688 33761
rect 4372 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4688 33760
rect 4372 33695 4688 33696
rect 7799 33760 8115 33761
rect 7799 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8115 33760
rect 7799 33695 8115 33696
rect 11226 33760 11542 33761
rect 11226 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11542 33760
rect 11226 33695 11542 33696
rect 14653 33760 14969 33761
rect 14653 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14969 33760
rect 15840 33736 16000 33766
rect 14653 33695 14969 33696
rect 13905 33554 13971 33557
rect 15840 33554 16000 33584
rect 13905 33552 16000 33554
rect 13905 33496 13910 33552
rect 13966 33496 16000 33552
rect 13905 33494 16000 33496
rect 13905 33491 13971 33494
rect 15840 33464 16000 33494
rect 0 33282 160 33312
rect 749 33282 815 33285
rect 0 33280 815 33282
rect 0 33224 754 33280
rect 810 33224 815 33280
rect 0 33222 815 33224
rect 0 33192 160 33222
rect 749 33219 815 33222
rect 14365 33282 14431 33285
rect 15840 33282 16000 33312
rect 14365 33280 16000 33282
rect 14365 33224 14370 33280
rect 14426 33224 16000 33280
rect 14365 33222 16000 33224
rect 14365 33219 14431 33222
rect 2659 33216 2975 33217
rect 2659 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2975 33216
rect 2659 33151 2975 33152
rect 6086 33216 6402 33217
rect 6086 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6402 33216
rect 6086 33151 6402 33152
rect 9513 33216 9829 33217
rect 9513 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9829 33216
rect 9513 33151 9829 33152
rect 12940 33216 13256 33217
rect 12940 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13256 33216
rect 15840 33192 16000 33222
rect 12940 33151 13256 33152
rect 11421 33146 11487 33149
rect 12617 33146 12683 33149
rect 11421 33144 12683 33146
rect 11421 33088 11426 33144
rect 11482 33088 12622 33144
rect 12678 33088 12683 33144
rect 11421 33086 12683 33088
rect 11421 33083 11487 33086
rect 12617 33083 12683 33086
rect 13629 33010 13695 33013
rect 14181 33010 14247 33013
rect 15840 33010 16000 33040
rect 13629 33008 14106 33010
rect 13629 32952 13634 33008
rect 13690 32952 14106 33008
rect 13629 32950 14106 32952
rect 13629 32947 13695 32950
rect 14046 32874 14106 32950
rect 14181 33008 16000 33010
rect 14181 32952 14186 33008
rect 14242 32952 16000 33008
rect 14181 32950 16000 32952
rect 14181 32947 14247 32950
rect 15840 32920 16000 32950
rect 14046 32814 15164 32874
rect 15104 32738 15164 32814
rect 15840 32738 16000 32768
rect 15104 32678 16000 32738
rect 4372 32672 4688 32673
rect 4372 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4688 32672
rect 4372 32607 4688 32608
rect 7799 32672 8115 32673
rect 7799 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8115 32672
rect 7799 32607 8115 32608
rect 11226 32672 11542 32673
rect 11226 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11542 32672
rect 11226 32607 11542 32608
rect 14653 32672 14969 32673
rect 14653 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14969 32672
rect 15840 32648 16000 32678
rect 14653 32607 14969 32608
rect 0 32466 160 32496
rect 749 32466 815 32469
rect 0 32464 815 32466
rect 0 32408 754 32464
rect 810 32408 815 32464
rect 0 32406 815 32408
rect 0 32376 160 32406
rect 749 32403 815 32406
rect 11053 32466 11119 32469
rect 12014 32466 12020 32468
rect 11053 32464 12020 32466
rect 11053 32408 11058 32464
rect 11114 32408 12020 32464
rect 11053 32406 12020 32408
rect 11053 32403 11119 32406
rect 12014 32404 12020 32406
rect 12084 32466 12090 32468
rect 14273 32466 14339 32469
rect 15840 32466 16000 32496
rect 12084 32406 12450 32466
rect 12084 32404 12090 32406
rect 11789 32332 11855 32333
rect 11789 32330 11836 32332
rect 11744 32328 11836 32330
rect 11744 32272 11794 32328
rect 11744 32270 11836 32272
rect 11789 32268 11836 32270
rect 11900 32268 11906 32332
rect 12390 32330 12450 32406
rect 14273 32464 16000 32466
rect 14273 32408 14278 32464
rect 14334 32408 16000 32464
rect 14273 32406 16000 32408
rect 14273 32403 14339 32406
rect 15840 32376 16000 32406
rect 13537 32330 13603 32333
rect 12390 32328 13603 32330
rect 12390 32272 13542 32328
rect 13598 32272 13603 32328
rect 12390 32270 13603 32272
rect 11789 32267 11855 32268
rect 13537 32267 13603 32270
rect 14365 32194 14431 32197
rect 15840 32194 16000 32224
rect 14365 32192 16000 32194
rect 14365 32136 14370 32192
rect 14426 32136 16000 32192
rect 14365 32134 16000 32136
rect 14365 32131 14431 32134
rect 2659 32128 2975 32129
rect 2659 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2975 32128
rect 2659 32063 2975 32064
rect 6086 32128 6402 32129
rect 6086 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6402 32128
rect 6086 32063 6402 32064
rect 9513 32128 9829 32129
rect 9513 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9829 32128
rect 9513 32063 9829 32064
rect 12940 32128 13256 32129
rect 12940 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13256 32128
rect 15840 32104 16000 32134
rect 12940 32063 13256 32064
rect 10961 31922 11027 31925
rect 13721 31922 13787 31925
rect 10961 31920 13787 31922
rect 10961 31864 10966 31920
rect 11022 31864 13726 31920
rect 13782 31864 13787 31920
rect 10961 31862 13787 31864
rect 10961 31859 11027 31862
rect 13721 31859 13787 31862
rect 13905 31922 13971 31925
rect 15840 31922 16000 31952
rect 13905 31920 16000 31922
rect 13905 31864 13910 31920
rect 13966 31864 16000 31920
rect 13905 31862 16000 31864
rect 13905 31859 13971 31862
rect 15840 31832 16000 31862
rect 12617 31788 12683 31789
rect 12566 31786 12572 31788
rect 12526 31726 12572 31786
rect 12636 31784 12683 31788
rect 12678 31728 12683 31784
rect 12566 31724 12572 31726
rect 12636 31724 12683 31728
rect 12617 31723 12683 31724
rect 0 31650 160 31680
rect 1393 31650 1459 31653
rect 0 31648 1459 31650
rect 0 31592 1398 31648
rect 1454 31592 1459 31648
rect 0 31590 1459 31592
rect 0 31560 160 31590
rect 1393 31587 1459 31590
rect 15101 31650 15167 31653
rect 15840 31650 16000 31680
rect 15101 31648 16000 31650
rect 15101 31592 15106 31648
rect 15162 31592 16000 31648
rect 15101 31590 16000 31592
rect 15101 31587 15167 31590
rect 4372 31584 4688 31585
rect 4372 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4688 31584
rect 4372 31519 4688 31520
rect 7799 31584 8115 31585
rect 7799 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8115 31584
rect 7799 31519 8115 31520
rect 11226 31584 11542 31585
rect 11226 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11542 31584
rect 11226 31519 11542 31520
rect 14653 31584 14969 31585
rect 14653 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14969 31584
rect 15840 31560 16000 31590
rect 14653 31519 14969 31520
rect 10317 31378 10383 31381
rect 12985 31378 13051 31381
rect 10317 31376 13051 31378
rect 10317 31320 10322 31376
rect 10378 31320 12990 31376
rect 13046 31320 13051 31376
rect 10317 31318 13051 31320
rect 10317 31315 10383 31318
rect 12985 31315 13051 31318
rect 13997 31378 14063 31381
rect 15840 31378 16000 31408
rect 13997 31376 16000 31378
rect 13997 31320 14002 31376
rect 14058 31320 16000 31376
rect 13997 31318 16000 31320
rect 13997 31315 14063 31318
rect 15840 31288 16000 31318
rect 8753 31242 8819 31245
rect 13445 31242 13511 31245
rect 8753 31240 13511 31242
rect 8753 31184 8758 31240
rect 8814 31184 13450 31240
rect 13506 31184 13511 31240
rect 8753 31182 13511 31184
rect 8753 31179 8819 31182
rect 13445 31179 13511 31182
rect 11513 31106 11579 31109
rect 12433 31106 12499 31109
rect 11513 31104 12499 31106
rect 11513 31048 11518 31104
rect 11574 31048 12438 31104
rect 12494 31048 12499 31104
rect 11513 31046 12499 31048
rect 11513 31043 11579 31046
rect 12433 31043 12499 31046
rect 13353 31106 13419 31109
rect 15840 31106 16000 31136
rect 13353 31104 16000 31106
rect 13353 31048 13358 31104
rect 13414 31048 16000 31104
rect 13353 31046 16000 31048
rect 13353 31043 13419 31046
rect 2659 31040 2975 31041
rect 2659 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2975 31040
rect 2659 30975 2975 30976
rect 6086 31040 6402 31041
rect 6086 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6402 31040
rect 6086 30975 6402 30976
rect 9513 31040 9829 31041
rect 9513 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9829 31040
rect 9513 30975 9829 30976
rect 12940 31040 13256 31041
rect 12940 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13256 31040
rect 15840 31016 16000 31046
rect 12940 30975 13256 30976
rect 0 30834 160 30864
rect 749 30834 815 30837
rect 0 30832 815 30834
rect 0 30776 754 30832
rect 810 30776 815 30832
rect 0 30774 815 30776
rect 0 30744 160 30774
rect 749 30771 815 30774
rect 13905 30834 13971 30837
rect 15840 30834 16000 30864
rect 13905 30832 16000 30834
rect 13905 30776 13910 30832
rect 13966 30776 16000 30832
rect 13905 30774 16000 30776
rect 13905 30771 13971 30774
rect 15840 30744 16000 30774
rect 15101 30562 15167 30565
rect 15840 30562 16000 30592
rect 15101 30560 16000 30562
rect 15101 30504 15106 30560
rect 15162 30504 16000 30560
rect 15101 30502 16000 30504
rect 15101 30499 15167 30502
rect 4372 30496 4688 30497
rect 4372 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4688 30496
rect 4372 30431 4688 30432
rect 7799 30496 8115 30497
rect 7799 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8115 30496
rect 7799 30431 8115 30432
rect 11226 30496 11542 30497
rect 11226 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11542 30496
rect 11226 30431 11542 30432
rect 14653 30496 14969 30497
rect 14653 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14969 30496
rect 15840 30472 16000 30502
rect 14653 30431 14969 30432
rect 12893 30290 12959 30293
rect 13353 30290 13419 30293
rect 15840 30290 16000 30320
rect 12893 30288 13186 30290
rect 12893 30232 12898 30288
rect 12954 30232 13186 30288
rect 12893 30230 13186 30232
rect 12893 30227 12959 30230
rect 13126 30154 13186 30230
rect 13353 30288 16000 30290
rect 13353 30232 13358 30288
rect 13414 30232 16000 30288
rect 13353 30230 16000 30232
rect 13353 30227 13419 30230
rect 15840 30200 16000 30230
rect 13126 30094 14290 30154
rect 0 30018 160 30048
rect 749 30018 815 30021
rect 0 30016 815 30018
rect 0 29960 754 30016
rect 810 29960 815 30016
rect 0 29958 815 29960
rect 14230 30018 14290 30094
rect 15840 30018 16000 30048
rect 14230 29958 16000 30018
rect 0 29928 160 29958
rect 749 29955 815 29958
rect 2659 29952 2975 29953
rect 2659 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2975 29952
rect 2659 29887 2975 29888
rect 6086 29952 6402 29953
rect 6086 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6402 29952
rect 6086 29887 6402 29888
rect 9513 29952 9829 29953
rect 9513 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9829 29952
rect 9513 29887 9829 29888
rect 12940 29952 13256 29953
rect 12940 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13256 29952
rect 15840 29928 16000 29958
rect 12940 29887 13256 29888
rect 11605 29882 11671 29885
rect 11605 29880 12450 29882
rect 11605 29824 11610 29880
rect 11666 29824 12450 29880
rect 11605 29822 12450 29824
rect 11605 29819 11671 29822
rect 12390 29610 12450 29822
rect 13629 29746 13695 29749
rect 15285 29746 15351 29749
rect 15840 29746 16000 29776
rect 13629 29744 15164 29746
rect 13629 29688 13634 29744
rect 13690 29688 15164 29744
rect 13629 29686 15164 29688
rect 13629 29683 13695 29686
rect 13905 29610 13971 29613
rect 12390 29608 13971 29610
rect 12390 29552 13910 29608
rect 13966 29552 13971 29608
rect 12390 29550 13971 29552
rect 13905 29547 13971 29550
rect 15104 29474 15164 29686
rect 15285 29744 16000 29746
rect 15285 29688 15290 29744
rect 15346 29688 16000 29744
rect 15285 29686 16000 29688
rect 15285 29683 15351 29686
rect 15840 29656 16000 29686
rect 15840 29474 16000 29504
rect 15104 29414 16000 29474
rect 4372 29408 4688 29409
rect 4372 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4688 29408
rect 4372 29343 4688 29344
rect 7799 29408 8115 29409
rect 7799 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8115 29408
rect 7799 29343 8115 29344
rect 11226 29408 11542 29409
rect 11226 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11542 29408
rect 11226 29343 11542 29344
rect 14653 29408 14969 29409
rect 14653 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14969 29408
rect 15840 29384 16000 29414
rect 14653 29343 14969 29344
rect 0 29202 160 29232
rect 749 29202 815 29205
rect 0 29200 815 29202
rect 0 29144 754 29200
rect 810 29144 815 29200
rect 0 29142 815 29144
rect 0 29112 160 29142
rect 749 29139 815 29142
rect 3969 29202 4035 29205
rect 12893 29202 12959 29205
rect 3969 29200 12959 29202
rect 3969 29144 3974 29200
rect 4030 29144 12898 29200
rect 12954 29144 12959 29200
rect 3969 29142 12959 29144
rect 3969 29139 4035 29142
rect 12893 29139 12959 29142
rect 14273 29202 14339 29205
rect 15840 29202 16000 29232
rect 14273 29200 16000 29202
rect 14273 29144 14278 29200
rect 14334 29144 16000 29200
rect 14273 29142 16000 29144
rect 14273 29139 14339 29142
rect 15840 29112 16000 29142
rect 8937 29066 9003 29069
rect 9213 29068 9279 29069
rect 9070 29066 9076 29068
rect 8937 29064 9076 29066
rect 8937 29008 8942 29064
rect 8998 29008 9076 29064
rect 8937 29006 9076 29008
rect 8937 29003 9003 29006
rect 9070 29004 9076 29006
rect 9140 29004 9146 29068
rect 9213 29064 9260 29068
rect 9324 29066 9330 29068
rect 9213 29008 9218 29064
rect 9213 29004 9260 29008
rect 9324 29006 9370 29066
rect 9324 29004 9330 29006
rect 9213 29003 9279 29004
rect 11973 28932 12039 28933
rect 11973 28928 12020 28932
rect 12084 28930 12090 28932
rect 14549 28930 14615 28933
rect 15840 28930 16000 28960
rect 11973 28872 11978 28928
rect 11973 28868 12020 28872
rect 12084 28870 12130 28930
rect 14549 28928 16000 28930
rect 14549 28872 14554 28928
rect 14610 28872 16000 28928
rect 14549 28870 16000 28872
rect 12084 28868 12090 28870
rect 11973 28867 12039 28868
rect 14549 28867 14615 28870
rect 2659 28864 2975 28865
rect 2659 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2975 28864
rect 2659 28799 2975 28800
rect 6086 28864 6402 28865
rect 6086 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6402 28864
rect 6086 28799 6402 28800
rect 9513 28864 9829 28865
rect 9513 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9829 28864
rect 9513 28799 9829 28800
rect 12940 28864 13256 28865
rect 12940 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13256 28864
rect 15840 28840 16000 28870
rect 12940 28799 13256 28800
rect 13629 28658 13695 28661
rect 14181 28658 14247 28661
rect 15840 28658 16000 28688
rect 13629 28656 14106 28658
rect 13629 28600 13634 28656
rect 13690 28600 14106 28656
rect 13629 28598 14106 28600
rect 13629 28595 13695 28598
rect 14046 28522 14106 28598
rect 14181 28656 16000 28658
rect 14181 28600 14186 28656
rect 14242 28600 16000 28656
rect 14181 28598 16000 28600
rect 14181 28595 14247 28598
rect 15840 28568 16000 28598
rect 14046 28462 15164 28522
rect 0 28386 160 28416
rect 749 28386 815 28389
rect 0 28384 815 28386
rect 0 28328 754 28384
rect 810 28328 815 28384
rect 0 28326 815 28328
rect 15104 28386 15164 28462
rect 15840 28386 16000 28416
rect 15104 28326 16000 28386
rect 0 28296 160 28326
rect 749 28323 815 28326
rect 4372 28320 4688 28321
rect 4372 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4688 28320
rect 4372 28255 4688 28256
rect 7799 28320 8115 28321
rect 7799 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8115 28320
rect 7799 28255 8115 28256
rect 11226 28320 11542 28321
rect 11226 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11542 28320
rect 11226 28255 11542 28256
rect 14653 28320 14969 28321
rect 14653 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14969 28320
rect 15840 28296 16000 28326
rect 14653 28255 14969 28256
rect 13813 28114 13879 28117
rect 15840 28114 16000 28144
rect 13813 28112 16000 28114
rect 13813 28056 13818 28112
rect 13874 28056 16000 28112
rect 13813 28054 16000 28056
rect 13813 28051 13879 28054
rect 15840 28024 16000 28054
rect 11789 27842 11855 27845
rect 14365 27842 14431 27845
rect 15840 27842 16000 27872
rect 11789 27840 12450 27842
rect 11789 27784 11794 27840
rect 11850 27784 12450 27840
rect 11789 27782 12450 27784
rect 11789 27779 11855 27782
rect 2659 27776 2975 27777
rect 2659 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2975 27776
rect 2659 27711 2975 27712
rect 6086 27776 6402 27777
rect 6086 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6402 27776
rect 6086 27711 6402 27712
rect 9513 27776 9829 27777
rect 9513 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9829 27776
rect 9513 27711 9829 27712
rect 1669 27708 1735 27709
rect 1669 27706 1716 27708
rect 1624 27704 1716 27706
rect 1624 27648 1674 27704
rect 1624 27646 1716 27648
rect 1669 27644 1716 27646
rect 1780 27644 1786 27708
rect 1669 27643 1735 27644
rect 0 27570 160 27600
rect 1485 27570 1551 27573
rect 0 27568 1551 27570
rect 0 27512 1490 27568
rect 1546 27512 1551 27568
rect 0 27510 1551 27512
rect 0 27480 160 27510
rect 1485 27507 1551 27510
rect 12390 27298 12450 27782
rect 14365 27840 16000 27842
rect 14365 27784 14370 27840
rect 14426 27784 16000 27840
rect 14365 27782 16000 27784
rect 14365 27779 14431 27782
rect 12940 27776 13256 27777
rect 12940 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13256 27776
rect 15840 27752 16000 27782
rect 12940 27711 13256 27712
rect 13629 27570 13695 27573
rect 14181 27570 14247 27573
rect 15840 27570 16000 27600
rect 13629 27568 14106 27570
rect 13629 27512 13634 27568
rect 13690 27512 14106 27568
rect 13629 27510 14106 27512
rect 13629 27507 13695 27510
rect 14046 27434 14106 27510
rect 14181 27568 16000 27570
rect 14181 27512 14186 27568
rect 14242 27512 16000 27568
rect 14181 27510 16000 27512
rect 14181 27507 14247 27510
rect 15840 27480 16000 27510
rect 14046 27374 15164 27434
rect 12985 27298 13051 27301
rect 12390 27296 13051 27298
rect 12390 27240 12990 27296
rect 13046 27240 13051 27296
rect 12390 27238 13051 27240
rect 15104 27298 15164 27374
rect 15840 27298 16000 27328
rect 15104 27238 16000 27298
rect 12985 27235 13051 27238
rect 4372 27232 4688 27233
rect 4372 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4688 27232
rect 4372 27167 4688 27168
rect 7799 27232 8115 27233
rect 7799 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8115 27232
rect 7799 27167 8115 27168
rect 11226 27232 11542 27233
rect 11226 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11542 27232
rect 11226 27167 11542 27168
rect 14653 27232 14969 27233
rect 14653 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14969 27232
rect 15840 27208 16000 27238
rect 14653 27167 14969 27168
rect 12525 27026 12591 27029
rect 13353 27026 13419 27029
rect 12525 27024 13419 27026
rect 12525 26968 12530 27024
rect 12586 26968 13358 27024
rect 13414 26968 13419 27024
rect 12525 26966 13419 26968
rect 12525 26963 12591 26966
rect 13353 26963 13419 26966
rect 13905 27026 13971 27029
rect 15840 27026 16000 27056
rect 13905 27024 16000 27026
rect 13905 26968 13910 27024
rect 13966 26968 16000 27024
rect 13905 26966 16000 26968
rect 13905 26963 13971 26966
rect 15840 26936 16000 26966
rect 0 26754 160 26784
rect 749 26754 815 26757
rect 0 26752 815 26754
rect 0 26696 754 26752
rect 810 26696 815 26752
rect 0 26694 815 26696
rect 0 26664 160 26694
rect 749 26691 815 26694
rect 13813 26754 13879 26757
rect 15840 26754 16000 26784
rect 13813 26752 16000 26754
rect 13813 26696 13818 26752
rect 13874 26696 16000 26752
rect 13813 26694 16000 26696
rect 13813 26691 13879 26694
rect 2659 26688 2975 26689
rect 2659 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2975 26688
rect 2659 26623 2975 26624
rect 6086 26688 6402 26689
rect 6086 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6402 26688
rect 6086 26623 6402 26624
rect 9513 26688 9829 26689
rect 9513 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9829 26688
rect 9513 26623 9829 26624
rect 12940 26688 13256 26689
rect 12940 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13256 26688
rect 15840 26664 16000 26694
rect 12940 26623 13256 26624
rect 5206 26420 5212 26484
rect 5276 26482 5282 26484
rect 12157 26482 12223 26485
rect 5276 26480 12223 26482
rect 5276 26424 12162 26480
rect 12218 26424 12223 26480
rect 5276 26422 12223 26424
rect 5276 26420 5282 26422
rect 12157 26419 12223 26422
rect 14917 26482 14983 26485
rect 15840 26482 16000 26512
rect 14917 26480 16000 26482
rect 14917 26424 14922 26480
rect 14978 26424 16000 26480
rect 14917 26422 16000 26424
rect 14917 26419 14983 26422
rect 15840 26392 16000 26422
rect 8753 26346 8819 26349
rect 8886 26346 8892 26348
rect 8753 26344 8892 26346
rect 8753 26288 8758 26344
rect 8814 26288 8892 26344
rect 8753 26286 8892 26288
rect 8753 26283 8819 26286
rect 8886 26284 8892 26286
rect 8956 26284 8962 26348
rect 14414 26286 15164 26346
rect 1485 26210 1551 26213
rect 798 26208 1551 26210
rect 798 26152 1490 26208
rect 1546 26152 1551 26208
rect 798 26150 1551 26152
rect 0 25938 160 25968
rect 798 25938 858 26150
rect 1485 26147 1551 26150
rect 13261 26210 13327 26213
rect 14414 26210 14474 26286
rect 13261 26208 14474 26210
rect 13261 26152 13266 26208
rect 13322 26152 14474 26208
rect 13261 26150 14474 26152
rect 15104 26210 15164 26286
rect 15840 26210 16000 26240
rect 15104 26150 16000 26210
rect 13261 26147 13327 26150
rect 4372 26144 4688 26145
rect 4372 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4688 26144
rect 4372 26079 4688 26080
rect 7799 26144 8115 26145
rect 7799 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8115 26144
rect 7799 26079 8115 26080
rect 11226 26144 11542 26145
rect 11226 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11542 26144
rect 11226 26079 11542 26080
rect 14653 26144 14969 26145
rect 14653 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14969 26144
rect 15840 26120 16000 26150
rect 14653 26079 14969 26080
rect 12801 26074 12867 26077
rect 11654 26072 12867 26074
rect 11654 26016 12806 26072
rect 12862 26016 12867 26072
rect 11654 26014 12867 26016
rect 0 25878 858 25938
rect 9949 25938 10015 25941
rect 11654 25938 11714 26014
rect 12801 26011 12867 26014
rect 9949 25936 11714 25938
rect 9949 25880 9954 25936
rect 10010 25880 11714 25936
rect 9949 25878 11714 25880
rect 12341 25938 12407 25941
rect 15840 25938 16000 25968
rect 12341 25936 16000 25938
rect 12341 25880 12346 25936
rect 12402 25880 16000 25936
rect 12341 25878 16000 25880
rect 0 25848 160 25878
rect 9949 25875 10015 25878
rect 12341 25875 12407 25878
rect 15840 25848 16000 25878
rect 15285 25666 15351 25669
rect 15840 25666 16000 25696
rect 15285 25664 16000 25666
rect 15285 25608 15290 25664
rect 15346 25608 16000 25664
rect 15285 25606 16000 25608
rect 15285 25603 15351 25606
rect 2659 25600 2975 25601
rect 2659 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2975 25600
rect 2659 25535 2975 25536
rect 6086 25600 6402 25601
rect 6086 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6402 25600
rect 6086 25535 6402 25536
rect 9513 25600 9829 25601
rect 9513 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9829 25600
rect 9513 25535 9829 25536
rect 12940 25600 13256 25601
rect 12940 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13256 25600
rect 15840 25576 16000 25606
rect 12940 25535 13256 25536
rect 13813 25394 13879 25397
rect 15840 25394 16000 25424
rect 13813 25392 16000 25394
rect 13813 25336 13818 25392
rect 13874 25336 16000 25392
rect 13813 25334 16000 25336
rect 13813 25331 13879 25334
rect 15840 25304 16000 25334
rect 14365 25258 14431 25261
rect 14365 25256 15210 25258
rect 14365 25200 14370 25256
rect 14426 25200 15210 25256
rect 14365 25198 15210 25200
rect 14365 25195 14431 25198
rect 0 25122 160 25152
rect 749 25122 815 25125
rect 0 25120 815 25122
rect 0 25064 754 25120
rect 810 25064 815 25120
rect 0 25062 815 25064
rect 15150 25122 15210 25198
rect 15840 25122 16000 25152
rect 15150 25062 16000 25122
rect 0 25032 160 25062
rect 749 25059 815 25062
rect 4372 25056 4688 25057
rect 4372 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4688 25056
rect 4372 24991 4688 24992
rect 7799 25056 8115 25057
rect 7799 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8115 25056
rect 7799 24991 8115 24992
rect 11226 25056 11542 25057
rect 11226 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11542 25056
rect 11226 24991 11542 24992
rect 14653 25056 14969 25057
rect 14653 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14969 25056
rect 15840 25032 16000 25062
rect 14653 24991 14969 24992
rect 9765 24850 9831 24853
rect 10409 24850 10475 24853
rect 9765 24848 10475 24850
rect 9765 24792 9770 24848
rect 9826 24792 10414 24848
rect 10470 24792 10475 24848
rect 9765 24790 10475 24792
rect 9765 24787 9831 24790
rect 10409 24787 10475 24790
rect 15101 24850 15167 24853
rect 15840 24850 16000 24880
rect 15101 24848 16000 24850
rect 15101 24792 15106 24848
rect 15162 24792 16000 24848
rect 15101 24790 16000 24792
rect 15101 24787 15167 24790
rect 15840 24760 16000 24790
rect 9857 24714 9923 24717
rect 13721 24714 13787 24717
rect 9857 24712 13787 24714
rect 9857 24656 9862 24712
rect 9918 24656 13726 24712
rect 13782 24656 13787 24712
rect 9857 24654 13787 24656
rect 9857 24651 9923 24654
rect 13721 24651 13787 24654
rect 14181 24578 14247 24581
rect 15840 24578 16000 24608
rect 14181 24576 16000 24578
rect 14181 24520 14186 24576
rect 14242 24520 16000 24576
rect 14181 24518 16000 24520
rect 14181 24515 14247 24518
rect 2659 24512 2975 24513
rect 2659 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2975 24512
rect 2659 24447 2975 24448
rect 6086 24512 6402 24513
rect 6086 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6402 24512
rect 6086 24447 6402 24448
rect 9513 24512 9829 24513
rect 9513 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9829 24512
rect 9513 24447 9829 24448
rect 12940 24512 13256 24513
rect 12940 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13256 24512
rect 15840 24488 16000 24518
rect 12940 24447 13256 24448
rect 0 24306 160 24336
rect 749 24306 815 24309
rect 0 24304 815 24306
rect 0 24248 754 24304
rect 810 24248 815 24304
rect 0 24246 815 24248
rect 0 24216 160 24246
rect 749 24243 815 24246
rect 14365 24306 14431 24309
rect 15840 24306 16000 24336
rect 14365 24304 16000 24306
rect 14365 24248 14370 24304
rect 14426 24248 16000 24304
rect 14365 24246 16000 24248
rect 14365 24243 14431 24246
rect 15840 24216 16000 24246
rect 15101 24034 15167 24037
rect 15840 24034 16000 24064
rect 15101 24032 16000 24034
rect 15101 23976 15106 24032
rect 15162 23976 16000 24032
rect 15101 23974 16000 23976
rect 15101 23971 15167 23974
rect 4372 23968 4688 23969
rect 4372 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4688 23968
rect 4372 23903 4688 23904
rect 7799 23968 8115 23969
rect 7799 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8115 23968
rect 7799 23903 8115 23904
rect 11226 23968 11542 23969
rect 11226 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11542 23968
rect 11226 23903 11542 23904
rect 14653 23968 14969 23969
rect 14653 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14969 23968
rect 15840 23944 16000 23974
rect 14653 23903 14969 23904
rect 12065 23898 12131 23901
rect 13486 23898 13492 23900
rect 12065 23896 13492 23898
rect 12065 23840 12070 23896
rect 12126 23840 13492 23896
rect 12065 23838 13492 23840
rect 12065 23835 12131 23838
rect 13486 23836 13492 23838
rect 13556 23836 13562 23900
rect 14365 23762 14431 23765
rect 15840 23762 16000 23792
rect 14365 23760 16000 23762
rect 14365 23704 14370 23760
rect 14426 23704 16000 23760
rect 14365 23702 16000 23704
rect 14365 23699 14431 23702
rect 15840 23672 16000 23702
rect 0 23490 160 23520
rect 749 23490 815 23493
rect 0 23488 815 23490
rect 0 23432 754 23488
rect 810 23432 815 23488
rect 0 23430 815 23432
rect 0 23400 160 23430
rect 749 23427 815 23430
rect 14365 23490 14431 23493
rect 15840 23490 16000 23520
rect 14365 23488 16000 23490
rect 14365 23432 14370 23488
rect 14426 23432 16000 23488
rect 14365 23430 16000 23432
rect 14365 23427 14431 23430
rect 2659 23424 2975 23425
rect 2659 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2975 23424
rect 2659 23359 2975 23360
rect 6086 23424 6402 23425
rect 6086 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6402 23424
rect 6086 23359 6402 23360
rect 9513 23424 9829 23425
rect 9513 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9829 23424
rect 9513 23359 9829 23360
rect 12940 23424 13256 23425
rect 12940 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13256 23424
rect 15840 23400 16000 23430
rect 12940 23359 13256 23360
rect 8477 23218 8543 23221
rect 11145 23218 11211 23221
rect 8477 23216 11211 23218
rect 8477 23160 8482 23216
rect 8538 23160 11150 23216
rect 11206 23160 11211 23216
rect 8477 23158 11211 23160
rect 8477 23155 8543 23158
rect 11145 23155 11211 23158
rect 14365 23218 14431 23221
rect 15840 23218 16000 23248
rect 14365 23216 16000 23218
rect 14365 23160 14370 23216
rect 14426 23160 16000 23216
rect 14365 23158 16000 23160
rect 14365 23155 14431 23158
rect 15840 23128 16000 23158
rect 8477 23082 8543 23085
rect 13445 23082 13511 23085
rect 8477 23080 13511 23082
rect 8477 23024 8482 23080
rect 8538 23024 13450 23080
rect 13506 23024 13511 23080
rect 8477 23022 13511 23024
rect 8477 23019 8543 23022
rect 13445 23019 13511 23022
rect 15101 22946 15167 22949
rect 15840 22946 16000 22976
rect 15101 22944 16000 22946
rect 15101 22888 15106 22944
rect 15162 22888 16000 22944
rect 15101 22886 16000 22888
rect 15101 22883 15167 22886
rect 4372 22880 4688 22881
rect 4372 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4688 22880
rect 4372 22815 4688 22816
rect 7799 22880 8115 22881
rect 7799 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8115 22880
rect 7799 22815 8115 22816
rect 11226 22880 11542 22881
rect 11226 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11542 22880
rect 11226 22815 11542 22816
rect 14653 22880 14969 22881
rect 14653 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14969 22880
rect 15840 22856 16000 22886
rect 14653 22815 14969 22816
rect 0 22674 160 22704
rect 749 22674 815 22677
rect 15840 22674 16000 22704
rect 0 22672 815 22674
rect 0 22616 754 22672
rect 810 22616 815 22672
rect 0 22614 815 22616
rect 0 22584 160 22614
rect 749 22611 815 22614
rect 15104 22614 16000 22674
rect 15104 22538 15164 22614
rect 15840 22584 16000 22614
rect 14598 22478 15164 22538
rect 13721 22402 13787 22405
rect 13854 22402 13860 22404
rect 13721 22400 13860 22402
rect 13721 22344 13726 22400
rect 13782 22344 13860 22400
rect 13721 22342 13860 22344
rect 13721 22339 13787 22342
rect 13854 22340 13860 22342
rect 13924 22340 13930 22404
rect 14457 22402 14523 22405
rect 14598 22402 14658 22478
rect 14457 22400 14658 22402
rect 14457 22344 14462 22400
rect 14518 22344 14658 22400
rect 14457 22342 14658 22344
rect 14917 22402 14983 22405
rect 15840 22402 16000 22432
rect 14917 22400 16000 22402
rect 14917 22344 14922 22400
rect 14978 22344 16000 22400
rect 14917 22342 16000 22344
rect 14457 22339 14523 22342
rect 14917 22339 14983 22342
rect 2659 22336 2975 22337
rect 2659 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2975 22336
rect 2659 22271 2975 22272
rect 6086 22336 6402 22337
rect 6086 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6402 22336
rect 6086 22271 6402 22272
rect 9513 22336 9829 22337
rect 9513 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9829 22336
rect 9513 22271 9829 22272
rect 12940 22336 13256 22337
rect 12940 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13256 22336
rect 15840 22312 16000 22342
rect 12940 22271 13256 22272
rect 13445 22266 13511 22269
rect 15653 22266 15719 22269
rect 13445 22264 15719 22266
rect 13445 22208 13450 22264
rect 13506 22208 15658 22264
rect 15714 22208 15719 22264
rect 13445 22206 15719 22208
rect 13445 22203 13511 22206
rect 15653 22203 15719 22206
rect 14457 22130 14523 22133
rect 15840 22130 16000 22160
rect 14457 22128 16000 22130
rect 14457 22072 14462 22128
rect 14518 22072 16000 22128
rect 14457 22070 16000 22072
rect 14457 22067 14523 22070
rect 15840 22040 16000 22070
rect 9949 21994 10015 21997
rect 11830 21994 11836 21996
rect 9949 21992 11836 21994
rect 9949 21936 9954 21992
rect 10010 21936 11836 21992
rect 9949 21934 11836 21936
rect 9949 21931 10015 21934
rect 11830 21932 11836 21934
rect 11900 21932 11906 21996
rect 12065 21994 12131 21997
rect 15377 21996 15443 21997
rect 12566 21994 12572 21996
rect 12065 21992 12572 21994
rect 12065 21936 12070 21992
rect 12126 21936 12572 21992
rect 12065 21934 12572 21936
rect 12065 21931 12131 21934
rect 12566 21932 12572 21934
rect 12636 21932 12642 21996
rect 15326 21994 15332 21996
rect 15286 21934 15332 21994
rect 15396 21992 15443 21996
rect 15438 21936 15443 21992
rect 15326 21932 15332 21934
rect 15396 21932 15443 21936
rect 15377 21931 15443 21932
rect 0 21858 160 21888
rect 749 21858 815 21861
rect 0 21856 815 21858
rect 0 21800 754 21856
rect 810 21800 815 21856
rect 0 21798 815 21800
rect 0 21768 160 21798
rect 749 21795 815 21798
rect 8477 21858 8543 21861
rect 8845 21858 8911 21861
rect 8477 21856 8911 21858
rect 8477 21800 8482 21856
rect 8538 21800 8850 21856
rect 8906 21800 8911 21856
rect 8477 21798 8911 21800
rect 8477 21795 8543 21798
rect 8845 21795 8911 21798
rect 15101 21858 15167 21861
rect 15840 21858 16000 21888
rect 15101 21856 16000 21858
rect 15101 21800 15106 21856
rect 15162 21800 16000 21856
rect 15101 21798 16000 21800
rect 15101 21795 15167 21798
rect 4372 21792 4688 21793
rect 4372 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4688 21792
rect 4372 21727 4688 21728
rect 7799 21792 8115 21793
rect 7799 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8115 21792
rect 7799 21727 8115 21728
rect 11226 21792 11542 21793
rect 11226 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11542 21792
rect 11226 21727 11542 21728
rect 14653 21792 14969 21793
rect 14653 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14969 21792
rect 15840 21768 16000 21798
rect 14653 21727 14969 21728
rect 7281 21720 7347 21725
rect 7281 21664 7286 21720
rect 7342 21664 7347 21720
rect 7281 21659 7347 21664
rect 7284 21589 7344 21659
rect 7281 21584 7347 21589
rect 7281 21528 7286 21584
rect 7342 21528 7347 21584
rect 7281 21523 7347 21528
rect 14273 21586 14339 21589
rect 15840 21586 16000 21616
rect 14273 21584 16000 21586
rect 14273 21528 14278 21584
rect 14334 21528 16000 21584
rect 14273 21526 16000 21528
rect 14273 21523 14339 21526
rect 15840 21496 16000 21526
rect 1577 21450 1643 21453
rect 9489 21450 9555 21453
rect 1577 21448 9555 21450
rect 1577 21392 1582 21448
rect 1638 21392 9494 21448
rect 9550 21392 9555 21448
rect 1577 21390 9555 21392
rect 1577 21387 1643 21390
rect 9489 21387 9555 21390
rect 9857 21450 9923 21453
rect 11053 21450 11119 21453
rect 9857 21448 11119 21450
rect 9857 21392 9862 21448
rect 9918 21392 11058 21448
rect 11114 21392 11119 21448
rect 9857 21390 11119 21392
rect 9857 21387 9923 21390
rect 11053 21387 11119 21390
rect 13721 21314 13787 21317
rect 15840 21314 16000 21344
rect 13721 21312 16000 21314
rect 13721 21256 13726 21312
rect 13782 21256 16000 21312
rect 13721 21254 16000 21256
rect 13721 21251 13787 21254
rect 2659 21248 2975 21249
rect 2659 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2975 21248
rect 2659 21183 2975 21184
rect 6086 21248 6402 21249
rect 6086 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6402 21248
rect 6086 21183 6402 21184
rect 9513 21248 9829 21249
rect 9513 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9829 21248
rect 9513 21183 9829 21184
rect 12940 21248 13256 21249
rect 12940 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13256 21248
rect 15840 21224 16000 21254
rect 12940 21183 13256 21184
rect 13537 21180 13603 21181
rect 13486 21116 13492 21180
rect 13556 21178 13603 21180
rect 13556 21176 13648 21178
rect 13598 21120 13648 21176
rect 13556 21118 13648 21120
rect 13556 21116 13603 21118
rect 13537 21115 13603 21116
rect 0 21042 160 21072
rect 749 21042 815 21045
rect 0 21040 815 21042
rect 0 20984 754 21040
rect 810 20984 815 21040
rect 0 20982 815 20984
rect 0 20952 160 20982
rect 749 20979 815 20982
rect 13813 21042 13879 21045
rect 15840 21042 16000 21072
rect 13813 21040 16000 21042
rect 13813 20984 13818 21040
rect 13874 20984 16000 21040
rect 13813 20982 16000 20984
rect 13813 20979 13879 20982
rect 15840 20952 16000 20982
rect 12617 20906 12683 20909
rect 9630 20904 12683 20906
rect 9630 20848 12622 20904
rect 12678 20848 12683 20904
rect 9630 20846 12683 20848
rect 4372 20704 4688 20705
rect 4372 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4688 20704
rect 4372 20639 4688 20640
rect 7799 20704 8115 20705
rect 7799 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8115 20704
rect 7799 20639 8115 20640
rect 8201 20634 8267 20637
rect 9630 20634 9690 20846
rect 12617 20843 12683 20846
rect 11789 20770 11855 20773
rect 12750 20770 12756 20772
rect 11789 20768 12756 20770
rect 11789 20712 11794 20768
rect 11850 20712 12756 20768
rect 11789 20710 12756 20712
rect 11789 20707 11855 20710
rect 12750 20708 12756 20710
rect 12820 20708 12826 20772
rect 15285 20770 15351 20773
rect 15840 20770 16000 20800
rect 15285 20768 16000 20770
rect 15285 20712 15290 20768
rect 15346 20712 16000 20768
rect 15285 20710 16000 20712
rect 15285 20707 15351 20710
rect 11226 20704 11542 20705
rect 11226 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11542 20704
rect 11226 20639 11542 20640
rect 14653 20704 14969 20705
rect 14653 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14969 20704
rect 15840 20680 16000 20710
rect 14653 20639 14969 20640
rect 8201 20632 9690 20634
rect 8201 20576 8206 20632
rect 8262 20576 9690 20632
rect 8201 20574 9690 20576
rect 8201 20571 8267 20574
rect 5257 20498 5323 20501
rect 8702 20498 8708 20500
rect 5257 20496 8708 20498
rect 5257 20440 5262 20496
rect 5318 20440 8708 20496
rect 5257 20438 8708 20440
rect 5257 20435 5323 20438
rect 8702 20436 8708 20438
rect 8772 20436 8778 20500
rect 14089 20498 14155 20501
rect 15840 20498 16000 20528
rect 14089 20496 16000 20498
rect 14089 20440 14094 20496
rect 14150 20440 16000 20496
rect 14089 20438 16000 20440
rect 14089 20435 14155 20438
rect 15840 20408 16000 20438
rect 7281 20364 7347 20365
rect 7230 20362 7236 20364
rect 7190 20302 7236 20362
rect 7300 20360 7347 20364
rect 7342 20304 7347 20360
rect 7230 20300 7236 20302
rect 7300 20300 7347 20304
rect 7281 20299 7347 20300
rect 12433 20362 12499 20365
rect 12433 20360 13692 20362
rect 12433 20304 12438 20360
rect 12494 20304 13692 20360
rect 12433 20302 13692 20304
rect 12433 20299 12499 20302
rect 0 20226 160 20256
rect 13632 20229 13692 20302
rect 749 20226 815 20229
rect 0 20224 815 20226
rect 0 20168 754 20224
rect 810 20168 815 20224
rect 0 20166 815 20168
rect 0 20136 160 20166
rect 749 20163 815 20166
rect 13629 20224 13695 20229
rect 13629 20168 13634 20224
rect 13690 20168 13695 20224
rect 13629 20163 13695 20168
rect 14365 20226 14431 20229
rect 15840 20226 16000 20256
rect 14365 20224 16000 20226
rect 14365 20168 14370 20224
rect 14426 20168 16000 20224
rect 14365 20166 16000 20168
rect 14365 20163 14431 20166
rect 2659 20160 2975 20161
rect 2659 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2975 20160
rect 2659 20095 2975 20096
rect 6086 20160 6402 20161
rect 6086 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6402 20160
rect 6086 20095 6402 20096
rect 9513 20160 9829 20161
rect 9513 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9829 20160
rect 9513 20095 9829 20096
rect 12940 20160 13256 20161
rect 12940 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13256 20160
rect 15840 20136 16000 20166
rect 12940 20095 13256 20096
rect 9070 20090 9076 20092
rect 6502 20030 9076 20090
rect 5441 19954 5507 19957
rect 6502 19954 6562 20030
rect 9070 20028 9076 20030
rect 9140 20028 9146 20092
rect 5441 19952 6562 19954
rect 5441 19896 5446 19952
rect 5502 19896 6562 19952
rect 5441 19894 6562 19896
rect 7097 19954 7163 19957
rect 9254 19954 9260 19956
rect 7097 19952 9260 19954
rect 7097 19896 7102 19952
rect 7158 19896 9260 19952
rect 7097 19894 9260 19896
rect 5441 19891 5507 19894
rect 7097 19891 7163 19894
rect 9254 19892 9260 19894
rect 9324 19892 9330 19956
rect 15561 19954 15627 19957
rect 15840 19954 16000 19984
rect 15561 19952 16000 19954
rect 15561 19896 15566 19952
rect 15622 19896 16000 19952
rect 15561 19894 16000 19896
rect 15561 19891 15627 19894
rect 15840 19864 16000 19894
rect 7005 19818 7071 19821
rect 8201 19818 8267 19821
rect 7005 19816 8267 19818
rect 7005 19760 7010 19816
rect 7066 19760 8206 19816
rect 8262 19760 8267 19816
rect 7005 19758 8267 19760
rect 7005 19755 7071 19758
rect 8201 19755 8267 19758
rect 8702 19756 8708 19820
rect 8772 19818 8778 19820
rect 11237 19818 11303 19821
rect 8772 19816 11303 19818
rect 8772 19760 11242 19816
rect 11298 19760 11303 19816
rect 8772 19758 11303 19760
rect 8772 19756 8778 19758
rect 11237 19755 11303 19758
rect 11513 19818 11579 19821
rect 14641 19818 14707 19821
rect 11513 19816 11714 19818
rect 11513 19760 11518 19816
rect 11574 19760 11714 19816
rect 11513 19758 11714 19760
rect 11513 19755 11579 19758
rect 9121 19684 9187 19685
rect 9070 19620 9076 19684
rect 9140 19682 9187 19684
rect 9140 19680 9232 19682
rect 9182 19624 9232 19680
rect 9140 19622 9232 19624
rect 9140 19620 9187 19622
rect 9121 19619 9187 19620
rect 4372 19616 4688 19617
rect 4372 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4688 19616
rect 4372 19551 4688 19552
rect 7799 19616 8115 19617
rect 7799 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8115 19616
rect 7799 19551 8115 19552
rect 11226 19616 11542 19617
rect 11226 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11542 19616
rect 11226 19551 11542 19552
rect 0 19410 160 19440
rect 749 19410 815 19413
rect 0 19408 815 19410
rect 0 19352 754 19408
rect 810 19352 815 19408
rect 0 19350 815 19352
rect 0 19320 160 19350
rect 749 19347 815 19350
rect 11513 19410 11579 19413
rect 11654 19410 11714 19758
rect 14641 19816 15210 19818
rect 14641 19760 14646 19816
rect 14702 19760 15210 19816
rect 14641 19758 15210 19760
rect 14641 19755 14707 19758
rect 15150 19682 15210 19758
rect 15840 19682 16000 19712
rect 15150 19622 16000 19682
rect 14653 19616 14969 19617
rect 14653 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14969 19616
rect 15840 19592 16000 19622
rect 14653 19551 14969 19552
rect 11513 19408 11714 19410
rect 11513 19352 11518 19408
rect 11574 19352 11714 19408
rect 11513 19350 11714 19352
rect 12249 19410 12315 19413
rect 15840 19410 16000 19440
rect 12249 19408 16000 19410
rect 12249 19352 12254 19408
rect 12310 19352 16000 19408
rect 12249 19350 16000 19352
rect 11513 19347 11579 19350
rect 12249 19347 12315 19350
rect 15840 19320 16000 19350
rect 9673 19274 9739 19277
rect 10501 19276 10567 19277
rect 10501 19274 10548 19276
rect 9673 19272 10548 19274
rect 10612 19274 10618 19276
rect 9673 19216 9678 19272
rect 9734 19216 10506 19272
rect 9673 19214 10548 19216
rect 9673 19211 9739 19214
rect 10501 19212 10548 19214
rect 10612 19214 10694 19274
rect 10612 19212 10618 19214
rect 10501 19211 10567 19212
rect 11237 19138 11303 19141
rect 11789 19138 11855 19141
rect 11237 19136 11855 19138
rect 11237 19080 11242 19136
rect 11298 19080 11794 19136
rect 11850 19080 11855 19136
rect 11237 19078 11855 19080
rect 11237 19075 11303 19078
rect 11789 19075 11855 19078
rect 14365 19138 14431 19141
rect 15840 19138 16000 19168
rect 14365 19136 16000 19138
rect 14365 19080 14370 19136
rect 14426 19080 16000 19136
rect 14365 19078 16000 19080
rect 14365 19075 14431 19078
rect 2659 19072 2975 19073
rect 2659 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2975 19072
rect 2659 19007 2975 19008
rect 6086 19072 6402 19073
rect 6086 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6402 19072
rect 6086 19007 6402 19008
rect 9513 19072 9829 19073
rect 9513 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9829 19072
rect 9513 19007 9829 19008
rect 12940 19072 13256 19073
rect 12940 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13256 19072
rect 15840 19048 16000 19078
rect 12940 19007 13256 19008
rect 10133 19002 10199 19005
rect 12709 19002 12775 19005
rect 10133 19000 12775 19002
rect 10133 18944 10138 19000
rect 10194 18944 12714 19000
rect 12770 18944 12775 19000
rect 10133 18942 12775 18944
rect 10133 18939 10199 18942
rect 12709 18939 12775 18942
rect 9673 18866 9739 18869
rect 12801 18866 12867 18869
rect 9673 18864 12867 18866
rect 9673 18808 9678 18864
rect 9734 18808 12806 18864
rect 12862 18808 12867 18864
rect 9673 18806 12867 18808
rect 9673 18803 9739 18806
rect 12801 18803 12867 18806
rect 14457 18866 14523 18869
rect 15840 18866 16000 18896
rect 14457 18864 16000 18866
rect 14457 18808 14462 18864
rect 14518 18808 16000 18864
rect 14457 18806 16000 18808
rect 14457 18803 14523 18806
rect 15840 18776 16000 18806
rect 3693 18730 3759 18733
rect 6085 18730 6151 18733
rect 3693 18728 6151 18730
rect 3693 18672 3698 18728
rect 3754 18672 6090 18728
rect 6146 18672 6151 18728
rect 3693 18670 6151 18672
rect 3693 18667 3759 18670
rect 6085 18667 6151 18670
rect 10041 18730 10107 18733
rect 13169 18730 13235 18733
rect 10041 18728 13235 18730
rect 10041 18672 10046 18728
rect 10102 18672 13174 18728
rect 13230 18672 13235 18728
rect 10041 18670 13235 18672
rect 10041 18667 10107 18670
rect 13169 18667 13235 18670
rect 0 18594 160 18624
rect 749 18594 815 18597
rect 0 18592 815 18594
rect 0 18536 754 18592
rect 810 18536 815 18592
rect 0 18534 815 18536
rect 0 18504 160 18534
rect 749 18531 815 18534
rect 15101 18594 15167 18597
rect 15840 18594 16000 18624
rect 15101 18592 16000 18594
rect 15101 18536 15106 18592
rect 15162 18536 16000 18592
rect 15101 18534 16000 18536
rect 15101 18531 15167 18534
rect 4372 18528 4688 18529
rect 4372 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4688 18528
rect 4372 18463 4688 18464
rect 7799 18528 8115 18529
rect 7799 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8115 18528
rect 7799 18463 8115 18464
rect 11226 18528 11542 18529
rect 11226 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11542 18528
rect 11226 18463 11542 18464
rect 14653 18528 14969 18529
rect 14653 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14969 18528
rect 15840 18504 16000 18534
rect 14653 18463 14969 18464
rect 15840 18322 16000 18352
rect 15334 18262 16000 18322
rect 10358 18124 10364 18188
rect 10428 18186 10434 18188
rect 10501 18186 10567 18189
rect 10428 18184 10567 18186
rect 10428 18128 10506 18184
rect 10562 18128 10567 18184
rect 10428 18126 10567 18128
rect 10428 18124 10434 18126
rect 10501 18123 10567 18126
rect 13169 18186 13235 18189
rect 13486 18186 13492 18188
rect 13169 18184 13492 18186
rect 13169 18128 13174 18184
rect 13230 18128 13492 18184
rect 13169 18126 13492 18128
rect 13169 18123 13235 18126
rect 13486 18124 13492 18126
rect 13556 18124 13562 18188
rect 15193 18186 15259 18189
rect 15334 18186 15394 18262
rect 15840 18232 16000 18262
rect 15193 18184 15394 18186
rect 15193 18128 15198 18184
rect 15254 18128 15394 18184
rect 15193 18126 15394 18128
rect 15193 18123 15259 18126
rect 13353 18050 13419 18053
rect 15840 18050 16000 18080
rect 13353 18048 16000 18050
rect 13353 17992 13358 18048
rect 13414 17992 16000 18048
rect 13353 17990 16000 17992
rect 13353 17987 13419 17990
rect 2659 17984 2975 17985
rect 2659 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2975 17984
rect 2659 17919 2975 17920
rect 6086 17984 6402 17985
rect 6086 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6402 17984
rect 6086 17919 6402 17920
rect 9513 17984 9829 17985
rect 9513 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9829 17984
rect 9513 17919 9829 17920
rect 12940 17984 13256 17985
rect 12940 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13256 17984
rect 15840 17960 16000 17990
rect 12940 17919 13256 17920
rect 1485 17914 1551 17917
rect 798 17912 1551 17914
rect 798 17856 1490 17912
rect 1546 17856 1551 17912
rect 798 17854 1551 17856
rect 0 17778 160 17808
rect 798 17778 858 17854
rect 1485 17851 1551 17854
rect 11053 17914 11119 17917
rect 11830 17914 11836 17916
rect 11053 17912 11836 17914
rect 11053 17856 11058 17912
rect 11114 17856 11836 17912
rect 11053 17854 11836 17856
rect 11053 17851 11119 17854
rect 11830 17852 11836 17854
rect 11900 17852 11906 17916
rect 0 17718 858 17778
rect 11237 17776 11303 17781
rect 11237 17720 11242 17776
rect 11298 17720 11303 17776
rect 0 17688 160 17718
rect 11237 17715 11303 17720
rect 11421 17778 11487 17781
rect 15840 17778 16000 17808
rect 11421 17776 16000 17778
rect 11421 17720 11426 17776
rect 11482 17720 16000 17776
rect 11421 17718 16000 17720
rect 11421 17715 11487 17718
rect 11240 17642 11300 17715
rect 15840 17688 16000 17718
rect 11240 17582 15164 17642
rect 15104 17506 15164 17582
rect 15840 17506 16000 17536
rect 15104 17446 16000 17506
rect 4372 17440 4688 17441
rect 4372 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4688 17440
rect 4372 17375 4688 17376
rect 7799 17440 8115 17441
rect 7799 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8115 17440
rect 7799 17375 8115 17376
rect 11226 17440 11542 17441
rect 11226 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11542 17440
rect 11226 17375 11542 17376
rect 14653 17440 14969 17441
rect 14653 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14969 17440
rect 15840 17416 16000 17446
rect 14653 17375 14969 17376
rect 8201 17370 8267 17373
rect 8201 17368 11162 17370
rect 8201 17312 8206 17368
rect 8262 17312 11162 17368
rect 8201 17310 11162 17312
rect 8201 17307 8267 17310
rect 11102 17234 11162 17310
rect 11102 17174 12450 17234
rect 12390 17098 12450 17174
rect 13854 17172 13860 17236
rect 13924 17234 13930 17236
rect 14089 17234 14155 17237
rect 13924 17232 14155 17234
rect 13924 17176 14094 17232
rect 14150 17176 14155 17232
rect 13924 17174 14155 17176
rect 13924 17172 13930 17174
rect 14089 17171 14155 17174
rect 14273 17234 14339 17237
rect 15840 17234 16000 17264
rect 14273 17232 16000 17234
rect 14273 17176 14278 17232
rect 14334 17176 16000 17232
rect 14273 17174 16000 17176
rect 14273 17171 14339 17174
rect 15840 17144 16000 17174
rect 13629 17098 13695 17101
rect 12390 17096 13695 17098
rect 12390 17040 13634 17096
rect 13690 17040 13695 17096
rect 12390 17038 13695 17040
rect 13629 17035 13695 17038
rect 0 16962 160 16992
rect 749 16962 815 16965
rect 0 16960 815 16962
rect 0 16904 754 16960
rect 810 16904 815 16960
rect 0 16902 815 16904
rect 0 16872 160 16902
rect 749 16899 815 16902
rect 13813 16962 13879 16965
rect 15840 16962 16000 16992
rect 13813 16960 16000 16962
rect 13813 16904 13818 16960
rect 13874 16904 16000 16960
rect 13813 16902 16000 16904
rect 13813 16899 13879 16902
rect 2659 16896 2975 16897
rect 2659 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2975 16896
rect 2659 16831 2975 16832
rect 6086 16896 6402 16897
rect 6086 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6402 16896
rect 6086 16831 6402 16832
rect 9513 16896 9829 16897
rect 9513 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9829 16896
rect 9513 16831 9829 16832
rect 12940 16896 13256 16897
rect 12940 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13256 16896
rect 15840 16872 16000 16902
rect 12940 16831 13256 16832
rect 10869 16826 10935 16829
rect 12709 16826 12775 16829
rect 10869 16824 12775 16826
rect 10869 16768 10874 16824
rect 10930 16768 12714 16824
rect 12770 16768 12775 16824
rect 10869 16766 12775 16768
rect 10869 16763 10935 16766
rect 12709 16763 12775 16766
rect 10777 16690 10843 16693
rect 12985 16690 13051 16693
rect 10777 16688 13051 16690
rect 10777 16632 10782 16688
rect 10838 16632 12990 16688
rect 13046 16632 13051 16688
rect 10777 16630 13051 16632
rect 10777 16627 10843 16630
rect 12985 16627 13051 16630
rect 14273 16690 14339 16693
rect 15840 16690 16000 16720
rect 14273 16688 16000 16690
rect 14273 16632 14278 16688
rect 14334 16632 16000 16688
rect 14273 16630 16000 16632
rect 14273 16627 14339 16630
rect 15840 16600 16000 16630
rect 10542 16492 10548 16556
rect 10612 16554 10618 16556
rect 12065 16554 12131 16557
rect 10612 16552 12131 16554
rect 10612 16496 12070 16552
rect 12126 16496 12131 16552
rect 10612 16494 12131 16496
rect 10612 16492 10618 16494
rect 12065 16491 12131 16494
rect 12249 16554 12315 16557
rect 15193 16554 15259 16557
rect 12249 16552 15259 16554
rect 12249 16496 12254 16552
rect 12310 16496 15198 16552
rect 15254 16496 15259 16552
rect 12249 16494 15259 16496
rect 12249 16491 12315 16494
rect 15193 16491 15259 16494
rect 15101 16418 15167 16421
rect 15840 16418 16000 16448
rect 15101 16416 16000 16418
rect 15101 16360 15106 16416
rect 15162 16360 16000 16416
rect 15101 16358 16000 16360
rect 15101 16355 15167 16358
rect 4372 16352 4688 16353
rect 4372 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4688 16352
rect 4372 16287 4688 16288
rect 7799 16352 8115 16353
rect 7799 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8115 16352
rect 7799 16287 8115 16288
rect 11226 16352 11542 16353
rect 11226 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11542 16352
rect 11226 16287 11542 16288
rect 14653 16352 14969 16353
rect 14653 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14969 16352
rect 15840 16328 16000 16358
rect 14653 16287 14969 16288
rect 13077 16282 13143 16285
rect 13813 16284 13879 16285
rect 13486 16282 13492 16284
rect 13077 16280 13492 16282
rect 13077 16224 13082 16280
rect 13138 16224 13492 16280
rect 13077 16222 13492 16224
rect 13077 16219 13143 16222
rect 13486 16220 13492 16222
rect 13556 16220 13562 16284
rect 13813 16282 13860 16284
rect 13768 16280 13860 16282
rect 13768 16224 13818 16280
rect 13768 16222 13860 16224
rect 13813 16220 13860 16222
rect 13924 16220 13930 16284
rect 13813 16219 13879 16220
rect 0 16146 160 16176
rect 749 16146 815 16149
rect 0 16144 815 16146
rect 0 16088 754 16144
rect 810 16088 815 16144
rect 0 16086 815 16088
rect 0 16056 160 16086
rect 749 16083 815 16086
rect 7189 16146 7255 16149
rect 12709 16148 12775 16149
rect 8886 16146 8892 16148
rect 7189 16144 8892 16146
rect 7189 16088 7194 16144
rect 7250 16088 8892 16144
rect 7189 16086 8892 16088
rect 7189 16083 7255 16086
rect 8886 16084 8892 16086
rect 8956 16084 8962 16148
rect 12709 16146 12756 16148
rect 12664 16144 12756 16146
rect 12664 16088 12714 16144
rect 12664 16086 12756 16088
rect 12709 16084 12756 16086
rect 12820 16084 12826 16148
rect 13537 16146 13603 16149
rect 15840 16146 16000 16176
rect 13537 16144 16000 16146
rect 13537 16088 13542 16144
rect 13598 16088 16000 16144
rect 13537 16086 16000 16088
rect 12709 16083 12775 16084
rect 13537 16083 13603 16086
rect 15840 16056 16000 16086
rect 11789 15874 11855 15877
rect 12566 15874 12572 15876
rect 11789 15872 12572 15874
rect 11789 15816 11794 15872
rect 11850 15816 12572 15872
rect 11789 15814 12572 15816
rect 11789 15811 11855 15814
rect 12566 15812 12572 15814
rect 12636 15812 12642 15876
rect 13721 15874 13787 15877
rect 15840 15874 16000 15904
rect 13721 15872 16000 15874
rect 13721 15816 13726 15872
rect 13782 15816 16000 15872
rect 13721 15814 16000 15816
rect 13721 15811 13787 15814
rect 2659 15808 2975 15809
rect 2659 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2975 15808
rect 2659 15743 2975 15744
rect 6086 15808 6402 15809
rect 6086 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6402 15808
rect 6086 15743 6402 15744
rect 9513 15808 9829 15809
rect 9513 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9829 15808
rect 9513 15743 9829 15744
rect 12940 15808 13256 15809
rect 12940 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13256 15808
rect 15840 15784 16000 15814
rect 12940 15743 13256 15744
rect 11513 15602 11579 15605
rect 11646 15602 11652 15604
rect 11513 15600 11652 15602
rect 11513 15544 11518 15600
rect 11574 15544 11652 15600
rect 11513 15542 11652 15544
rect 11513 15539 11579 15542
rect 11646 15540 11652 15542
rect 11716 15540 11722 15604
rect 12341 15602 12407 15605
rect 14825 15602 14891 15605
rect 15840 15602 16000 15632
rect 12341 15600 14704 15602
rect 12341 15544 12346 15600
rect 12402 15544 14704 15600
rect 12341 15542 14704 15544
rect 12341 15539 12407 15542
rect 10409 15466 10475 15469
rect 14644 15466 14704 15542
rect 14825 15600 16000 15602
rect 14825 15544 14830 15600
rect 14886 15544 16000 15600
rect 14825 15542 16000 15544
rect 14825 15539 14891 15542
rect 15840 15512 16000 15542
rect 10409 15464 12450 15466
rect 10409 15408 10414 15464
rect 10470 15408 12450 15464
rect 10409 15406 12450 15408
rect 14644 15406 15164 15466
rect 10409 15403 10475 15406
rect 0 15330 160 15360
rect 841 15330 907 15333
rect 0 15328 907 15330
rect 0 15272 846 15328
rect 902 15272 907 15328
rect 0 15270 907 15272
rect 12390 15330 12450 15406
rect 13537 15330 13603 15333
rect 12390 15328 13603 15330
rect 12390 15272 13542 15328
rect 13598 15272 13603 15328
rect 12390 15270 13603 15272
rect 15104 15330 15164 15406
rect 15840 15330 16000 15360
rect 15104 15270 16000 15330
rect 0 15240 160 15270
rect 841 15267 907 15270
rect 13537 15267 13603 15270
rect 4372 15264 4688 15265
rect 4372 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4688 15264
rect 4372 15199 4688 15200
rect 7799 15264 8115 15265
rect 7799 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8115 15264
rect 7799 15199 8115 15200
rect 11226 15264 11542 15265
rect 11226 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11542 15264
rect 11226 15199 11542 15200
rect 14653 15264 14969 15265
rect 14653 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14969 15264
rect 15840 15240 16000 15270
rect 14653 15199 14969 15200
rect 12433 15194 12499 15197
rect 12433 15192 13692 15194
rect 12433 15136 12438 15192
rect 12494 15136 13692 15192
rect 12433 15134 13692 15136
rect 12433 15131 12499 15134
rect 10225 15058 10291 15061
rect 12893 15058 12959 15061
rect 10225 15056 12959 15058
rect 10225 15000 10230 15056
rect 10286 15000 12898 15056
rect 12954 15000 12959 15056
rect 10225 14998 12959 15000
rect 10225 14995 10291 14998
rect 12893 14995 12959 14998
rect 9121 14922 9187 14925
rect 11145 14922 11211 14925
rect 12709 14922 12775 14925
rect 9121 14920 12775 14922
rect 9121 14864 9126 14920
rect 9182 14864 11150 14920
rect 11206 14864 12714 14920
rect 12770 14864 12775 14920
rect 9121 14862 12775 14864
rect 9121 14859 9187 14862
rect 11145 14859 11211 14862
rect 12709 14859 12775 14862
rect 2659 14720 2975 14721
rect 2659 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2975 14720
rect 2659 14655 2975 14656
rect 6086 14720 6402 14721
rect 6086 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6402 14720
rect 6086 14655 6402 14656
rect 9513 14720 9829 14721
rect 9513 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9829 14720
rect 9513 14655 9829 14656
rect 12940 14720 13256 14721
rect 12940 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13256 14720
rect 12940 14655 13256 14656
rect 13632 14653 13692 15134
rect 14273 15058 14339 15061
rect 15840 15058 16000 15088
rect 14273 15056 16000 15058
rect 14273 15000 14278 15056
rect 14334 15000 16000 15056
rect 14273 14998 16000 15000
rect 14273 14995 14339 14998
rect 15840 14968 16000 14998
rect 14825 14786 14891 14789
rect 15840 14786 16000 14816
rect 14825 14784 16000 14786
rect 14825 14728 14830 14784
rect 14886 14728 16000 14784
rect 14825 14726 16000 14728
rect 14825 14723 14891 14726
rect 15840 14696 16000 14726
rect 13629 14648 13695 14653
rect 13629 14592 13634 14648
rect 13690 14592 13695 14648
rect 13629 14587 13695 14592
rect 0 14514 160 14544
rect 841 14514 907 14517
rect 0 14512 907 14514
rect 0 14456 846 14512
rect 902 14456 907 14512
rect 0 14454 907 14456
rect 0 14424 160 14454
rect 841 14451 907 14454
rect 10225 14514 10291 14517
rect 10358 14514 10364 14516
rect 10225 14512 10364 14514
rect 10225 14456 10230 14512
rect 10286 14456 10364 14512
rect 10225 14454 10364 14456
rect 10225 14451 10291 14454
rect 10358 14452 10364 14454
rect 10428 14452 10434 14516
rect 14181 14514 14247 14517
rect 15840 14514 16000 14544
rect 14181 14512 16000 14514
rect 14181 14456 14186 14512
rect 14242 14456 16000 14512
rect 14181 14454 16000 14456
rect 14181 14451 14247 14454
rect 15840 14424 16000 14454
rect 8201 14378 8267 14381
rect 15285 14378 15351 14381
rect 8201 14376 15351 14378
rect 8201 14320 8206 14376
rect 8262 14320 15290 14376
rect 15346 14320 15351 14376
rect 8201 14318 15351 14320
rect 8201 14315 8267 14318
rect 15285 14315 15351 14318
rect 8477 14242 8543 14245
rect 8937 14242 9003 14245
rect 8477 14240 9003 14242
rect 8477 14184 8482 14240
rect 8538 14184 8942 14240
rect 8998 14184 9003 14240
rect 8477 14182 9003 14184
rect 8477 14179 8543 14182
rect 8937 14179 9003 14182
rect 15101 14242 15167 14245
rect 15840 14242 16000 14272
rect 15101 14240 16000 14242
rect 15101 14184 15106 14240
rect 15162 14184 16000 14240
rect 15101 14182 16000 14184
rect 15101 14179 15167 14182
rect 4372 14176 4688 14177
rect 4372 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4688 14176
rect 4372 14111 4688 14112
rect 7799 14176 8115 14177
rect 7799 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8115 14176
rect 7799 14111 8115 14112
rect 11226 14176 11542 14177
rect 11226 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11542 14176
rect 11226 14111 11542 14112
rect 14653 14176 14969 14177
rect 14653 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14969 14176
rect 15840 14152 16000 14182
rect 14653 14111 14969 14112
rect 1669 14108 1735 14109
rect 1669 14106 1716 14108
rect 1624 14104 1716 14106
rect 1624 14048 1674 14104
rect 1624 14046 1716 14048
rect 1669 14044 1716 14046
rect 1780 14044 1786 14108
rect 1669 14043 1735 14044
rect 8293 13970 8359 13973
rect 15840 13970 16000 14000
rect 8250 13968 8359 13970
rect 8250 13912 8298 13968
rect 8354 13912 8359 13968
rect 8250 13907 8359 13912
rect 15150 13910 16000 13970
rect 0 13698 160 13728
rect 8250 13701 8310 13907
rect 9029 13834 9095 13837
rect 12525 13834 12591 13837
rect 13721 13836 13787 13837
rect 9029 13832 12591 13834
rect 9029 13776 9034 13832
rect 9090 13776 12530 13832
rect 12586 13776 12591 13832
rect 9029 13774 12591 13776
rect 9029 13771 9095 13774
rect 12525 13771 12591 13774
rect 13670 13772 13676 13836
rect 13740 13834 13787 13836
rect 14273 13834 14339 13837
rect 15150 13834 15210 13910
rect 15840 13880 16000 13910
rect 13740 13832 13832 13834
rect 13782 13776 13832 13832
rect 13740 13774 13832 13776
rect 14273 13832 15210 13834
rect 14273 13776 14278 13832
rect 14334 13776 15210 13832
rect 14273 13774 15210 13776
rect 13740 13772 13787 13774
rect 13721 13771 13787 13772
rect 14273 13771 14339 13774
rect 2497 13698 2563 13701
rect 0 13696 2563 13698
rect 0 13640 2502 13696
rect 2558 13640 2563 13696
rect 0 13638 2563 13640
rect 8250 13696 8359 13701
rect 8250 13640 8298 13696
rect 8354 13640 8359 13696
rect 8250 13638 8359 13640
rect 0 13608 160 13638
rect 2497 13635 2563 13638
rect 8293 13635 8359 13638
rect 13629 13698 13695 13701
rect 13997 13698 14063 13701
rect 15840 13698 16000 13728
rect 13629 13696 13738 13698
rect 13629 13640 13634 13696
rect 13690 13640 13738 13696
rect 13629 13635 13738 13640
rect 13997 13696 16000 13698
rect 13997 13640 14002 13696
rect 14058 13640 16000 13696
rect 13997 13638 16000 13640
rect 13997 13635 14063 13638
rect 2659 13632 2975 13633
rect 2659 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2975 13632
rect 2659 13567 2975 13568
rect 6086 13632 6402 13633
rect 6086 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6402 13632
rect 6086 13567 6402 13568
rect 9513 13632 9829 13633
rect 9513 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9829 13632
rect 9513 13567 9829 13568
rect 12940 13632 13256 13633
rect 12940 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13256 13632
rect 12940 13567 13256 13568
rect 10726 13500 10732 13564
rect 10796 13562 10802 13564
rect 11830 13562 11836 13564
rect 10796 13502 11836 13562
rect 10796 13500 10802 13502
rect 11830 13500 11836 13502
rect 11900 13500 11906 13564
rect 5257 13426 5323 13429
rect 9949 13426 10015 13429
rect 13077 13426 13143 13429
rect 5257 13424 9690 13426
rect 5257 13368 5262 13424
rect 5318 13368 9690 13424
rect 5257 13366 9690 13368
rect 5257 13363 5323 13366
rect 4372 13088 4688 13089
rect 4372 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4688 13088
rect 4372 13023 4688 13024
rect 7799 13088 8115 13089
rect 7799 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8115 13088
rect 7799 13023 8115 13024
rect 1945 13018 2011 13021
rect 982 13016 2011 13018
rect 982 12960 1950 13016
rect 2006 12960 2011 13016
rect 982 12958 2011 12960
rect 0 12882 160 12912
rect 982 12882 1042 12958
rect 1945 12955 2011 12958
rect 0 12822 1042 12882
rect 0 12792 160 12822
rect 3918 12820 3924 12884
rect 3988 12882 3994 12884
rect 7097 12882 7163 12885
rect 3988 12880 7163 12882
rect 3988 12824 7102 12880
rect 7158 12824 7163 12880
rect 3988 12822 7163 12824
rect 9630 12882 9690 13366
rect 9949 13424 13143 13426
rect 9949 13368 9954 13424
rect 10010 13368 13082 13424
rect 13138 13368 13143 13424
rect 9949 13366 13143 13368
rect 9949 13363 10015 13366
rect 13077 13363 13143 13366
rect 11421 13290 11487 13293
rect 12341 13290 12407 13293
rect 13077 13290 13143 13293
rect 11421 13288 12266 13290
rect 11421 13232 11426 13288
rect 11482 13232 12266 13288
rect 11421 13230 12266 13232
rect 11421 13227 11487 13230
rect 12206 13154 12266 13230
rect 12341 13288 13143 13290
rect 12341 13232 12346 13288
rect 12402 13232 13082 13288
rect 13138 13232 13143 13288
rect 12341 13230 13143 13232
rect 13678 13290 13738 13635
rect 15840 13608 16000 13638
rect 14181 13562 14247 13565
rect 15326 13562 15332 13564
rect 14181 13560 15332 13562
rect 14181 13504 14186 13560
rect 14242 13504 15332 13560
rect 14181 13502 15332 13504
rect 14181 13499 14247 13502
rect 15326 13500 15332 13502
rect 15396 13500 15402 13564
rect 13905 13426 13971 13429
rect 15840 13426 16000 13456
rect 13905 13424 16000 13426
rect 13905 13368 13910 13424
rect 13966 13368 16000 13424
rect 13905 13366 16000 13368
rect 13905 13363 13971 13366
rect 15840 13336 16000 13366
rect 13678 13230 14520 13290
rect 12341 13227 12407 13230
rect 13077 13227 13143 13230
rect 13261 13154 13327 13157
rect 12206 13152 13327 13154
rect 12206 13096 13266 13152
rect 13322 13096 13327 13152
rect 12206 13094 13327 13096
rect 13261 13091 13327 13094
rect 11226 13088 11542 13089
rect 11226 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11542 13088
rect 11226 13023 11542 13024
rect 14181 13018 14247 13021
rect 11608 13016 14247 13018
rect 11608 12960 14186 13016
rect 14242 12960 14247 13016
rect 11608 12958 14247 12960
rect 9765 12882 9831 12885
rect 11608 12882 11668 12958
rect 14181 12955 14247 12958
rect 9630 12880 11668 12882
rect 9630 12824 9770 12880
rect 9826 12824 11668 12880
rect 9630 12822 11668 12824
rect 13077 12882 13143 12885
rect 14460 12882 14520 13230
rect 15193 13154 15259 13157
rect 15840 13154 16000 13184
rect 15193 13152 16000 13154
rect 15193 13096 15198 13152
rect 15254 13096 16000 13152
rect 15193 13094 16000 13096
rect 15193 13091 15259 13094
rect 14653 13088 14969 13089
rect 14653 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14969 13088
rect 15840 13064 16000 13094
rect 14653 13023 14969 13024
rect 15840 12882 16000 12912
rect 13077 12880 14106 12882
rect 13077 12824 13082 12880
rect 13138 12824 14106 12880
rect 13077 12822 14106 12824
rect 14460 12822 16000 12882
rect 3988 12820 3994 12822
rect 7097 12819 7163 12822
rect 9765 12819 9831 12822
rect 13077 12819 13143 12822
rect 7649 12746 7715 12749
rect 13905 12746 13971 12749
rect 7649 12744 13971 12746
rect 7649 12688 7654 12744
rect 7710 12688 13910 12744
rect 13966 12688 13971 12744
rect 7649 12686 13971 12688
rect 7649 12683 7715 12686
rect 13905 12683 13971 12686
rect 12249 12610 12315 12613
rect 12566 12610 12572 12612
rect 12249 12608 12572 12610
rect 12249 12552 12254 12608
rect 12310 12552 12572 12608
rect 12249 12550 12572 12552
rect 12249 12547 12315 12550
rect 12566 12548 12572 12550
rect 12636 12548 12642 12612
rect 14046 12610 14106 12822
rect 15840 12792 16000 12822
rect 15840 12610 16000 12640
rect 14046 12550 16000 12610
rect 2659 12544 2975 12545
rect 2659 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2975 12544
rect 2659 12479 2975 12480
rect 6086 12544 6402 12545
rect 6086 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6402 12544
rect 6086 12479 6402 12480
rect 9513 12544 9829 12545
rect 9513 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9829 12544
rect 9513 12479 9829 12480
rect 12940 12544 13256 12545
rect 12940 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13256 12544
rect 15840 12520 16000 12550
rect 12940 12479 13256 12480
rect 12617 12474 12683 12477
rect 12750 12474 12756 12476
rect 12617 12472 12756 12474
rect 12617 12416 12622 12472
rect 12678 12416 12756 12472
rect 12617 12414 12756 12416
rect 12617 12411 12683 12414
rect 12750 12412 12756 12414
rect 12820 12412 12826 12476
rect 13854 12412 13860 12476
rect 13924 12474 13930 12476
rect 13997 12474 14063 12477
rect 13924 12472 14063 12474
rect 13924 12416 14002 12472
rect 14058 12416 14063 12472
rect 13924 12414 14063 12416
rect 13924 12412 13930 12414
rect 13997 12411 14063 12414
rect 9673 12338 9739 12341
rect 10777 12338 10843 12341
rect 11605 12340 11671 12341
rect 11605 12338 11652 12340
rect 9673 12336 10843 12338
rect 9673 12280 9678 12336
rect 9734 12280 10782 12336
rect 10838 12280 10843 12336
rect 9673 12278 10843 12280
rect 11560 12336 11652 12338
rect 11560 12280 11610 12336
rect 11560 12278 11652 12280
rect 9673 12275 9739 12278
rect 10777 12275 10843 12278
rect 11605 12276 11652 12278
rect 11716 12276 11722 12340
rect 11789 12338 11855 12341
rect 15840 12338 16000 12368
rect 11789 12336 16000 12338
rect 11789 12280 11794 12336
rect 11850 12280 16000 12336
rect 11789 12278 16000 12280
rect 11605 12275 11671 12276
rect 11789 12275 11855 12278
rect 15840 12248 16000 12278
rect 5901 12202 5967 12205
rect 9949 12202 10015 12205
rect 5901 12200 10015 12202
rect 5901 12144 5906 12200
rect 5962 12144 9954 12200
rect 10010 12144 10015 12200
rect 5901 12142 10015 12144
rect 5901 12139 5967 12142
rect 9949 12139 10015 12142
rect 0 12066 160 12096
rect 841 12066 907 12069
rect 15840 12066 16000 12096
rect 0 12064 907 12066
rect 0 12008 846 12064
rect 902 12008 907 12064
rect 0 12006 907 12008
rect 0 11976 160 12006
rect 841 12003 907 12006
rect 15150 12006 16000 12066
rect 4372 12000 4688 12001
rect 4372 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4688 12000
rect 4372 11935 4688 11936
rect 7799 12000 8115 12001
rect 7799 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8115 12000
rect 7799 11935 8115 11936
rect 11226 12000 11542 12001
rect 11226 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11542 12000
rect 11226 11935 11542 11936
rect 14653 12000 14969 12001
rect 14653 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14969 12000
rect 14653 11935 14969 11936
rect 15150 11933 15210 12006
rect 15840 11976 16000 12006
rect 15101 11928 15210 11933
rect 15101 11872 15106 11928
rect 15162 11872 15210 11928
rect 15101 11870 15210 11872
rect 15101 11867 15167 11870
rect 7230 11732 7236 11796
rect 7300 11794 7306 11796
rect 8753 11794 8819 11797
rect 12617 11794 12683 11797
rect 7300 11792 12683 11794
rect 7300 11736 8758 11792
rect 8814 11736 12622 11792
rect 12678 11736 12683 11792
rect 7300 11734 12683 11736
rect 7300 11732 7306 11734
rect 8753 11731 8819 11734
rect 12617 11731 12683 11734
rect 14089 11794 14155 11797
rect 15840 11794 16000 11824
rect 14089 11792 16000 11794
rect 14089 11736 14094 11792
rect 14150 11736 16000 11792
rect 14089 11734 16000 11736
rect 14089 11731 14155 11734
rect 15840 11704 16000 11734
rect 14273 11522 14339 11525
rect 15840 11522 16000 11552
rect 14273 11520 16000 11522
rect 14273 11464 14278 11520
rect 14334 11464 16000 11520
rect 14273 11462 16000 11464
rect 14273 11459 14339 11462
rect 2659 11456 2975 11457
rect 2659 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2975 11456
rect 2659 11391 2975 11392
rect 6086 11456 6402 11457
rect 6086 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6402 11456
rect 6086 11391 6402 11392
rect 9513 11456 9829 11457
rect 9513 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9829 11456
rect 9513 11391 9829 11392
rect 12940 11456 13256 11457
rect 12940 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13256 11456
rect 15840 11432 16000 11462
rect 12940 11391 13256 11392
rect 0 11250 160 11280
rect 841 11250 907 11253
rect 0 11248 907 11250
rect 0 11192 846 11248
rect 902 11192 907 11248
rect 0 11190 907 11192
rect 0 11160 160 11190
rect 841 11187 907 11190
rect 12341 11250 12407 11253
rect 15840 11250 16000 11280
rect 12341 11248 16000 11250
rect 12341 11192 12346 11248
rect 12402 11192 16000 11248
rect 12341 11190 16000 11192
rect 12341 11187 12407 11190
rect 15840 11160 16000 11190
rect 15193 10978 15259 10981
rect 15840 10978 16000 11008
rect 15193 10976 16000 10978
rect 15193 10920 15198 10976
rect 15254 10920 16000 10976
rect 15193 10918 16000 10920
rect 15193 10915 15259 10918
rect 4372 10912 4688 10913
rect 4372 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4688 10912
rect 4372 10847 4688 10848
rect 7799 10912 8115 10913
rect 7799 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8115 10912
rect 7799 10847 8115 10848
rect 11226 10912 11542 10913
rect 11226 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11542 10912
rect 11226 10847 11542 10848
rect 14653 10912 14969 10913
rect 14653 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14969 10912
rect 15840 10888 16000 10918
rect 14653 10847 14969 10848
rect 14181 10706 14247 10709
rect 15840 10706 16000 10736
rect 14181 10704 16000 10706
rect 14181 10648 14186 10704
rect 14242 10648 16000 10704
rect 14181 10646 16000 10648
rect 14181 10643 14247 10646
rect 15840 10616 16000 10646
rect 9949 10570 10015 10573
rect 14089 10570 14155 10573
rect 9949 10568 14155 10570
rect 9949 10512 9954 10568
rect 10010 10512 14094 10568
rect 14150 10512 14155 10568
rect 9949 10510 14155 10512
rect 9949 10507 10015 10510
rect 14089 10507 14155 10510
rect 0 10434 160 10464
rect 841 10434 907 10437
rect 0 10432 907 10434
rect 0 10376 846 10432
rect 902 10376 907 10432
rect 0 10374 907 10376
rect 0 10344 160 10374
rect 841 10371 907 10374
rect 11973 10434 12039 10437
rect 12198 10434 12204 10436
rect 11973 10432 12204 10434
rect 11973 10376 11978 10432
rect 12034 10376 12204 10432
rect 11973 10374 12204 10376
rect 11973 10371 12039 10374
rect 12198 10372 12204 10374
rect 12268 10372 12274 10436
rect 14641 10434 14707 10437
rect 15840 10434 16000 10464
rect 14641 10432 16000 10434
rect 14641 10376 14646 10432
rect 14702 10376 16000 10432
rect 14641 10374 16000 10376
rect 14641 10371 14707 10374
rect 2659 10368 2975 10369
rect 2659 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2975 10368
rect 2659 10303 2975 10304
rect 6086 10368 6402 10369
rect 6086 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6402 10368
rect 6086 10303 6402 10304
rect 9513 10368 9829 10369
rect 9513 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9829 10368
rect 9513 10303 9829 10304
rect 12940 10368 13256 10369
rect 12940 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13256 10368
rect 15840 10344 16000 10374
rect 12940 10303 13256 10304
rect 10225 10298 10291 10301
rect 12433 10298 12499 10301
rect 10225 10296 12499 10298
rect 10225 10240 10230 10296
rect 10286 10240 12438 10296
rect 12494 10240 12499 10296
rect 10225 10238 12499 10240
rect 10225 10235 10291 10238
rect 12433 10235 12499 10238
rect 9397 10162 9463 10165
rect 11973 10162 12039 10165
rect 12709 10162 12775 10165
rect 9397 10160 12775 10162
rect 9397 10104 9402 10160
rect 9458 10104 11978 10160
rect 12034 10104 12714 10160
rect 12770 10104 12775 10160
rect 9397 10102 12775 10104
rect 9397 10099 9463 10102
rect 11973 10099 12039 10102
rect 12709 10099 12775 10102
rect 13721 10162 13787 10165
rect 15840 10162 16000 10192
rect 13721 10160 16000 10162
rect 13721 10104 13726 10160
rect 13782 10104 16000 10160
rect 13721 10102 16000 10104
rect 13721 10099 13787 10102
rect 15840 10072 16000 10102
rect 9305 10026 9371 10029
rect 13445 10026 13511 10029
rect 9305 10024 13511 10026
rect 9305 9968 9310 10024
rect 9366 9968 13450 10024
rect 13506 9968 13511 10024
rect 9305 9966 13511 9968
rect 9305 9963 9371 9966
rect 13445 9963 13511 9966
rect 10501 9890 10567 9893
rect 10726 9890 10732 9892
rect 10501 9888 10732 9890
rect 10501 9832 10506 9888
rect 10562 9832 10732 9888
rect 10501 9830 10732 9832
rect 10501 9827 10567 9830
rect 10726 9828 10732 9830
rect 10796 9828 10802 9892
rect 11697 9890 11763 9893
rect 13905 9890 13971 9893
rect 11697 9888 13971 9890
rect 11697 9832 11702 9888
rect 11758 9832 13910 9888
rect 13966 9832 13971 9888
rect 11697 9830 13971 9832
rect 11697 9827 11763 9830
rect 13905 9827 13971 9830
rect 15101 9890 15167 9893
rect 15840 9890 16000 9920
rect 15101 9888 16000 9890
rect 15101 9832 15106 9888
rect 15162 9832 16000 9888
rect 15101 9830 16000 9832
rect 15101 9827 15167 9830
rect 4372 9824 4688 9825
rect 4372 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4688 9824
rect 4372 9759 4688 9760
rect 7799 9824 8115 9825
rect 7799 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8115 9824
rect 7799 9759 8115 9760
rect 11226 9824 11542 9825
rect 11226 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11542 9824
rect 11226 9759 11542 9760
rect 14653 9824 14969 9825
rect 14653 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14969 9824
rect 15840 9800 16000 9830
rect 14653 9759 14969 9760
rect 4981 9754 5047 9757
rect 5717 9754 5783 9757
rect 4981 9752 5783 9754
rect 4981 9696 4986 9752
rect 5042 9696 5722 9752
rect 5778 9696 5783 9752
rect 4981 9694 5783 9696
rect 4981 9691 5047 9694
rect 5717 9691 5783 9694
rect 11789 9754 11855 9757
rect 12525 9754 12591 9757
rect 11789 9752 12591 9754
rect 11789 9696 11794 9752
rect 11850 9696 12530 9752
rect 12586 9696 12591 9752
rect 11789 9694 12591 9696
rect 11789 9691 11855 9694
rect 12525 9691 12591 9694
rect 0 9618 160 9648
rect 933 9618 999 9621
rect 0 9616 999 9618
rect 0 9560 938 9616
rect 994 9560 999 9616
rect 0 9558 999 9560
rect 0 9528 160 9558
rect 933 9555 999 9558
rect 10225 9618 10291 9621
rect 10961 9618 11027 9621
rect 10225 9616 11027 9618
rect 10225 9560 10230 9616
rect 10286 9560 10966 9616
rect 11022 9560 11027 9616
rect 10225 9558 11027 9560
rect 10225 9555 10291 9558
rect 10961 9555 11027 9558
rect 11329 9618 11395 9621
rect 12709 9618 12775 9621
rect 15840 9618 16000 9648
rect 11329 9616 12128 9618
rect 11329 9560 11334 9616
rect 11390 9560 12128 9616
rect 11329 9558 12128 9560
rect 11329 9555 11395 9558
rect 10409 9346 10475 9349
rect 11053 9346 11119 9349
rect 11329 9346 11395 9349
rect 10409 9344 10978 9346
rect 10409 9288 10414 9344
rect 10470 9288 10978 9344
rect 10409 9286 10978 9288
rect 10409 9283 10475 9286
rect 2659 9280 2975 9281
rect 2659 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2975 9280
rect 2659 9215 2975 9216
rect 6086 9280 6402 9281
rect 6086 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6402 9280
rect 6086 9215 6402 9216
rect 9513 9280 9829 9281
rect 9513 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9829 9280
rect 9513 9215 9829 9216
rect 10317 9210 10383 9213
rect 10542 9210 10548 9212
rect 10317 9208 10548 9210
rect 10317 9152 10322 9208
rect 10378 9152 10548 9208
rect 10317 9150 10548 9152
rect 10317 9147 10383 9150
rect 10542 9148 10548 9150
rect 10612 9148 10618 9212
rect 10918 9210 10978 9286
rect 11053 9344 11395 9346
rect 11053 9288 11058 9344
rect 11114 9288 11334 9344
rect 11390 9288 11395 9344
rect 11053 9286 11395 9288
rect 11053 9283 11119 9286
rect 11329 9283 11395 9286
rect 11513 9346 11579 9349
rect 11646 9346 11652 9348
rect 11513 9344 11652 9346
rect 11513 9288 11518 9344
rect 11574 9288 11652 9344
rect 11513 9286 11652 9288
rect 11513 9283 11579 9286
rect 11646 9284 11652 9286
rect 11716 9284 11722 9348
rect 12068 9346 12128 9558
rect 12709 9616 16000 9618
rect 12709 9560 12714 9616
rect 12770 9560 16000 9616
rect 12709 9558 16000 9560
rect 12709 9555 12775 9558
rect 15840 9528 16000 9558
rect 12249 9484 12315 9485
rect 12198 9420 12204 9484
rect 12268 9482 12315 9484
rect 13261 9482 13327 9485
rect 13813 9482 13879 9485
rect 12268 9480 12360 9482
rect 12310 9424 12360 9480
rect 12268 9422 12360 9424
rect 13261 9480 13879 9482
rect 13261 9424 13266 9480
rect 13322 9424 13818 9480
rect 13874 9424 13879 9480
rect 13261 9422 13879 9424
rect 12268 9420 12315 9422
rect 12249 9419 12315 9420
rect 13261 9419 13327 9422
rect 13813 9419 13879 9422
rect 12198 9346 12204 9348
rect 12068 9286 12204 9346
rect 12198 9284 12204 9286
rect 12268 9284 12274 9348
rect 14457 9346 14523 9349
rect 15840 9346 16000 9376
rect 14457 9344 16000 9346
rect 14457 9288 14462 9344
rect 14518 9288 16000 9344
rect 14457 9286 16000 9288
rect 14457 9283 14523 9286
rect 12940 9280 13256 9281
rect 12940 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13256 9280
rect 15840 9256 16000 9286
rect 12940 9215 13256 9216
rect 11973 9210 12039 9213
rect 10918 9208 12039 9210
rect 10918 9152 11978 9208
rect 12034 9152 12039 9208
rect 10918 9150 12039 9152
rect 11973 9147 12039 9150
rect 12617 9210 12683 9213
rect 12750 9210 12756 9212
rect 12617 9208 12756 9210
rect 12617 9152 12622 9208
rect 12678 9152 12756 9208
rect 12617 9150 12756 9152
rect 12617 9147 12683 9150
rect 12750 9148 12756 9150
rect 12820 9148 12826 9212
rect 1393 9074 1459 9077
rect 11697 9074 11763 9077
rect 1393 9072 11763 9074
rect 1393 9016 1398 9072
rect 1454 9016 11702 9072
rect 11758 9016 11763 9072
rect 1393 9014 11763 9016
rect 1393 9011 1459 9014
rect 11697 9011 11763 9014
rect 14365 9074 14431 9077
rect 15840 9074 16000 9104
rect 14365 9072 16000 9074
rect 14365 9016 14370 9072
rect 14426 9016 16000 9072
rect 14365 9014 16000 9016
rect 14365 9011 14431 9014
rect 15840 8984 16000 9014
rect 9673 8938 9739 8941
rect 11237 8938 11303 8941
rect 13353 8938 13419 8941
rect 9673 8936 13419 8938
rect 9673 8880 9678 8936
rect 9734 8880 11242 8936
rect 11298 8880 13358 8936
rect 13414 8880 13419 8936
rect 9673 8878 13419 8880
rect 9673 8875 9739 8878
rect 11237 8875 11303 8878
rect 13353 8875 13419 8878
rect 0 8802 160 8832
rect 9489 8802 9555 8805
rect 10685 8802 10751 8805
rect 0 8742 858 8802
rect 0 8712 160 8742
rect 798 8394 858 8742
rect 9489 8800 10751 8802
rect 9489 8744 9494 8800
rect 9550 8744 10690 8800
rect 10746 8744 10751 8800
rect 9489 8742 10751 8744
rect 9489 8739 9555 8742
rect 10685 8739 10751 8742
rect 11830 8740 11836 8804
rect 11900 8802 11906 8804
rect 12433 8802 12499 8805
rect 11900 8800 12499 8802
rect 11900 8744 12438 8800
rect 12494 8744 12499 8800
rect 11900 8742 12499 8744
rect 11900 8740 11906 8742
rect 12433 8739 12499 8742
rect 15101 8802 15167 8805
rect 15840 8802 16000 8832
rect 15101 8800 16000 8802
rect 15101 8744 15106 8800
rect 15162 8744 16000 8800
rect 15101 8742 16000 8744
rect 15101 8739 15167 8742
rect 4372 8736 4688 8737
rect 4372 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4688 8736
rect 4372 8671 4688 8672
rect 7799 8736 8115 8737
rect 7799 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8115 8736
rect 7799 8671 8115 8672
rect 10133 8530 10199 8533
rect 10688 8530 10748 8739
rect 11226 8736 11542 8737
rect 11226 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11542 8736
rect 11226 8671 11542 8672
rect 14653 8736 14969 8737
rect 14653 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14969 8736
rect 15840 8712 16000 8742
rect 14653 8671 14969 8672
rect 12198 8604 12204 8668
rect 12268 8666 12274 8668
rect 12525 8666 12591 8669
rect 12268 8664 12591 8666
rect 12268 8608 12530 8664
rect 12586 8608 12591 8664
rect 12268 8606 12591 8608
rect 12268 8604 12274 8606
rect 12525 8603 12591 8606
rect 12985 8530 13051 8533
rect 10133 8528 10242 8530
rect 10133 8472 10138 8528
rect 10194 8472 10242 8528
rect 10133 8467 10242 8472
rect 10688 8528 13051 8530
rect 10688 8472 12990 8528
rect 13046 8472 13051 8528
rect 10688 8470 13051 8472
rect 12985 8467 13051 8470
rect 13905 8530 13971 8533
rect 15840 8530 16000 8560
rect 13905 8528 16000 8530
rect 13905 8472 13910 8528
rect 13966 8472 16000 8528
rect 13905 8470 16000 8472
rect 13905 8467 13971 8470
rect 1577 8394 1643 8397
rect 798 8392 1643 8394
rect 798 8336 1582 8392
rect 1638 8336 1643 8392
rect 798 8334 1643 8336
rect 1577 8331 1643 8334
rect 10182 8261 10242 8467
rect 15840 8440 16000 8470
rect 1853 8258 1919 8261
rect 982 8256 1919 8258
rect 982 8200 1858 8256
rect 1914 8200 1919 8256
rect 982 8198 1919 8200
rect 0 7986 160 8016
rect 982 7986 1042 8198
rect 1853 8195 1919 8198
rect 10133 8256 10242 8261
rect 10133 8200 10138 8256
rect 10194 8200 10242 8256
rect 10133 8198 10242 8200
rect 10317 8258 10383 8261
rect 11973 8258 12039 8261
rect 13721 8260 13787 8261
rect 13670 8258 13676 8260
rect 10317 8256 12039 8258
rect 10317 8200 10322 8256
rect 10378 8200 11978 8256
rect 12034 8200 12039 8256
rect 10317 8198 12039 8200
rect 13630 8198 13676 8258
rect 13740 8256 13787 8260
rect 13782 8200 13787 8256
rect 10133 8195 10199 8198
rect 10317 8195 10383 8198
rect 11973 8195 12039 8198
rect 13670 8196 13676 8198
rect 13740 8196 13787 8200
rect 13721 8195 13787 8196
rect 14273 8258 14339 8261
rect 15840 8258 16000 8288
rect 14273 8256 16000 8258
rect 14273 8200 14278 8256
rect 14334 8200 16000 8256
rect 14273 8198 16000 8200
rect 14273 8195 14339 8198
rect 2659 8192 2975 8193
rect 2659 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2975 8192
rect 2659 8127 2975 8128
rect 6086 8192 6402 8193
rect 6086 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6402 8192
rect 6086 8127 6402 8128
rect 9513 8192 9829 8193
rect 9513 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9829 8192
rect 9513 8127 9829 8128
rect 12940 8192 13256 8193
rect 12940 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13256 8192
rect 15840 8168 16000 8198
rect 12940 8127 13256 8128
rect 0 7926 1042 7986
rect 7005 7986 7071 7989
rect 9765 7986 9831 7989
rect 7005 7984 9831 7986
rect 7005 7928 7010 7984
rect 7066 7928 9770 7984
rect 9826 7928 9831 7984
rect 7005 7926 9831 7928
rect 0 7896 160 7926
rect 7005 7923 7071 7926
rect 9765 7923 9831 7926
rect 11237 7986 11303 7989
rect 13353 7986 13419 7989
rect 11237 7984 13419 7986
rect 11237 7928 11242 7984
rect 11298 7928 13358 7984
rect 13414 7928 13419 7984
rect 11237 7926 13419 7928
rect 11237 7923 11303 7926
rect 13353 7923 13419 7926
rect 14273 7986 14339 7989
rect 15840 7986 16000 8016
rect 14273 7984 16000 7986
rect 14273 7928 14278 7984
rect 14334 7928 16000 7984
rect 14273 7926 16000 7928
rect 14273 7923 14339 7926
rect 15840 7896 16000 7926
rect 6545 7850 6611 7853
rect 9581 7850 9647 7853
rect 10593 7852 10659 7853
rect 10542 7850 10548 7852
rect 6545 7848 9647 7850
rect 6545 7792 6550 7848
rect 6606 7792 9586 7848
rect 9642 7792 9647 7848
rect 6545 7790 9647 7792
rect 10502 7790 10548 7850
rect 10612 7848 10659 7852
rect 10654 7792 10659 7848
rect 6545 7787 6611 7790
rect 9581 7787 9647 7790
rect 10542 7788 10548 7790
rect 10612 7788 10659 7792
rect 12566 7788 12572 7852
rect 12636 7850 12642 7852
rect 12893 7850 12959 7853
rect 12636 7848 12959 7850
rect 12636 7792 12898 7848
rect 12954 7792 12959 7848
rect 12636 7790 12959 7792
rect 12636 7788 12642 7790
rect 10593 7787 10659 7788
rect 12893 7787 12959 7790
rect 14181 7850 14247 7853
rect 14181 7848 15210 7850
rect 14181 7792 14186 7848
rect 14242 7792 15210 7848
rect 14181 7790 15210 7792
rect 14181 7787 14247 7790
rect 15150 7714 15210 7790
rect 15840 7714 16000 7744
rect 15150 7654 16000 7714
rect 4372 7648 4688 7649
rect 4372 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4688 7648
rect 4372 7583 4688 7584
rect 7799 7648 8115 7649
rect 7799 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8115 7648
rect 7799 7583 8115 7584
rect 11226 7648 11542 7649
rect 11226 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11542 7648
rect 11226 7583 11542 7584
rect 14653 7648 14969 7649
rect 14653 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14969 7648
rect 15840 7624 16000 7654
rect 14653 7583 14969 7584
rect 14549 7442 14615 7445
rect 15840 7442 16000 7472
rect 14549 7440 16000 7442
rect 14549 7384 14554 7440
rect 14610 7384 16000 7440
rect 14549 7382 16000 7384
rect 14549 7379 14615 7382
rect 15840 7352 16000 7382
rect 0 7170 160 7200
rect 841 7170 907 7173
rect 0 7168 907 7170
rect 0 7112 846 7168
rect 902 7112 907 7168
rect 0 7110 907 7112
rect 0 7080 160 7110
rect 841 7107 907 7110
rect 14273 7170 14339 7173
rect 15840 7170 16000 7200
rect 14273 7168 16000 7170
rect 14273 7112 14278 7168
rect 14334 7112 16000 7168
rect 14273 7110 16000 7112
rect 14273 7107 14339 7110
rect 2659 7104 2975 7105
rect 2659 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2975 7104
rect 2659 7039 2975 7040
rect 6086 7104 6402 7105
rect 6086 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6402 7104
rect 6086 7039 6402 7040
rect 9513 7104 9829 7105
rect 9513 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9829 7104
rect 9513 7039 9829 7040
rect 12940 7104 13256 7105
rect 12940 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13256 7104
rect 15840 7080 16000 7110
rect 12940 7039 13256 7040
rect 5206 6836 5212 6900
rect 5276 6898 5282 6900
rect 12893 6898 12959 6901
rect 13629 6898 13695 6901
rect 5276 6838 12450 6898
rect 5276 6836 5282 6838
rect 12390 6762 12450 6838
rect 12893 6896 13695 6898
rect 12893 6840 12898 6896
rect 12954 6840 13634 6896
rect 13690 6840 13695 6896
rect 12893 6838 13695 6840
rect 12893 6835 12959 6838
rect 13629 6835 13695 6838
rect 15101 6898 15167 6901
rect 15840 6898 16000 6928
rect 15101 6896 16000 6898
rect 15101 6840 15106 6896
rect 15162 6840 16000 6896
rect 15101 6838 16000 6840
rect 15101 6835 15167 6838
rect 15840 6808 16000 6838
rect 13905 6762 13971 6765
rect 12390 6760 13971 6762
rect 12390 6704 13910 6760
rect 13966 6704 13971 6760
rect 12390 6702 13971 6704
rect 13905 6699 13971 6702
rect 15840 6626 16000 6656
rect 15150 6566 16000 6626
rect 4372 6560 4688 6561
rect 4372 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4688 6560
rect 4372 6495 4688 6496
rect 7799 6560 8115 6561
rect 7799 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8115 6560
rect 7799 6495 8115 6496
rect 11226 6560 11542 6561
rect 11226 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11542 6560
rect 11226 6495 11542 6496
rect 14653 6560 14969 6561
rect 14653 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14969 6560
rect 14653 6495 14969 6496
rect 12157 6490 12223 6493
rect 12985 6490 13051 6493
rect 12157 6488 13051 6490
rect 12157 6432 12162 6488
rect 12218 6432 12990 6488
rect 13046 6432 13051 6488
rect 12157 6430 13051 6432
rect 12157 6427 12223 6430
rect 12985 6427 13051 6430
rect 0 6354 160 6384
rect 841 6354 907 6357
rect 0 6352 907 6354
rect 0 6296 846 6352
rect 902 6296 907 6352
rect 0 6294 907 6296
rect 0 6264 160 6294
rect 841 6291 907 6294
rect 8293 6354 8359 6357
rect 13537 6354 13603 6357
rect 8293 6352 13603 6354
rect 8293 6296 8298 6352
rect 8354 6296 13542 6352
rect 13598 6296 13603 6352
rect 8293 6294 13603 6296
rect 8293 6291 8359 6294
rect 13537 6291 13603 6294
rect 13721 6354 13787 6357
rect 15150 6354 15210 6566
rect 15840 6536 16000 6566
rect 15840 6354 16000 6384
rect 13721 6352 15210 6354
rect 13721 6296 13726 6352
rect 13782 6296 15210 6352
rect 13721 6294 15210 6296
rect 15334 6294 16000 6354
rect 13721 6291 13787 6294
rect 3325 6218 3391 6221
rect 14365 6218 14431 6221
rect 3325 6216 14431 6218
rect 3325 6160 3330 6216
rect 3386 6160 14370 6216
rect 14426 6160 14431 6216
rect 3325 6158 14431 6160
rect 3325 6155 3391 6158
rect 14365 6155 14431 6158
rect 15193 6218 15259 6221
rect 15334 6218 15394 6294
rect 15840 6264 16000 6294
rect 15193 6216 15394 6218
rect 15193 6160 15198 6216
rect 15254 6160 15394 6216
rect 15193 6158 15394 6160
rect 15193 6155 15259 6158
rect 11881 6082 11947 6085
rect 11881 6080 12450 6082
rect 11881 6024 11886 6080
rect 11942 6024 12450 6080
rect 11881 6022 12450 6024
rect 11881 6019 11947 6022
rect 2659 6016 2975 6017
rect 2659 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2975 6016
rect 2659 5951 2975 5952
rect 6086 6016 6402 6017
rect 6086 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6402 6016
rect 6086 5951 6402 5952
rect 9513 6016 9829 6017
rect 9513 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9829 6016
rect 9513 5951 9829 5952
rect 11646 5884 11652 5948
rect 11716 5946 11722 5948
rect 11881 5946 11947 5949
rect 11716 5944 11947 5946
rect 11716 5888 11886 5944
rect 11942 5888 11947 5944
rect 11716 5886 11947 5888
rect 11716 5884 11722 5886
rect 11881 5883 11947 5886
rect 12390 5810 12450 6022
rect 12566 6020 12572 6084
rect 12636 6082 12642 6084
rect 12709 6082 12775 6085
rect 15840 6082 16000 6112
rect 12636 6080 12775 6082
rect 12636 6024 12714 6080
rect 12770 6024 12775 6080
rect 12636 6022 12775 6024
rect 12636 6020 12642 6022
rect 12709 6019 12775 6022
rect 14184 6022 16000 6082
rect 12940 6016 13256 6017
rect 12940 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13256 6016
rect 12940 5951 13256 5952
rect 14184 5810 14244 6022
rect 15840 5992 16000 6022
rect 8710 5750 11898 5810
rect 12390 5750 14244 5810
rect 14825 5810 14891 5813
rect 15840 5810 16000 5840
rect 14825 5808 16000 5810
rect 14825 5752 14830 5808
rect 14886 5752 16000 5808
rect 14825 5750 16000 5752
rect 8201 5674 8267 5677
rect 8710 5674 8770 5750
rect 8201 5672 8770 5674
rect 8201 5616 8206 5672
rect 8262 5616 8770 5672
rect 8201 5614 8770 5616
rect 9765 5674 9831 5677
rect 11838 5674 11898 5750
rect 14825 5747 14891 5750
rect 15840 5720 16000 5750
rect 12617 5674 12683 5677
rect 9765 5672 11714 5674
rect 9765 5616 9770 5672
rect 9826 5616 11714 5672
rect 9765 5614 11714 5616
rect 11838 5672 12683 5674
rect 11838 5616 12622 5672
rect 12678 5616 12683 5672
rect 11838 5614 12683 5616
rect 8201 5611 8267 5614
rect 9765 5611 9831 5614
rect 0 5538 160 5568
rect 841 5538 907 5541
rect 0 5536 907 5538
rect 0 5480 846 5536
rect 902 5480 907 5536
rect 0 5478 907 5480
rect 11654 5538 11714 5614
rect 12617 5611 12683 5614
rect 13905 5538 13971 5541
rect 11654 5536 13971 5538
rect 11654 5480 13910 5536
rect 13966 5480 13971 5536
rect 11654 5478 13971 5480
rect 0 5448 160 5478
rect 841 5475 907 5478
rect 13905 5475 13971 5478
rect 14273 5538 14339 5541
rect 15101 5538 15167 5541
rect 15840 5538 16000 5568
rect 14273 5536 14474 5538
rect 14273 5480 14278 5536
rect 14334 5480 14474 5536
rect 14273 5478 14474 5480
rect 14273 5475 14339 5478
rect 4372 5472 4688 5473
rect 4372 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4688 5472
rect 4372 5407 4688 5408
rect 7799 5472 8115 5473
rect 7799 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8115 5472
rect 7799 5407 8115 5408
rect 11226 5472 11542 5473
rect 11226 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11542 5472
rect 11226 5407 11542 5408
rect 10726 5204 10732 5268
rect 10796 5204 10802 5268
rect 10961 5266 11027 5269
rect 13997 5266 14063 5269
rect 10961 5264 14063 5266
rect 10961 5208 10966 5264
rect 11022 5208 14002 5264
rect 14058 5208 14063 5264
rect 10961 5206 14063 5208
rect 14414 5266 14474 5478
rect 15101 5536 16000 5538
rect 15101 5480 15106 5536
rect 15162 5480 16000 5536
rect 15101 5478 16000 5480
rect 15101 5475 15167 5478
rect 14653 5472 14969 5473
rect 14653 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14969 5472
rect 15840 5448 16000 5478
rect 14653 5407 14969 5408
rect 15840 5266 16000 5296
rect 14414 5206 16000 5266
rect 10734 5130 10794 5204
rect 10961 5203 11027 5206
rect 13997 5203 14063 5206
rect 15840 5176 16000 5206
rect 12065 5130 12131 5133
rect 10734 5128 12131 5130
rect 10734 5072 12070 5128
rect 12126 5072 12131 5128
rect 10734 5070 12131 5072
rect 12065 5067 12131 5070
rect 14273 4994 14339 4997
rect 15840 4994 16000 5024
rect 14273 4992 16000 4994
rect 14273 4936 14278 4992
rect 14334 4936 16000 4992
rect 14273 4934 16000 4936
rect 14273 4931 14339 4934
rect 2659 4928 2975 4929
rect 2659 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2975 4928
rect 2659 4863 2975 4864
rect 6086 4928 6402 4929
rect 6086 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6402 4928
rect 6086 4863 6402 4864
rect 9513 4928 9829 4929
rect 9513 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9829 4928
rect 9513 4863 9829 4864
rect 12940 4928 13256 4929
rect 12940 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13256 4928
rect 15840 4904 16000 4934
rect 12940 4863 13256 4864
rect 0 4722 160 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 160 4662
rect 933 4659 999 4662
rect 4372 4384 4688 4385
rect 4372 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4688 4384
rect 4372 4319 4688 4320
rect 7799 4384 8115 4385
rect 7799 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8115 4384
rect 7799 4319 8115 4320
rect 11226 4384 11542 4385
rect 11226 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11542 4384
rect 11226 4319 11542 4320
rect 14653 4384 14969 4385
rect 14653 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14969 4384
rect 14653 4319 14969 4320
rect 8702 3980 8708 4044
rect 8772 4042 8778 4044
rect 14365 4042 14431 4045
rect 8772 4040 14431 4042
rect 8772 3984 14370 4040
rect 14426 3984 14431 4040
rect 8772 3982 14431 3984
rect 8772 3980 8778 3982
rect 14365 3979 14431 3982
rect 0 3906 160 3936
rect 749 3906 815 3909
rect 0 3904 815 3906
rect 0 3848 754 3904
rect 810 3848 815 3904
rect 0 3846 815 3848
rect 0 3816 160 3846
rect 749 3843 815 3846
rect 2659 3840 2975 3841
rect 2659 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2975 3840
rect 2659 3775 2975 3776
rect 6086 3840 6402 3841
rect 6086 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6402 3840
rect 6086 3775 6402 3776
rect 9513 3840 9829 3841
rect 9513 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9829 3840
rect 9513 3775 9829 3776
rect 12940 3840 13256 3841
rect 12940 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13256 3840
rect 12940 3775 13256 3776
rect 4372 3296 4688 3297
rect 4372 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4688 3296
rect 4372 3231 4688 3232
rect 7799 3296 8115 3297
rect 7799 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8115 3296
rect 7799 3231 8115 3232
rect 11226 3296 11542 3297
rect 11226 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11542 3296
rect 11226 3231 11542 3232
rect 14653 3296 14969 3297
rect 14653 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14969 3296
rect 14653 3231 14969 3232
rect 2659 2752 2975 2753
rect 2659 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2975 2752
rect 2659 2687 2975 2688
rect 6086 2752 6402 2753
rect 6086 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6402 2752
rect 6086 2687 6402 2688
rect 9513 2752 9829 2753
rect 9513 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9829 2752
rect 9513 2687 9829 2688
rect 12940 2752 13256 2753
rect 12940 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13256 2752
rect 12940 2687 13256 2688
rect 5809 2684 5875 2685
rect 5758 2682 5764 2684
rect 5718 2622 5764 2682
rect 5828 2680 5875 2684
rect 6637 2684 6703 2685
rect 6637 2682 6684 2684
rect 5870 2624 5875 2680
rect 5758 2620 5764 2622
rect 5828 2620 5875 2624
rect 6592 2680 6684 2682
rect 6592 2624 6642 2680
rect 6592 2622 6684 2624
rect 5809 2619 5875 2620
rect 6637 2620 6684 2622
rect 6748 2620 6754 2684
rect 7414 2620 7420 2684
rect 7484 2682 7490 2684
rect 7649 2682 7715 2685
rect 10869 2684 10935 2685
rect 10869 2682 10916 2684
rect 7484 2680 7715 2682
rect 7484 2624 7654 2680
rect 7710 2624 7715 2680
rect 7484 2622 7715 2624
rect 10824 2680 10916 2682
rect 10824 2624 10874 2680
rect 10824 2622 10916 2624
rect 7484 2620 7490 2622
rect 6637 2619 6703 2620
rect 7649 2619 7715 2622
rect 10869 2620 10916 2622
rect 10980 2620 10986 2684
rect 10869 2619 10935 2620
rect 4372 2208 4688 2209
rect 4372 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4688 2208
rect 4372 2143 4688 2144
rect 7799 2208 8115 2209
rect 7799 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8115 2208
rect 7799 2143 8115 2144
rect 11226 2208 11542 2209
rect 11226 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11542 2208
rect 11226 2143 11542 2144
rect 14653 2208 14969 2209
rect 14653 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14969 2208
rect 14653 2143 14969 2144
rect 5390 1804 5396 1868
rect 5460 1866 5466 1868
rect 11697 1866 11763 1869
rect 5460 1864 11763 1866
rect 5460 1808 11702 1864
rect 11758 1808 11763 1864
rect 5460 1806 11763 1808
rect 5460 1804 5466 1806
rect 11697 1803 11763 1806
rect 2659 1664 2975 1665
rect 2659 1600 2665 1664
rect 2729 1600 2745 1664
rect 2809 1600 2825 1664
rect 2889 1600 2905 1664
rect 2969 1600 2975 1664
rect 2659 1599 2975 1600
rect 6086 1664 6402 1665
rect 6086 1600 6092 1664
rect 6156 1600 6172 1664
rect 6236 1600 6252 1664
rect 6316 1600 6332 1664
rect 6396 1600 6402 1664
rect 6086 1599 6402 1600
rect 9513 1664 9829 1665
rect 9513 1600 9519 1664
rect 9583 1600 9599 1664
rect 9663 1600 9679 1664
rect 9743 1600 9759 1664
rect 9823 1600 9829 1664
rect 9513 1599 9829 1600
rect 12940 1664 13256 1665
rect 12940 1600 12946 1664
rect 13010 1600 13026 1664
rect 13090 1600 13106 1664
rect 13170 1600 13186 1664
rect 13250 1600 13256 1664
rect 12940 1599 13256 1600
rect 4372 1120 4688 1121
rect 4372 1056 4378 1120
rect 4442 1056 4458 1120
rect 4522 1056 4538 1120
rect 4602 1056 4618 1120
rect 4682 1056 4688 1120
rect 4372 1055 4688 1056
rect 7799 1120 8115 1121
rect 7799 1056 7805 1120
rect 7869 1056 7885 1120
rect 7949 1056 7965 1120
rect 8029 1056 8045 1120
rect 8109 1056 8115 1120
rect 7799 1055 8115 1056
rect 11226 1120 11542 1121
rect 11226 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11392 1120
rect 11456 1056 11472 1120
rect 11536 1056 11542 1120
rect 11226 1055 11542 1056
rect 14653 1120 14969 1121
rect 14653 1056 14659 1120
rect 14723 1056 14739 1120
rect 14803 1056 14819 1120
rect 14883 1056 14899 1120
rect 14963 1056 14969 1120
rect 14653 1055 14969 1056
<< via3 >>
rect 4378 43548 4442 43552
rect 4378 43492 4382 43548
rect 4382 43492 4438 43548
rect 4438 43492 4442 43548
rect 4378 43488 4442 43492
rect 4458 43548 4522 43552
rect 4458 43492 4462 43548
rect 4462 43492 4518 43548
rect 4518 43492 4522 43548
rect 4458 43488 4522 43492
rect 4538 43548 4602 43552
rect 4538 43492 4542 43548
rect 4542 43492 4598 43548
rect 4598 43492 4602 43548
rect 4538 43488 4602 43492
rect 4618 43548 4682 43552
rect 4618 43492 4622 43548
rect 4622 43492 4678 43548
rect 4678 43492 4682 43548
rect 4618 43488 4682 43492
rect 7805 43548 7869 43552
rect 7805 43492 7809 43548
rect 7809 43492 7865 43548
rect 7865 43492 7869 43548
rect 7805 43488 7869 43492
rect 7885 43548 7949 43552
rect 7885 43492 7889 43548
rect 7889 43492 7945 43548
rect 7945 43492 7949 43548
rect 7885 43488 7949 43492
rect 7965 43548 8029 43552
rect 7965 43492 7969 43548
rect 7969 43492 8025 43548
rect 8025 43492 8029 43548
rect 7965 43488 8029 43492
rect 8045 43548 8109 43552
rect 8045 43492 8049 43548
rect 8049 43492 8105 43548
rect 8105 43492 8109 43548
rect 8045 43488 8109 43492
rect 11232 43548 11296 43552
rect 11232 43492 11236 43548
rect 11236 43492 11292 43548
rect 11292 43492 11296 43548
rect 11232 43488 11296 43492
rect 11312 43548 11376 43552
rect 11312 43492 11316 43548
rect 11316 43492 11372 43548
rect 11372 43492 11376 43548
rect 11312 43488 11376 43492
rect 11392 43548 11456 43552
rect 11392 43492 11396 43548
rect 11396 43492 11452 43548
rect 11452 43492 11456 43548
rect 11392 43488 11456 43492
rect 11472 43548 11536 43552
rect 11472 43492 11476 43548
rect 11476 43492 11532 43548
rect 11532 43492 11536 43548
rect 11472 43488 11536 43492
rect 14659 43548 14723 43552
rect 14659 43492 14663 43548
rect 14663 43492 14719 43548
rect 14719 43492 14723 43548
rect 14659 43488 14723 43492
rect 14739 43548 14803 43552
rect 14739 43492 14743 43548
rect 14743 43492 14799 43548
rect 14799 43492 14803 43548
rect 14739 43488 14803 43492
rect 14819 43548 14883 43552
rect 14819 43492 14823 43548
rect 14823 43492 14879 43548
rect 14879 43492 14883 43548
rect 14819 43488 14883 43492
rect 14899 43548 14963 43552
rect 14899 43492 14903 43548
rect 14903 43492 14959 43548
rect 14959 43492 14963 43548
rect 14899 43488 14963 43492
rect 2665 43004 2729 43008
rect 2665 42948 2669 43004
rect 2669 42948 2725 43004
rect 2725 42948 2729 43004
rect 2665 42944 2729 42948
rect 2745 43004 2809 43008
rect 2745 42948 2749 43004
rect 2749 42948 2805 43004
rect 2805 42948 2809 43004
rect 2745 42944 2809 42948
rect 2825 43004 2889 43008
rect 2825 42948 2829 43004
rect 2829 42948 2885 43004
rect 2885 42948 2889 43004
rect 2825 42944 2889 42948
rect 2905 43004 2969 43008
rect 2905 42948 2909 43004
rect 2909 42948 2965 43004
rect 2965 42948 2969 43004
rect 2905 42944 2969 42948
rect 6092 43004 6156 43008
rect 6092 42948 6096 43004
rect 6096 42948 6152 43004
rect 6152 42948 6156 43004
rect 6092 42944 6156 42948
rect 6172 43004 6236 43008
rect 6172 42948 6176 43004
rect 6176 42948 6232 43004
rect 6232 42948 6236 43004
rect 6172 42944 6236 42948
rect 6252 43004 6316 43008
rect 6252 42948 6256 43004
rect 6256 42948 6312 43004
rect 6312 42948 6316 43004
rect 6252 42944 6316 42948
rect 6332 43004 6396 43008
rect 6332 42948 6336 43004
rect 6336 42948 6392 43004
rect 6392 42948 6396 43004
rect 6332 42944 6396 42948
rect 9519 43004 9583 43008
rect 9519 42948 9523 43004
rect 9523 42948 9579 43004
rect 9579 42948 9583 43004
rect 9519 42944 9583 42948
rect 9599 43004 9663 43008
rect 9599 42948 9603 43004
rect 9603 42948 9659 43004
rect 9659 42948 9663 43004
rect 9599 42944 9663 42948
rect 9679 43004 9743 43008
rect 9679 42948 9683 43004
rect 9683 42948 9739 43004
rect 9739 42948 9743 43004
rect 9679 42944 9743 42948
rect 9759 43004 9823 43008
rect 9759 42948 9763 43004
rect 9763 42948 9819 43004
rect 9819 42948 9823 43004
rect 9759 42944 9823 42948
rect 12946 43004 13010 43008
rect 12946 42948 12950 43004
rect 12950 42948 13006 43004
rect 13006 42948 13010 43004
rect 12946 42944 13010 42948
rect 13026 43004 13090 43008
rect 13026 42948 13030 43004
rect 13030 42948 13086 43004
rect 13086 42948 13090 43004
rect 13026 42944 13090 42948
rect 13106 43004 13170 43008
rect 13106 42948 13110 43004
rect 13110 42948 13166 43004
rect 13166 42948 13170 43004
rect 13106 42944 13170 42948
rect 13186 43004 13250 43008
rect 13186 42948 13190 43004
rect 13190 42948 13246 43004
rect 13246 42948 13250 43004
rect 13186 42944 13250 42948
rect 4378 42460 4442 42464
rect 4378 42404 4382 42460
rect 4382 42404 4438 42460
rect 4438 42404 4442 42460
rect 4378 42400 4442 42404
rect 4458 42460 4522 42464
rect 4458 42404 4462 42460
rect 4462 42404 4518 42460
rect 4518 42404 4522 42460
rect 4458 42400 4522 42404
rect 4538 42460 4602 42464
rect 4538 42404 4542 42460
rect 4542 42404 4598 42460
rect 4598 42404 4602 42460
rect 4538 42400 4602 42404
rect 4618 42460 4682 42464
rect 4618 42404 4622 42460
rect 4622 42404 4678 42460
rect 4678 42404 4682 42460
rect 4618 42400 4682 42404
rect 7805 42460 7869 42464
rect 7805 42404 7809 42460
rect 7809 42404 7865 42460
rect 7865 42404 7869 42460
rect 7805 42400 7869 42404
rect 7885 42460 7949 42464
rect 7885 42404 7889 42460
rect 7889 42404 7945 42460
rect 7945 42404 7949 42460
rect 7885 42400 7949 42404
rect 7965 42460 8029 42464
rect 7965 42404 7969 42460
rect 7969 42404 8025 42460
rect 8025 42404 8029 42460
rect 7965 42400 8029 42404
rect 8045 42460 8109 42464
rect 8045 42404 8049 42460
rect 8049 42404 8105 42460
rect 8105 42404 8109 42460
rect 8045 42400 8109 42404
rect 11232 42460 11296 42464
rect 11232 42404 11236 42460
rect 11236 42404 11292 42460
rect 11292 42404 11296 42460
rect 11232 42400 11296 42404
rect 11312 42460 11376 42464
rect 11312 42404 11316 42460
rect 11316 42404 11372 42460
rect 11372 42404 11376 42460
rect 11312 42400 11376 42404
rect 11392 42460 11456 42464
rect 11392 42404 11396 42460
rect 11396 42404 11452 42460
rect 11452 42404 11456 42460
rect 11392 42400 11456 42404
rect 11472 42460 11536 42464
rect 11472 42404 11476 42460
rect 11476 42404 11532 42460
rect 11532 42404 11536 42460
rect 11472 42400 11536 42404
rect 14659 42460 14723 42464
rect 14659 42404 14663 42460
rect 14663 42404 14719 42460
rect 14719 42404 14723 42460
rect 14659 42400 14723 42404
rect 14739 42460 14803 42464
rect 14739 42404 14743 42460
rect 14743 42404 14799 42460
rect 14799 42404 14803 42460
rect 14739 42400 14803 42404
rect 14819 42460 14883 42464
rect 14819 42404 14823 42460
rect 14823 42404 14879 42460
rect 14879 42404 14883 42460
rect 14819 42400 14883 42404
rect 14899 42460 14963 42464
rect 14899 42404 14903 42460
rect 14903 42404 14959 42460
rect 14959 42404 14963 42460
rect 14899 42400 14963 42404
rect 5396 42060 5460 42124
rect 2665 41916 2729 41920
rect 2665 41860 2669 41916
rect 2669 41860 2725 41916
rect 2725 41860 2729 41916
rect 2665 41856 2729 41860
rect 2745 41916 2809 41920
rect 2745 41860 2749 41916
rect 2749 41860 2805 41916
rect 2805 41860 2809 41916
rect 2745 41856 2809 41860
rect 2825 41916 2889 41920
rect 2825 41860 2829 41916
rect 2829 41860 2885 41916
rect 2885 41860 2889 41916
rect 2825 41856 2889 41860
rect 2905 41916 2969 41920
rect 2905 41860 2909 41916
rect 2909 41860 2965 41916
rect 2965 41860 2969 41916
rect 2905 41856 2969 41860
rect 6092 41916 6156 41920
rect 6092 41860 6096 41916
rect 6096 41860 6152 41916
rect 6152 41860 6156 41916
rect 6092 41856 6156 41860
rect 6172 41916 6236 41920
rect 6172 41860 6176 41916
rect 6176 41860 6232 41916
rect 6232 41860 6236 41916
rect 6172 41856 6236 41860
rect 6252 41916 6316 41920
rect 6252 41860 6256 41916
rect 6256 41860 6312 41916
rect 6312 41860 6316 41916
rect 6252 41856 6316 41860
rect 6332 41916 6396 41920
rect 6332 41860 6336 41916
rect 6336 41860 6392 41916
rect 6392 41860 6396 41916
rect 6332 41856 6396 41860
rect 9519 41916 9583 41920
rect 9519 41860 9523 41916
rect 9523 41860 9579 41916
rect 9579 41860 9583 41916
rect 9519 41856 9583 41860
rect 9599 41916 9663 41920
rect 9599 41860 9603 41916
rect 9603 41860 9659 41916
rect 9659 41860 9663 41916
rect 9599 41856 9663 41860
rect 9679 41916 9743 41920
rect 9679 41860 9683 41916
rect 9683 41860 9739 41916
rect 9739 41860 9743 41916
rect 9679 41856 9743 41860
rect 9759 41916 9823 41920
rect 9759 41860 9763 41916
rect 9763 41860 9819 41916
rect 9819 41860 9823 41916
rect 9759 41856 9823 41860
rect 12946 41916 13010 41920
rect 12946 41860 12950 41916
rect 12950 41860 13006 41916
rect 13006 41860 13010 41916
rect 12946 41856 13010 41860
rect 13026 41916 13090 41920
rect 13026 41860 13030 41916
rect 13030 41860 13086 41916
rect 13086 41860 13090 41916
rect 13026 41856 13090 41860
rect 13106 41916 13170 41920
rect 13106 41860 13110 41916
rect 13110 41860 13166 41916
rect 13166 41860 13170 41916
rect 13106 41856 13170 41860
rect 13186 41916 13250 41920
rect 13186 41860 13190 41916
rect 13190 41860 13246 41916
rect 13246 41860 13250 41916
rect 13186 41856 13250 41860
rect 5764 41848 5828 41852
rect 5764 41792 5778 41848
rect 5778 41792 5828 41848
rect 5764 41788 5828 41792
rect 6684 41788 6748 41852
rect 7420 41788 7484 41852
rect 10916 41848 10980 41852
rect 10916 41792 10966 41848
rect 10966 41792 10980 41848
rect 10916 41788 10980 41792
rect 3924 41516 3988 41580
rect 10732 41516 10796 41580
rect 4378 41372 4442 41376
rect 4378 41316 4382 41372
rect 4382 41316 4438 41372
rect 4438 41316 4442 41372
rect 4378 41312 4442 41316
rect 4458 41372 4522 41376
rect 4458 41316 4462 41372
rect 4462 41316 4518 41372
rect 4518 41316 4522 41372
rect 4458 41312 4522 41316
rect 4538 41372 4602 41376
rect 4538 41316 4542 41372
rect 4542 41316 4598 41372
rect 4598 41316 4602 41372
rect 4538 41312 4602 41316
rect 4618 41372 4682 41376
rect 4618 41316 4622 41372
rect 4622 41316 4678 41372
rect 4678 41316 4682 41372
rect 4618 41312 4682 41316
rect 7805 41372 7869 41376
rect 7805 41316 7809 41372
rect 7809 41316 7865 41372
rect 7865 41316 7869 41372
rect 7805 41312 7869 41316
rect 7885 41372 7949 41376
rect 7885 41316 7889 41372
rect 7889 41316 7945 41372
rect 7945 41316 7949 41372
rect 7885 41312 7949 41316
rect 7965 41372 8029 41376
rect 7965 41316 7969 41372
rect 7969 41316 8025 41372
rect 8025 41316 8029 41372
rect 7965 41312 8029 41316
rect 8045 41372 8109 41376
rect 8045 41316 8049 41372
rect 8049 41316 8105 41372
rect 8105 41316 8109 41372
rect 8045 41312 8109 41316
rect 11232 41372 11296 41376
rect 11232 41316 11236 41372
rect 11236 41316 11292 41372
rect 11292 41316 11296 41372
rect 11232 41312 11296 41316
rect 11312 41372 11376 41376
rect 11312 41316 11316 41372
rect 11316 41316 11372 41372
rect 11372 41316 11376 41372
rect 11312 41312 11376 41316
rect 11392 41372 11456 41376
rect 11392 41316 11396 41372
rect 11396 41316 11452 41372
rect 11452 41316 11456 41372
rect 11392 41312 11456 41316
rect 11472 41372 11536 41376
rect 11472 41316 11476 41372
rect 11476 41316 11532 41372
rect 11532 41316 11536 41372
rect 11472 41312 11536 41316
rect 14659 41372 14723 41376
rect 14659 41316 14663 41372
rect 14663 41316 14719 41372
rect 14719 41316 14723 41372
rect 14659 41312 14723 41316
rect 14739 41372 14803 41376
rect 14739 41316 14743 41372
rect 14743 41316 14799 41372
rect 14799 41316 14803 41372
rect 14739 41312 14803 41316
rect 14819 41372 14883 41376
rect 14819 41316 14823 41372
rect 14823 41316 14879 41372
rect 14879 41316 14883 41372
rect 14819 41312 14883 41316
rect 14899 41372 14963 41376
rect 14899 41316 14903 41372
rect 14903 41316 14959 41372
rect 14959 41316 14963 41372
rect 14899 41312 14963 41316
rect 2665 40828 2729 40832
rect 2665 40772 2669 40828
rect 2669 40772 2725 40828
rect 2725 40772 2729 40828
rect 2665 40768 2729 40772
rect 2745 40828 2809 40832
rect 2745 40772 2749 40828
rect 2749 40772 2805 40828
rect 2805 40772 2809 40828
rect 2745 40768 2809 40772
rect 2825 40828 2889 40832
rect 2825 40772 2829 40828
rect 2829 40772 2885 40828
rect 2885 40772 2889 40828
rect 2825 40768 2889 40772
rect 2905 40828 2969 40832
rect 2905 40772 2909 40828
rect 2909 40772 2965 40828
rect 2965 40772 2969 40828
rect 2905 40768 2969 40772
rect 6092 40828 6156 40832
rect 6092 40772 6096 40828
rect 6096 40772 6152 40828
rect 6152 40772 6156 40828
rect 6092 40768 6156 40772
rect 6172 40828 6236 40832
rect 6172 40772 6176 40828
rect 6176 40772 6232 40828
rect 6232 40772 6236 40828
rect 6172 40768 6236 40772
rect 6252 40828 6316 40832
rect 6252 40772 6256 40828
rect 6256 40772 6312 40828
rect 6312 40772 6316 40828
rect 6252 40768 6316 40772
rect 6332 40828 6396 40832
rect 6332 40772 6336 40828
rect 6336 40772 6392 40828
rect 6392 40772 6396 40828
rect 6332 40768 6396 40772
rect 9519 40828 9583 40832
rect 9519 40772 9523 40828
rect 9523 40772 9579 40828
rect 9579 40772 9583 40828
rect 9519 40768 9583 40772
rect 9599 40828 9663 40832
rect 9599 40772 9603 40828
rect 9603 40772 9659 40828
rect 9659 40772 9663 40828
rect 9599 40768 9663 40772
rect 9679 40828 9743 40832
rect 9679 40772 9683 40828
rect 9683 40772 9739 40828
rect 9739 40772 9743 40828
rect 9679 40768 9743 40772
rect 9759 40828 9823 40832
rect 9759 40772 9763 40828
rect 9763 40772 9819 40828
rect 9819 40772 9823 40828
rect 9759 40768 9823 40772
rect 12946 40828 13010 40832
rect 12946 40772 12950 40828
rect 12950 40772 13006 40828
rect 13006 40772 13010 40828
rect 12946 40768 13010 40772
rect 13026 40828 13090 40832
rect 13026 40772 13030 40828
rect 13030 40772 13086 40828
rect 13086 40772 13090 40828
rect 13026 40768 13090 40772
rect 13106 40828 13170 40832
rect 13106 40772 13110 40828
rect 13110 40772 13166 40828
rect 13166 40772 13170 40828
rect 13106 40768 13170 40772
rect 13186 40828 13250 40832
rect 13186 40772 13190 40828
rect 13190 40772 13246 40828
rect 13246 40772 13250 40828
rect 13186 40768 13250 40772
rect 4378 40284 4442 40288
rect 4378 40228 4382 40284
rect 4382 40228 4438 40284
rect 4438 40228 4442 40284
rect 4378 40224 4442 40228
rect 4458 40284 4522 40288
rect 4458 40228 4462 40284
rect 4462 40228 4518 40284
rect 4518 40228 4522 40284
rect 4458 40224 4522 40228
rect 4538 40284 4602 40288
rect 4538 40228 4542 40284
rect 4542 40228 4598 40284
rect 4598 40228 4602 40284
rect 4538 40224 4602 40228
rect 4618 40284 4682 40288
rect 4618 40228 4622 40284
rect 4622 40228 4678 40284
rect 4678 40228 4682 40284
rect 4618 40224 4682 40228
rect 7805 40284 7869 40288
rect 7805 40228 7809 40284
rect 7809 40228 7865 40284
rect 7865 40228 7869 40284
rect 7805 40224 7869 40228
rect 7885 40284 7949 40288
rect 7885 40228 7889 40284
rect 7889 40228 7945 40284
rect 7945 40228 7949 40284
rect 7885 40224 7949 40228
rect 7965 40284 8029 40288
rect 7965 40228 7969 40284
rect 7969 40228 8025 40284
rect 8025 40228 8029 40284
rect 7965 40224 8029 40228
rect 8045 40284 8109 40288
rect 8045 40228 8049 40284
rect 8049 40228 8105 40284
rect 8105 40228 8109 40284
rect 8045 40224 8109 40228
rect 11232 40284 11296 40288
rect 11232 40228 11236 40284
rect 11236 40228 11292 40284
rect 11292 40228 11296 40284
rect 11232 40224 11296 40228
rect 11312 40284 11376 40288
rect 11312 40228 11316 40284
rect 11316 40228 11372 40284
rect 11372 40228 11376 40284
rect 11312 40224 11376 40228
rect 11392 40284 11456 40288
rect 11392 40228 11396 40284
rect 11396 40228 11452 40284
rect 11452 40228 11456 40284
rect 11392 40224 11456 40228
rect 11472 40284 11536 40288
rect 11472 40228 11476 40284
rect 11476 40228 11532 40284
rect 11532 40228 11536 40284
rect 11472 40224 11536 40228
rect 14659 40284 14723 40288
rect 14659 40228 14663 40284
rect 14663 40228 14719 40284
rect 14719 40228 14723 40284
rect 14659 40224 14723 40228
rect 14739 40284 14803 40288
rect 14739 40228 14743 40284
rect 14743 40228 14799 40284
rect 14799 40228 14803 40284
rect 14739 40224 14803 40228
rect 14819 40284 14883 40288
rect 14819 40228 14823 40284
rect 14823 40228 14879 40284
rect 14879 40228 14883 40284
rect 14819 40224 14883 40228
rect 14899 40284 14963 40288
rect 14899 40228 14903 40284
rect 14903 40228 14959 40284
rect 14959 40228 14963 40284
rect 14899 40224 14963 40228
rect 2665 39740 2729 39744
rect 2665 39684 2669 39740
rect 2669 39684 2725 39740
rect 2725 39684 2729 39740
rect 2665 39680 2729 39684
rect 2745 39740 2809 39744
rect 2745 39684 2749 39740
rect 2749 39684 2805 39740
rect 2805 39684 2809 39740
rect 2745 39680 2809 39684
rect 2825 39740 2889 39744
rect 2825 39684 2829 39740
rect 2829 39684 2885 39740
rect 2885 39684 2889 39740
rect 2825 39680 2889 39684
rect 2905 39740 2969 39744
rect 2905 39684 2909 39740
rect 2909 39684 2965 39740
rect 2965 39684 2969 39740
rect 2905 39680 2969 39684
rect 6092 39740 6156 39744
rect 6092 39684 6096 39740
rect 6096 39684 6152 39740
rect 6152 39684 6156 39740
rect 6092 39680 6156 39684
rect 6172 39740 6236 39744
rect 6172 39684 6176 39740
rect 6176 39684 6232 39740
rect 6232 39684 6236 39740
rect 6172 39680 6236 39684
rect 6252 39740 6316 39744
rect 6252 39684 6256 39740
rect 6256 39684 6312 39740
rect 6312 39684 6316 39740
rect 6252 39680 6316 39684
rect 6332 39740 6396 39744
rect 6332 39684 6336 39740
rect 6336 39684 6392 39740
rect 6392 39684 6396 39740
rect 6332 39680 6396 39684
rect 9519 39740 9583 39744
rect 9519 39684 9523 39740
rect 9523 39684 9579 39740
rect 9579 39684 9583 39740
rect 9519 39680 9583 39684
rect 9599 39740 9663 39744
rect 9599 39684 9603 39740
rect 9603 39684 9659 39740
rect 9659 39684 9663 39740
rect 9599 39680 9663 39684
rect 9679 39740 9743 39744
rect 9679 39684 9683 39740
rect 9683 39684 9739 39740
rect 9739 39684 9743 39740
rect 9679 39680 9743 39684
rect 9759 39740 9823 39744
rect 9759 39684 9763 39740
rect 9763 39684 9819 39740
rect 9819 39684 9823 39740
rect 9759 39680 9823 39684
rect 12946 39740 13010 39744
rect 12946 39684 12950 39740
rect 12950 39684 13006 39740
rect 13006 39684 13010 39740
rect 12946 39680 13010 39684
rect 13026 39740 13090 39744
rect 13026 39684 13030 39740
rect 13030 39684 13086 39740
rect 13086 39684 13090 39740
rect 13026 39680 13090 39684
rect 13106 39740 13170 39744
rect 13106 39684 13110 39740
rect 13110 39684 13166 39740
rect 13166 39684 13170 39740
rect 13106 39680 13170 39684
rect 13186 39740 13250 39744
rect 13186 39684 13190 39740
rect 13190 39684 13246 39740
rect 13246 39684 13250 39740
rect 13186 39680 13250 39684
rect 4378 39196 4442 39200
rect 4378 39140 4382 39196
rect 4382 39140 4438 39196
rect 4438 39140 4442 39196
rect 4378 39136 4442 39140
rect 4458 39196 4522 39200
rect 4458 39140 4462 39196
rect 4462 39140 4518 39196
rect 4518 39140 4522 39196
rect 4458 39136 4522 39140
rect 4538 39196 4602 39200
rect 4538 39140 4542 39196
rect 4542 39140 4598 39196
rect 4598 39140 4602 39196
rect 4538 39136 4602 39140
rect 4618 39196 4682 39200
rect 4618 39140 4622 39196
rect 4622 39140 4678 39196
rect 4678 39140 4682 39196
rect 4618 39136 4682 39140
rect 7805 39196 7869 39200
rect 7805 39140 7809 39196
rect 7809 39140 7865 39196
rect 7865 39140 7869 39196
rect 7805 39136 7869 39140
rect 7885 39196 7949 39200
rect 7885 39140 7889 39196
rect 7889 39140 7945 39196
rect 7945 39140 7949 39196
rect 7885 39136 7949 39140
rect 7965 39196 8029 39200
rect 7965 39140 7969 39196
rect 7969 39140 8025 39196
rect 8025 39140 8029 39196
rect 7965 39136 8029 39140
rect 8045 39196 8109 39200
rect 8045 39140 8049 39196
rect 8049 39140 8105 39196
rect 8105 39140 8109 39196
rect 8045 39136 8109 39140
rect 11232 39196 11296 39200
rect 11232 39140 11236 39196
rect 11236 39140 11292 39196
rect 11292 39140 11296 39196
rect 11232 39136 11296 39140
rect 11312 39196 11376 39200
rect 11312 39140 11316 39196
rect 11316 39140 11372 39196
rect 11372 39140 11376 39196
rect 11312 39136 11376 39140
rect 11392 39196 11456 39200
rect 11392 39140 11396 39196
rect 11396 39140 11452 39196
rect 11452 39140 11456 39196
rect 11392 39136 11456 39140
rect 11472 39196 11536 39200
rect 11472 39140 11476 39196
rect 11476 39140 11532 39196
rect 11532 39140 11536 39196
rect 11472 39136 11536 39140
rect 14659 39196 14723 39200
rect 14659 39140 14663 39196
rect 14663 39140 14719 39196
rect 14719 39140 14723 39196
rect 14659 39136 14723 39140
rect 14739 39196 14803 39200
rect 14739 39140 14743 39196
rect 14743 39140 14799 39196
rect 14799 39140 14803 39196
rect 14739 39136 14803 39140
rect 14819 39196 14883 39200
rect 14819 39140 14823 39196
rect 14823 39140 14879 39196
rect 14879 39140 14883 39196
rect 14819 39136 14883 39140
rect 14899 39196 14963 39200
rect 14899 39140 14903 39196
rect 14903 39140 14959 39196
rect 14959 39140 14963 39196
rect 14899 39136 14963 39140
rect 2665 38652 2729 38656
rect 2665 38596 2669 38652
rect 2669 38596 2725 38652
rect 2725 38596 2729 38652
rect 2665 38592 2729 38596
rect 2745 38652 2809 38656
rect 2745 38596 2749 38652
rect 2749 38596 2805 38652
rect 2805 38596 2809 38652
rect 2745 38592 2809 38596
rect 2825 38652 2889 38656
rect 2825 38596 2829 38652
rect 2829 38596 2885 38652
rect 2885 38596 2889 38652
rect 2825 38592 2889 38596
rect 2905 38652 2969 38656
rect 2905 38596 2909 38652
rect 2909 38596 2965 38652
rect 2965 38596 2969 38652
rect 2905 38592 2969 38596
rect 6092 38652 6156 38656
rect 6092 38596 6096 38652
rect 6096 38596 6152 38652
rect 6152 38596 6156 38652
rect 6092 38592 6156 38596
rect 6172 38652 6236 38656
rect 6172 38596 6176 38652
rect 6176 38596 6232 38652
rect 6232 38596 6236 38652
rect 6172 38592 6236 38596
rect 6252 38652 6316 38656
rect 6252 38596 6256 38652
rect 6256 38596 6312 38652
rect 6312 38596 6316 38652
rect 6252 38592 6316 38596
rect 6332 38652 6396 38656
rect 6332 38596 6336 38652
rect 6336 38596 6392 38652
rect 6392 38596 6396 38652
rect 6332 38592 6396 38596
rect 9519 38652 9583 38656
rect 9519 38596 9523 38652
rect 9523 38596 9579 38652
rect 9579 38596 9583 38652
rect 9519 38592 9583 38596
rect 9599 38652 9663 38656
rect 9599 38596 9603 38652
rect 9603 38596 9659 38652
rect 9659 38596 9663 38652
rect 9599 38592 9663 38596
rect 9679 38652 9743 38656
rect 9679 38596 9683 38652
rect 9683 38596 9739 38652
rect 9739 38596 9743 38652
rect 9679 38592 9743 38596
rect 9759 38652 9823 38656
rect 9759 38596 9763 38652
rect 9763 38596 9819 38652
rect 9819 38596 9823 38652
rect 9759 38592 9823 38596
rect 12946 38652 13010 38656
rect 12946 38596 12950 38652
rect 12950 38596 13006 38652
rect 13006 38596 13010 38652
rect 12946 38592 13010 38596
rect 13026 38652 13090 38656
rect 13026 38596 13030 38652
rect 13030 38596 13086 38652
rect 13086 38596 13090 38652
rect 13026 38592 13090 38596
rect 13106 38652 13170 38656
rect 13106 38596 13110 38652
rect 13110 38596 13166 38652
rect 13166 38596 13170 38652
rect 13106 38592 13170 38596
rect 13186 38652 13250 38656
rect 13186 38596 13190 38652
rect 13190 38596 13246 38652
rect 13246 38596 13250 38652
rect 13186 38592 13250 38596
rect 4378 38108 4442 38112
rect 4378 38052 4382 38108
rect 4382 38052 4438 38108
rect 4438 38052 4442 38108
rect 4378 38048 4442 38052
rect 4458 38108 4522 38112
rect 4458 38052 4462 38108
rect 4462 38052 4518 38108
rect 4518 38052 4522 38108
rect 4458 38048 4522 38052
rect 4538 38108 4602 38112
rect 4538 38052 4542 38108
rect 4542 38052 4598 38108
rect 4598 38052 4602 38108
rect 4538 38048 4602 38052
rect 4618 38108 4682 38112
rect 4618 38052 4622 38108
rect 4622 38052 4678 38108
rect 4678 38052 4682 38108
rect 4618 38048 4682 38052
rect 7805 38108 7869 38112
rect 7805 38052 7809 38108
rect 7809 38052 7865 38108
rect 7865 38052 7869 38108
rect 7805 38048 7869 38052
rect 7885 38108 7949 38112
rect 7885 38052 7889 38108
rect 7889 38052 7945 38108
rect 7945 38052 7949 38108
rect 7885 38048 7949 38052
rect 7965 38108 8029 38112
rect 7965 38052 7969 38108
rect 7969 38052 8025 38108
rect 8025 38052 8029 38108
rect 7965 38048 8029 38052
rect 8045 38108 8109 38112
rect 8045 38052 8049 38108
rect 8049 38052 8105 38108
rect 8105 38052 8109 38108
rect 8045 38048 8109 38052
rect 11232 38108 11296 38112
rect 11232 38052 11236 38108
rect 11236 38052 11292 38108
rect 11292 38052 11296 38108
rect 11232 38048 11296 38052
rect 11312 38108 11376 38112
rect 11312 38052 11316 38108
rect 11316 38052 11372 38108
rect 11372 38052 11376 38108
rect 11312 38048 11376 38052
rect 11392 38108 11456 38112
rect 11392 38052 11396 38108
rect 11396 38052 11452 38108
rect 11452 38052 11456 38108
rect 11392 38048 11456 38052
rect 11472 38108 11536 38112
rect 11472 38052 11476 38108
rect 11476 38052 11532 38108
rect 11532 38052 11536 38108
rect 11472 38048 11536 38052
rect 14659 38108 14723 38112
rect 14659 38052 14663 38108
rect 14663 38052 14719 38108
rect 14719 38052 14723 38108
rect 14659 38048 14723 38052
rect 14739 38108 14803 38112
rect 14739 38052 14743 38108
rect 14743 38052 14799 38108
rect 14799 38052 14803 38108
rect 14739 38048 14803 38052
rect 14819 38108 14883 38112
rect 14819 38052 14823 38108
rect 14823 38052 14879 38108
rect 14879 38052 14883 38108
rect 14819 38048 14883 38052
rect 14899 38108 14963 38112
rect 14899 38052 14903 38108
rect 14903 38052 14959 38108
rect 14959 38052 14963 38108
rect 14899 38048 14963 38052
rect 2665 37564 2729 37568
rect 2665 37508 2669 37564
rect 2669 37508 2725 37564
rect 2725 37508 2729 37564
rect 2665 37504 2729 37508
rect 2745 37564 2809 37568
rect 2745 37508 2749 37564
rect 2749 37508 2805 37564
rect 2805 37508 2809 37564
rect 2745 37504 2809 37508
rect 2825 37564 2889 37568
rect 2825 37508 2829 37564
rect 2829 37508 2885 37564
rect 2885 37508 2889 37564
rect 2825 37504 2889 37508
rect 2905 37564 2969 37568
rect 2905 37508 2909 37564
rect 2909 37508 2965 37564
rect 2965 37508 2969 37564
rect 2905 37504 2969 37508
rect 6092 37564 6156 37568
rect 6092 37508 6096 37564
rect 6096 37508 6152 37564
rect 6152 37508 6156 37564
rect 6092 37504 6156 37508
rect 6172 37564 6236 37568
rect 6172 37508 6176 37564
rect 6176 37508 6232 37564
rect 6232 37508 6236 37564
rect 6172 37504 6236 37508
rect 6252 37564 6316 37568
rect 6252 37508 6256 37564
rect 6256 37508 6312 37564
rect 6312 37508 6316 37564
rect 6252 37504 6316 37508
rect 6332 37564 6396 37568
rect 6332 37508 6336 37564
rect 6336 37508 6392 37564
rect 6392 37508 6396 37564
rect 6332 37504 6396 37508
rect 9519 37564 9583 37568
rect 9519 37508 9523 37564
rect 9523 37508 9579 37564
rect 9579 37508 9583 37564
rect 9519 37504 9583 37508
rect 9599 37564 9663 37568
rect 9599 37508 9603 37564
rect 9603 37508 9659 37564
rect 9659 37508 9663 37564
rect 9599 37504 9663 37508
rect 9679 37564 9743 37568
rect 9679 37508 9683 37564
rect 9683 37508 9739 37564
rect 9739 37508 9743 37564
rect 9679 37504 9743 37508
rect 9759 37564 9823 37568
rect 9759 37508 9763 37564
rect 9763 37508 9819 37564
rect 9819 37508 9823 37564
rect 9759 37504 9823 37508
rect 12946 37564 13010 37568
rect 12946 37508 12950 37564
rect 12950 37508 13006 37564
rect 13006 37508 13010 37564
rect 12946 37504 13010 37508
rect 13026 37564 13090 37568
rect 13026 37508 13030 37564
rect 13030 37508 13086 37564
rect 13086 37508 13090 37564
rect 13026 37504 13090 37508
rect 13106 37564 13170 37568
rect 13106 37508 13110 37564
rect 13110 37508 13166 37564
rect 13166 37508 13170 37564
rect 13106 37504 13170 37508
rect 13186 37564 13250 37568
rect 13186 37508 13190 37564
rect 13190 37508 13246 37564
rect 13246 37508 13250 37564
rect 13186 37504 13250 37508
rect 4378 37020 4442 37024
rect 4378 36964 4382 37020
rect 4382 36964 4438 37020
rect 4438 36964 4442 37020
rect 4378 36960 4442 36964
rect 4458 37020 4522 37024
rect 4458 36964 4462 37020
rect 4462 36964 4518 37020
rect 4518 36964 4522 37020
rect 4458 36960 4522 36964
rect 4538 37020 4602 37024
rect 4538 36964 4542 37020
rect 4542 36964 4598 37020
rect 4598 36964 4602 37020
rect 4538 36960 4602 36964
rect 4618 37020 4682 37024
rect 4618 36964 4622 37020
rect 4622 36964 4678 37020
rect 4678 36964 4682 37020
rect 4618 36960 4682 36964
rect 7805 37020 7869 37024
rect 7805 36964 7809 37020
rect 7809 36964 7865 37020
rect 7865 36964 7869 37020
rect 7805 36960 7869 36964
rect 7885 37020 7949 37024
rect 7885 36964 7889 37020
rect 7889 36964 7945 37020
rect 7945 36964 7949 37020
rect 7885 36960 7949 36964
rect 7965 37020 8029 37024
rect 7965 36964 7969 37020
rect 7969 36964 8025 37020
rect 8025 36964 8029 37020
rect 7965 36960 8029 36964
rect 8045 37020 8109 37024
rect 8045 36964 8049 37020
rect 8049 36964 8105 37020
rect 8105 36964 8109 37020
rect 8045 36960 8109 36964
rect 11232 37020 11296 37024
rect 11232 36964 11236 37020
rect 11236 36964 11292 37020
rect 11292 36964 11296 37020
rect 11232 36960 11296 36964
rect 11312 37020 11376 37024
rect 11312 36964 11316 37020
rect 11316 36964 11372 37020
rect 11372 36964 11376 37020
rect 11312 36960 11376 36964
rect 11392 37020 11456 37024
rect 11392 36964 11396 37020
rect 11396 36964 11452 37020
rect 11452 36964 11456 37020
rect 11392 36960 11456 36964
rect 11472 37020 11536 37024
rect 11472 36964 11476 37020
rect 11476 36964 11532 37020
rect 11532 36964 11536 37020
rect 11472 36960 11536 36964
rect 14659 37020 14723 37024
rect 14659 36964 14663 37020
rect 14663 36964 14719 37020
rect 14719 36964 14723 37020
rect 14659 36960 14723 36964
rect 14739 37020 14803 37024
rect 14739 36964 14743 37020
rect 14743 36964 14799 37020
rect 14799 36964 14803 37020
rect 14739 36960 14803 36964
rect 14819 37020 14883 37024
rect 14819 36964 14823 37020
rect 14823 36964 14879 37020
rect 14879 36964 14883 37020
rect 14819 36960 14883 36964
rect 14899 37020 14963 37024
rect 14899 36964 14903 37020
rect 14903 36964 14959 37020
rect 14959 36964 14963 37020
rect 14899 36960 14963 36964
rect 2665 36476 2729 36480
rect 2665 36420 2669 36476
rect 2669 36420 2725 36476
rect 2725 36420 2729 36476
rect 2665 36416 2729 36420
rect 2745 36476 2809 36480
rect 2745 36420 2749 36476
rect 2749 36420 2805 36476
rect 2805 36420 2809 36476
rect 2745 36416 2809 36420
rect 2825 36476 2889 36480
rect 2825 36420 2829 36476
rect 2829 36420 2885 36476
rect 2885 36420 2889 36476
rect 2825 36416 2889 36420
rect 2905 36476 2969 36480
rect 2905 36420 2909 36476
rect 2909 36420 2965 36476
rect 2965 36420 2969 36476
rect 2905 36416 2969 36420
rect 6092 36476 6156 36480
rect 6092 36420 6096 36476
rect 6096 36420 6152 36476
rect 6152 36420 6156 36476
rect 6092 36416 6156 36420
rect 6172 36476 6236 36480
rect 6172 36420 6176 36476
rect 6176 36420 6232 36476
rect 6232 36420 6236 36476
rect 6172 36416 6236 36420
rect 6252 36476 6316 36480
rect 6252 36420 6256 36476
rect 6256 36420 6312 36476
rect 6312 36420 6316 36476
rect 6252 36416 6316 36420
rect 6332 36476 6396 36480
rect 6332 36420 6336 36476
rect 6336 36420 6392 36476
rect 6392 36420 6396 36476
rect 6332 36416 6396 36420
rect 9519 36476 9583 36480
rect 9519 36420 9523 36476
rect 9523 36420 9579 36476
rect 9579 36420 9583 36476
rect 9519 36416 9583 36420
rect 9599 36476 9663 36480
rect 9599 36420 9603 36476
rect 9603 36420 9659 36476
rect 9659 36420 9663 36476
rect 9599 36416 9663 36420
rect 9679 36476 9743 36480
rect 9679 36420 9683 36476
rect 9683 36420 9739 36476
rect 9739 36420 9743 36476
rect 9679 36416 9743 36420
rect 9759 36476 9823 36480
rect 9759 36420 9763 36476
rect 9763 36420 9819 36476
rect 9819 36420 9823 36476
rect 9759 36416 9823 36420
rect 12946 36476 13010 36480
rect 12946 36420 12950 36476
rect 12950 36420 13006 36476
rect 13006 36420 13010 36476
rect 12946 36416 13010 36420
rect 13026 36476 13090 36480
rect 13026 36420 13030 36476
rect 13030 36420 13086 36476
rect 13086 36420 13090 36476
rect 13026 36416 13090 36420
rect 13106 36476 13170 36480
rect 13106 36420 13110 36476
rect 13110 36420 13166 36476
rect 13166 36420 13170 36476
rect 13106 36416 13170 36420
rect 13186 36476 13250 36480
rect 13186 36420 13190 36476
rect 13190 36420 13246 36476
rect 13246 36420 13250 36476
rect 13186 36416 13250 36420
rect 4378 35932 4442 35936
rect 4378 35876 4382 35932
rect 4382 35876 4438 35932
rect 4438 35876 4442 35932
rect 4378 35872 4442 35876
rect 4458 35932 4522 35936
rect 4458 35876 4462 35932
rect 4462 35876 4518 35932
rect 4518 35876 4522 35932
rect 4458 35872 4522 35876
rect 4538 35932 4602 35936
rect 4538 35876 4542 35932
rect 4542 35876 4598 35932
rect 4598 35876 4602 35932
rect 4538 35872 4602 35876
rect 4618 35932 4682 35936
rect 4618 35876 4622 35932
rect 4622 35876 4678 35932
rect 4678 35876 4682 35932
rect 4618 35872 4682 35876
rect 7805 35932 7869 35936
rect 7805 35876 7809 35932
rect 7809 35876 7865 35932
rect 7865 35876 7869 35932
rect 7805 35872 7869 35876
rect 7885 35932 7949 35936
rect 7885 35876 7889 35932
rect 7889 35876 7945 35932
rect 7945 35876 7949 35932
rect 7885 35872 7949 35876
rect 7965 35932 8029 35936
rect 7965 35876 7969 35932
rect 7969 35876 8025 35932
rect 8025 35876 8029 35932
rect 7965 35872 8029 35876
rect 8045 35932 8109 35936
rect 8045 35876 8049 35932
rect 8049 35876 8105 35932
rect 8105 35876 8109 35932
rect 8045 35872 8109 35876
rect 11232 35932 11296 35936
rect 11232 35876 11236 35932
rect 11236 35876 11292 35932
rect 11292 35876 11296 35932
rect 11232 35872 11296 35876
rect 11312 35932 11376 35936
rect 11312 35876 11316 35932
rect 11316 35876 11372 35932
rect 11372 35876 11376 35932
rect 11312 35872 11376 35876
rect 11392 35932 11456 35936
rect 11392 35876 11396 35932
rect 11396 35876 11452 35932
rect 11452 35876 11456 35932
rect 11392 35872 11456 35876
rect 11472 35932 11536 35936
rect 11472 35876 11476 35932
rect 11476 35876 11532 35932
rect 11532 35876 11536 35932
rect 11472 35872 11536 35876
rect 14659 35932 14723 35936
rect 14659 35876 14663 35932
rect 14663 35876 14719 35932
rect 14719 35876 14723 35932
rect 14659 35872 14723 35876
rect 14739 35932 14803 35936
rect 14739 35876 14743 35932
rect 14743 35876 14799 35932
rect 14799 35876 14803 35932
rect 14739 35872 14803 35876
rect 14819 35932 14883 35936
rect 14819 35876 14823 35932
rect 14823 35876 14879 35932
rect 14879 35876 14883 35932
rect 14819 35872 14883 35876
rect 14899 35932 14963 35936
rect 14899 35876 14903 35932
rect 14903 35876 14959 35932
rect 14959 35876 14963 35932
rect 14899 35872 14963 35876
rect 2665 35388 2729 35392
rect 2665 35332 2669 35388
rect 2669 35332 2725 35388
rect 2725 35332 2729 35388
rect 2665 35328 2729 35332
rect 2745 35388 2809 35392
rect 2745 35332 2749 35388
rect 2749 35332 2805 35388
rect 2805 35332 2809 35388
rect 2745 35328 2809 35332
rect 2825 35388 2889 35392
rect 2825 35332 2829 35388
rect 2829 35332 2885 35388
rect 2885 35332 2889 35388
rect 2825 35328 2889 35332
rect 2905 35388 2969 35392
rect 2905 35332 2909 35388
rect 2909 35332 2965 35388
rect 2965 35332 2969 35388
rect 2905 35328 2969 35332
rect 6092 35388 6156 35392
rect 6092 35332 6096 35388
rect 6096 35332 6152 35388
rect 6152 35332 6156 35388
rect 6092 35328 6156 35332
rect 6172 35388 6236 35392
rect 6172 35332 6176 35388
rect 6176 35332 6232 35388
rect 6232 35332 6236 35388
rect 6172 35328 6236 35332
rect 6252 35388 6316 35392
rect 6252 35332 6256 35388
rect 6256 35332 6312 35388
rect 6312 35332 6316 35388
rect 6252 35328 6316 35332
rect 6332 35388 6396 35392
rect 6332 35332 6336 35388
rect 6336 35332 6392 35388
rect 6392 35332 6396 35388
rect 6332 35328 6396 35332
rect 9519 35388 9583 35392
rect 9519 35332 9523 35388
rect 9523 35332 9579 35388
rect 9579 35332 9583 35388
rect 9519 35328 9583 35332
rect 9599 35388 9663 35392
rect 9599 35332 9603 35388
rect 9603 35332 9659 35388
rect 9659 35332 9663 35388
rect 9599 35328 9663 35332
rect 9679 35388 9743 35392
rect 9679 35332 9683 35388
rect 9683 35332 9739 35388
rect 9739 35332 9743 35388
rect 9679 35328 9743 35332
rect 9759 35388 9823 35392
rect 9759 35332 9763 35388
rect 9763 35332 9819 35388
rect 9819 35332 9823 35388
rect 9759 35328 9823 35332
rect 12946 35388 13010 35392
rect 12946 35332 12950 35388
rect 12950 35332 13006 35388
rect 13006 35332 13010 35388
rect 12946 35328 13010 35332
rect 13026 35388 13090 35392
rect 13026 35332 13030 35388
rect 13030 35332 13086 35388
rect 13086 35332 13090 35388
rect 13026 35328 13090 35332
rect 13106 35388 13170 35392
rect 13106 35332 13110 35388
rect 13110 35332 13166 35388
rect 13166 35332 13170 35388
rect 13106 35328 13170 35332
rect 13186 35388 13250 35392
rect 13186 35332 13190 35388
rect 13190 35332 13246 35388
rect 13246 35332 13250 35388
rect 13186 35328 13250 35332
rect 4378 34844 4442 34848
rect 4378 34788 4382 34844
rect 4382 34788 4438 34844
rect 4438 34788 4442 34844
rect 4378 34784 4442 34788
rect 4458 34844 4522 34848
rect 4458 34788 4462 34844
rect 4462 34788 4518 34844
rect 4518 34788 4522 34844
rect 4458 34784 4522 34788
rect 4538 34844 4602 34848
rect 4538 34788 4542 34844
rect 4542 34788 4598 34844
rect 4598 34788 4602 34844
rect 4538 34784 4602 34788
rect 4618 34844 4682 34848
rect 4618 34788 4622 34844
rect 4622 34788 4678 34844
rect 4678 34788 4682 34844
rect 4618 34784 4682 34788
rect 7805 34844 7869 34848
rect 7805 34788 7809 34844
rect 7809 34788 7865 34844
rect 7865 34788 7869 34844
rect 7805 34784 7869 34788
rect 7885 34844 7949 34848
rect 7885 34788 7889 34844
rect 7889 34788 7945 34844
rect 7945 34788 7949 34844
rect 7885 34784 7949 34788
rect 7965 34844 8029 34848
rect 7965 34788 7969 34844
rect 7969 34788 8025 34844
rect 8025 34788 8029 34844
rect 7965 34784 8029 34788
rect 8045 34844 8109 34848
rect 8045 34788 8049 34844
rect 8049 34788 8105 34844
rect 8105 34788 8109 34844
rect 8045 34784 8109 34788
rect 11232 34844 11296 34848
rect 11232 34788 11236 34844
rect 11236 34788 11292 34844
rect 11292 34788 11296 34844
rect 11232 34784 11296 34788
rect 11312 34844 11376 34848
rect 11312 34788 11316 34844
rect 11316 34788 11372 34844
rect 11372 34788 11376 34844
rect 11312 34784 11376 34788
rect 11392 34844 11456 34848
rect 11392 34788 11396 34844
rect 11396 34788 11452 34844
rect 11452 34788 11456 34844
rect 11392 34784 11456 34788
rect 11472 34844 11536 34848
rect 11472 34788 11476 34844
rect 11476 34788 11532 34844
rect 11532 34788 11536 34844
rect 11472 34784 11536 34788
rect 14659 34844 14723 34848
rect 14659 34788 14663 34844
rect 14663 34788 14719 34844
rect 14719 34788 14723 34844
rect 14659 34784 14723 34788
rect 14739 34844 14803 34848
rect 14739 34788 14743 34844
rect 14743 34788 14799 34844
rect 14799 34788 14803 34844
rect 14739 34784 14803 34788
rect 14819 34844 14883 34848
rect 14819 34788 14823 34844
rect 14823 34788 14879 34844
rect 14879 34788 14883 34844
rect 14819 34784 14883 34788
rect 14899 34844 14963 34848
rect 14899 34788 14903 34844
rect 14903 34788 14959 34844
rect 14959 34788 14963 34844
rect 14899 34784 14963 34788
rect 2665 34300 2729 34304
rect 2665 34244 2669 34300
rect 2669 34244 2725 34300
rect 2725 34244 2729 34300
rect 2665 34240 2729 34244
rect 2745 34300 2809 34304
rect 2745 34244 2749 34300
rect 2749 34244 2805 34300
rect 2805 34244 2809 34300
rect 2745 34240 2809 34244
rect 2825 34300 2889 34304
rect 2825 34244 2829 34300
rect 2829 34244 2885 34300
rect 2885 34244 2889 34300
rect 2825 34240 2889 34244
rect 2905 34300 2969 34304
rect 2905 34244 2909 34300
rect 2909 34244 2965 34300
rect 2965 34244 2969 34300
rect 2905 34240 2969 34244
rect 6092 34300 6156 34304
rect 6092 34244 6096 34300
rect 6096 34244 6152 34300
rect 6152 34244 6156 34300
rect 6092 34240 6156 34244
rect 6172 34300 6236 34304
rect 6172 34244 6176 34300
rect 6176 34244 6232 34300
rect 6232 34244 6236 34300
rect 6172 34240 6236 34244
rect 6252 34300 6316 34304
rect 6252 34244 6256 34300
rect 6256 34244 6312 34300
rect 6312 34244 6316 34300
rect 6252 34240 6316 34244
rect 6332 34300 6396 34304
rect 6332 34244 6336 34300
rect 6336 34244 6392 34300
rect 6392 34244 6396 34300
rect 6332 34240 6396 34244
rect 9519 34300 9583 34304
rect 9519 34244 9523 34300
rect 9523 34244 9579 34300
rect 9579 34244 9583 34300
rect 9519 34240 9583 34244
rect 9599 34300 9663 34304
rect 9599 34244 9603 34300
rect 9603 34244 9659 34300
rect 9659 34244 9663 34300
rect 9599 34240 9663 34244
rect 9679 34300 9743 34304
rect 9679 34244 9683 34300
rect 9683 34244 9739 34300
rect 9739 34244 9743 34300
rect 9679 34240 9743 34244
rect 9759 34300 9823 34304
rect 9759 34244 9763 34300
rect 9763 34244 9819 34300
rect 9819 34244 9823 34300
rect 9759 34240 9823 34244
rect 12946 34300 13010 34304
rect 12946 34244 12950 34300
rect 12950 34244 13006 34300
rect 13006 34244 13010 34300
rect 12946 34240 13010 34244
rect 13026 34300 13090 34304
rect 13026 34244 13030 34300
rect 13030 34244 13086 34300
rect 13086 34244 13090 34300
rect 13026 34240 13090 34244
rect 13106 34300 13170 34304
rect 13106 34244 13110 34300
rect 13110 34244 13166 34300
rect 13166 34244 13170 34300
rect 13106 34240 13170 34244
rect 13186 34300 13250 34304
rect 13186 34244 13190 34300
rect 13190 34244 13246 34300
rect 13246 34244 13250 34300
rect 13186 34240 13250 34244
rect 4378 33756 4442 33760
rect 4378 33700 4382 33756
rect 4382 33700 4438 33756
rect 4438 33700 4442 33756
rect 4378 33696 4442 33700
rect 4458 33756 4522 33760
rect 4458 33700 4462 33756
rect 4462 33700 4518 33756
rect 4518 33700 4522 33756
rect 4458 33696 4522 33700
rect 4538 33756 4602 33760
rect 4538 33700 4542 33756
rect 4542 33700 4598 33756
rect 4598 33700 4602 33756
rect 4538 33696 4602 33700
rect 4618 33756 4682 33760
rect 4618 33700 4622 33756
rect 4622 33700 4678 33756
rect 4678 33700 4682 33756
rect 4618 33696 4682 33700
rect 7805 33756 7869 33760
rect 7805 33700 7809 33756
rect 7809 33700 7865 33756
rect 7865 33700 7869 33756
rect 7805 33696 7869 33700
rect 7885 33756 7949 33760
rect 7885 33700 7889 33756
rect 7889 33700 7945 33756
rect 7945 33700 7949 33756
rect 7885 33696 7949 33700
rect 7965 33756 8029 33760
rect 7965 33700 7969 33756
rect 7969 33700 8025 33756
rect 8025 33700 8029 33756
rect 7965 33696 8029 33700
rect 8045 33756 8109 33760
rect 8045 33700 8049 33756
rect 8049 33700 8105 33756
rect 8105 33700 8109 33756
rect 8045 33696 8109 33700
rect 11232 33756 11296 33760
rect 11232 33700 11236 33756
rect 11236 33700 11292 33756
rect 11292 33700 11296 33756
rect 11232 33696 11296 33700
rect 11312 33756 11376 33760
rect 11312 33700 11316 33756
rect 11316 33700 11372 33756
rect 11372 33700 11376 33756
rect 11312 33696 11376 33700
rect 11392 33756 11456 33760
rect 11392 33700 11396 33756
rect 11396 33700 11452 33756
rect 11452 33700 11456 33756
rect 11392 33696 11456 33700
rect 11472 33756 11536 33760
rect 11472 33700 11476 33756
rect 11476 33700 11532 33756
rect 11532 33700 11536 33756
rect 11472 33696 11536 33700
rect 14659 33756 14723 33760
rect 14659 33700 14663 33756
rect 14663 33700 14719 33756
rect 14719 33700 14723 33756
rect 14659 33696 14723 33700
rect 14739 33756 14803 33760
rect 14739 33700 14743 33756
rect 14743 33700 14799 33756
rect 14799 33700 14803 33756
rect 14739 33696 14803 33700
rect 14819 33756 14883 33760
rect 14819 33700 14823 33756
rect 14823 33700 14879 33756
rect 14879 33700 14883 33756
rect 14819 33696 14883 33700
rect 14899 33756 14963 33760
rect 14899 33700 14903 33756
rect 14903 33700 14959 33756
rect 14959 33700 14963 33756
rect 14899 33696 14963 33700
rect 2665 33212 2729 33216
rect 2665 33156 2669 33212
rect 2669 33156 2725 33212
rect 2725 33156 2729 33212
rect 2665 33152 2729 33156
rect 2745 33212 2809 33216
rect 2745 33156 2749 33212
rect 2749 33156 2805 33212
rect 2805 33156 2809 33212
rect 2745 33152 2809 33156
rect 2825 33212 2889 33216
rect 2825 33156 2829 33212
rect 2829 33156 2885 33212
rect 2885 33156 2889 33212
rect 2825 33152 2889 33156
rect 2905 33212 2969 33216
rect 2905 33156 2909 33212
rect 2909 33156 2965 33212
rect 2965 33156 2969 33212
rect 2905 33152 2969 33156
rect 6092 33212 6156 33216
rect 6092 33156 6096 33212
rect 6096 33156 6152 33212
rect 6152 33156 6156 33212
rect 6092 33152 6156 33156
rect 6172 33212 6236 33216
rect 6172 33156 6176 33212
rect 6176 33156 6232 33212
rect 6232 33156 6236 33212
rect 6172 33152 6236 33156
rect 6252 33212 6316 33216
rect 6252 33156 6256 33212
rect 6256 33156 6312 33212
rect 6312 33156 6316 33212
rect 6252 33152 6316 33156
rect 6332 33212 6396 33216
rect 6332 33156 6336 33212
rect 6336 33156 6392 33212
rect 6392 33156 6396 33212
rect 6332 33152 6396 33156
rect 9519 33212 9583 33216
rect 9519 33156 9523 33212
rect 9523 33156 9579 33212
rect 9579 33156 9583 33212
rect 9519 33152 9583 33156
rect 9599 33212 9663 33216
rect 9599 33156 9603 33212
rect 9603 33156 9659 33212
rect 9659 33156 9663 33212
rect 9599 33152 9663 33156
rect 9679 33212 9743 33216
rect 9679 33156 9683 33212
rect 9683 33156 9739 33212
rect 9739 33156 9743 33212
rect 9679 33152 9743 33156
rect 9759 33212 9823 33216
rect 9759 33156 9763 33212
rect 9763 33156 9819 33212
rect 9819 33156 9823 33212
rect 9759 33152 9823 33156
rect 12946 33212 13010 33216
rect 12946 33156 12950 33212
rect 12950 33156 13006 33212
rect 13006 33156 13010 33212
rect 12946 33152 13010 33156
rect 13026 33212 13090 33216
rect 13026 33156 13030 33212
rect 13030 33156 13086 33212
rect 13086 33156 13090 33212
rect 13026 33152 13090 33156
rect 13106 33212 13170 33216
rect 13106 33156 13110 33212
rect 13110 33156 13166 33212
rect 13166 33156 13170 33212
rect 13106 33152 13170 33156
rect 13186 33212 13250 33216
rect 13186 33156 13190 33212
rect 13190 33156 13246 33212
rect 13246 33156 13250 33212
rect 13186 33152 13250 33156
rect 4378 32668 4442 32672
rect 4378 32612 4382 32668
rect 4382 32612 4438 32668
rect 4438 32612 4442 32668
rect 4378 32608 4442 32612
rect 4458 32668 4522 32672
rect 4458 32612 4462 32668
rect 4462 32612 4518 32668
rect 4518 32612 4522 32668
rect 4458 32608 4522 32612
rect 4538 32668 4602 32672
rect 4538 32612 4542 32668
rect 4542 32612 4598 32668
rect 4598 32612 4602 32668
rect 4538 32608 4602 32612
rect 4618 32668 4682 32672
rect 4618 32612 4622 32668
rect 4622 32612 4678 32668
rect 4678 32612 4682 32668
rect 4618 32608 4682 32612
rect 7805 32668 7869 32672
rect 7805 32612 7809 32668
rect 7809 32612 7865 32668
rect 7865 32612 7869 32668
rect 7805 32608 7869 32612
rect 7885 32668 7949 32672
rect 7885 32612 7889 32668
rect 7889 32612 7945 32668
rect 7945 32612 7949 32668
rect 7885 32608 7949 32612
rect 7965 32668 8029 32672
rect 7965 32612 7969 32668
rect 7969 32612 8025 32668
rect 8025 32612 8029 32668
rect 7965 32608 8029 32612
rect 8045 32668 8109 32672
rect 8045 32612 8049 32668
rect 8049 32612 8105 32668
rect 8105 32612 8109 32668
rect 8045 32608 8109 32612
rect 11232 32668 11296 32672
rect 11232 32612 11236 32668
rect 11236 32612 11292 32668
rect 11292 32612 11296 32668
rect 11232 32608 11296 32612
rect 11312 32668 11376 32672
rect 11312 32612 11316 32668
rect 11316 32612 11372 32668
rect 11372 32612 11376 32668
rect 11312 32608 11376 32612
rect 11392 32668 11456 32672
rect 11392 32612 11396 32668
rect 11396 32612 11452 32668
rect 11452 32612 11456 32668
rect 11392 32608 11456 32612
rect 11472 32668 11536 32672
rect 11472 32612 11476 32668
rect 11476 32612 11532 32668
rect 11532 32612 11536 32668
rect 11472 32608 11536 32612
rect 14659 32668 14723 32672
rect 14659 32612 14663 32668
rect 14663 32612 14719 32668
rect 14719 32612 14723 32668
rect 14659 32608 14723 32612
rect 14739 32668 14803 32672
rect 14739 32612 14743 32668
rect 14743 32612 14799 32668
rect 14799 32612 14803 32668
rect 14739 32608 14803 32612
rect 14819 32668 14883 32672
rect 14819 32612 14823 32668
rect 14823 32612 14879 32668
rect 14879 32612 14883 32668
rect 14819 32608 14883 32612
rect 14899 32668 14963 32672
rect 14899 32612 14903 32668
rect 14903 32612 14959 32668
rect 14959 32612 14963 32668
rect 14899 32608 14963 32612
rect 12020 32404 12084 32468
rect 11836 32328 11900 32332
rect 11836 32272 11850 32328
rect 11850 32272 11900 32328
rect 11836 32268 11900 32272
rect 2665 32124 2729 32128
rect 2665 32068 2669 32124
rect 2669 32068 2725 32124
rect 2725 32068 2729 32124
rect 2665 32064 2729 32068
rect 2745 32124 2809 32128
rect 2745 32068 2749 32124
rect 2749 32068 2805 32124
rect 2805 32068 2809 32124
rect 2745 32064 2809 32068
rect 2825 32124 2889 32128
rect 2825 32068 2829 32124
rect 2829 32068 2885 32124
rect 2885 32068 2889 32124
rect 2825 32064 2889 32068
rect 2905 32124 2969 32128
rect 2905 32068 2909 32124
rect 2909 32068 2965 32124
rect 2965 32068 2969 32124
rect 2905 32064 2969 32068
rect 6092 32124 6156 32128
rect 6092 32068 6096 32124
rect 6096 32068 6152 32124
rect 6152 32068 6156 32124
rect 6092 32064 6156 32068
rect 6172 32124 6236 32128
rect 6172 32068 6176 32124
rect 6176 32068 6232 32124
rect 6232 32068 6236 32124
rect 6172 32064 6236 32068
rect 6252 32124 6316 32128
rect 6252 32068 6256 32124
rect 6256 32068 6312 32124
rect 6312 32068 6316 32124
rect 6252 32064 6316 32068
rect 6332 32124 6396 32128
rect 6332 32068 6336 32124
rect 6336 32068 6392 32124
rect 6392 32068 6396 32124
rect 6332 32064 6396 32068
rect 9519 32124 9583 32128
rect 9519 32068 9523 32124
rect 9523 32068 9579 32124
rect 9579 32068 9583 32124
rect 9519 32064 9583 32068
rect 9599 32124 9663 32128
rect 9599 32068 9603 32124
rect 9603 32068 9659 32124
rect 9659 32068 9663 32124
rect 9599 32064 9663 32068
rect 9679 32124 9743 32128
rect 9679 32068 9683 32124
rect 9683 32068 9739 32124
rect 9739 32068 9743 32124
rect 9679 32064 9743 32068
rect 9759 32124 9823 32128
rect 9759 32068 9763 32124
rect 9763 32068 9819 32124
rect 9819 32068 9823 32124
rect 9759 32064 9823 32068
rect 12946 32124 13010 32128
rect 12946 32068 12950 32124
rect 12950 32068 13006 32124
rect 13006 32068 13010 32124
rect 12946 32064 13010 32068
rect 13026 32124 13090 32128
rect 13026 32068 13030 32124
rect 13030 32068 13086 32124
rect 13086 32068 13090 32124
rect 13026 32064 13090 32068
rect 13106 32124 13170 32128
rect 13106 32068 13110 32124
rect 13110 32068 13166 32124
rect 13166 32068 13170 32124
rect 13106 32064 13170 32068
rect 13186 32124 13250 32128
rect 13186 32068 13190 32124
rect 13190 32068 13246 32124
rect 13246 32068 13250 32124
rect 13186 32064 13250 32068
rect 12572 31784 12636 31788
rect 12572 31728 12622 31784
rect 12622 31728 12636 31784
rect 12572 31724 12636 31728
rect 4378 31580 4442 31584
rect 4378 31524 4382 31580
rect 4382 31524 4438 31580
rect 4438 31524 4442 31580
rect 4378 31520 4442 31524
rect 4458 31580 4522 31584
rect 4458 31524 4462 31580
rect 4462 31524 4518 31580
rect 4518 31524 4522 31580
rect 4458 31520 4522 31524
rect 4538 31580 4602 31584
rect 4538 31524 4542 31580
rect 4542 31524 4598 31580
rect 4598 31524 4602 31580
rect 4538 31520 4602 31524
rect 4618 31580 4682 31584
rect 4618 31524 4622 31580
rect 4622 31524 4678 31580
rect 4678 31524 4682 31580
rect 4618 31520 4682 31524
rect 7805 31580 7869 31584
rect 7805 31524 7809 31580
rect 7809 31524 7865 31580
rect 7865 31524 7869 31580
rect 7805 31520 7869 31524
rect 7885 31580 7949 31584
rect 7885 31524 7889 31580
rect 7889 31524 7945 31580
rect 7945 31524 7949 31580
rect 7885 31520 7949 31524
rect 7965 31580 8029 31584
rect 7965 31524 7969 31580
rect 7969 31524 8025 31580
rect 8025 31524 8029 31580
rect 7965 31520 8029 31524
rect 8045 31580 8109 31584
rect 8045 31524 8049 31580
rect 8049 31524 8105 31580
rect 8105 31524 8109 31580
rect 8045 31520 8109 31524
rect 11232 31580 11296 31584
rect 11232 31524 11236 31580
rect 11236 31524 11292 31580
rect 11292 31524 11296 31580
rect 11232 31520 11296 31524
rect 11312 31580 11376 31584
rect 11312 31524 11316 31580
rect 11316 31524 11372 31580
rect 11372 31524 11376 31580
rect 11312 31520 11376 31524
rect 11392 31580 11456 31584
rect 11392 31524 11396 31580
rect 11396 31524 11452 31580
rect 11452 31524 11456 31580
rect 11392 31520 11456 31524
rect 11472 31580 11536 31584
rect 11472 31524 11476 31580
rect 11476 31524 11532 31580
rect 11532 31524 11536 31580
rect 11472 31520 11536 31524
rect 14659 31580 14723 31584
rect 14659 31524 14663 31580
rect 14663 31524 14719 31580
rect 14719 31524 14723 31580
rect 14659 31520 14723 31524
rect 14739 31580 14803 31584
rect 14739 31524 14743 31580
rect 14743 31524 14799 31580
rect 14799 31524 14803 31580
rect 14739 31520 14803 31524
rect 14819 31580 14883 31584
rect 14819 31524 14823 31580
rect 14823 31524 14879 31580
rect 14879 31524 14883 31580
rect 14819 31520 14883 31524
rect 14899 31580 14963 31584
rect 14899 31524 14903 31580
rect 14903 31524 14959 31580
rect 14959 31524 14963 31580
rect 14899 31520 14963 31524
rect 2665 31036 2729 31040
rect 2665 30980 2669 31036
rect 2669 30980 2725 31036
rect 2725 30980 2729 31036
rect 2665 30976 2729 30980
rect 2745 31036 2809 31040
rect 2745 30980 2749 31036
rect 2749 30980 2805 31036
rect 2805 30980 2809 31036
rect 2745 30976 2809 30980
rect 2825 31036 2889 31040
rect 2825 30980 2829 31036
rect 2829 30980 2885 31036
rect 2885 30980 2889 31036
rect 2825 30976 2889 30980
rect 2905 31036 2969 31040
rect 2905 30980 2909 31036
rect 2909 30980 2965 31036
rect 2965 30980 2969 31036
rect 2905 30976 2969 30980
rect 6092 31036 6156 31040
rect 6092 30980 6096 31036
rect 6096 30980 6152 31036
rect 6152 30980 6156 31036
rect 6092 30976 6156 30980
rect 6172 31036 6236 31040
rect 6172 30980 6176 31036
rect 6176 30980 6232 31036
rect 6232 30980 6236 31036
rect 6172 30976 6236 30980
rect 6252 31036 6316 31040
rect 6252 30980 6256 31036
rect 6256 30980 6312 31036
rect 6312 30980 6316 31036
rect 6252 30976 6316 30980
rect 6332 31036 6396 31040
rect 6332 30980 6336 31036
rect 6336 30980 6392 31036
rect 6392 30980 6396 31036
rect 6332 30976 6396 30980
rect 9519 31036 9583 31040
rect 9519 30980 9523 31036
rect 9523 30980 9579 31036
rect 9579 30980 9583 31036
rect 9519 30976 9583 30980
rect 9599 31036 9663 31040
rect 9599 30980 9603 31036
rect 9603 30980 9659 31036
rect 9659 30980 9663 31036
rect 9599 30976 9663 30980
rect 9679 31036 9743 31040
rect 9679 30980 9683 31036
rect 9683 30980 9739 31036
rect 9739 30980 9743 31036
rect 9679 30976 9743 30980
rect 9759 31036 9823 31040
rect 9759 30980 9763 31036
rect 9763 30980 9819 31036
rect 9819 30980 9823 31036
rect 9759 30976 9823 30980
rect 12946 31036 13010 31040
rect 12946 30980 12950 31036
rect 12950 30980 13006 31036
rect 13006 30980 13010 31036
rect 12946 30976 13010 30980
rect 13026 31036 13090 31040
rect 13026 30980 13030 31036
rect 13030 30980 13086 31036
rect 13086 30980 13090 31036
rect 13026 30976 13090 30980
rect 13106 31036 13170 31040
rect 13106 30980 13110 31036
rect 13110 30980 13166 31036
rect 13166 30980 13170 31036
rect 13106 30976 13170 30980
rect 13186 31036 13250 31040
rect 13186 30980 13190 31036
rect 13190 30980 13246 31036
rect 13246 30980 13250 31036
rect 13186 30976 13250 30980
rect 4378 30492 4442 30496
rect 4378 30436 4382 30492
rect 4382 30436 4438 30492
rect 4438 30436 4442 30492
rect 4378 30432 4442 30436
rect 4458 30492 4522 30496
rect 4458 30436 4462 30492
rect 4462 30436 4518 30492
rect 4518 30436 4522 30492
rect 4458 30432 4522 30436
rect 4538 30492 4602 30496
rect 4538 30436 4542 30492
rect 4542 30436 4598 30492
rect 4598 30436 4602 30492
rect 4538 30432 4602 30436
rect 4618 30492 4682 30496
rect 4618 30436 4622 30492
rect 4622 30436 4678 30492
rect 4678 30436 4682 30492
rect 4618 30432 4682 30436
rect 7805 30492 7869 30496
rect 7805 30436 7809 30492
rect 7809 30436 7865 30492
rect 7865 30436 7869 30492
rect 7805 30432 7869 30436
rect 7885 30492 7949 30496
rect 7885 30436 7889 30492
rect 7889 30436 7945 30492
rect 7945 30436 7949 30492
rect 7885 30432 7949 30436
rect 7965 30492 8029 30496
rect 7965 30436 7969 30492
rect 7969 30436 8025 30492
rect 8025 30436 8029 30492
rect 7965 30432 8029 30436
rect 8045 30492 8109 30496
rect 8045 30436 8049 30492
rect 8049 30436 8105 30492
rect 8105 30436 8109 30492
rect 8045 30432 8109 30436
rect 11232 30492 11296 30496
rect 11232 30436 11236 30492
rect 11236 30436 11292 30492
rect 11292 30436 11296 30492
rect 11232 30432 11296 30436
rect 11312 30492 11376 30496
rect 11312 30436 11316 30492
rect 11316 30436 11372 30492
rect 11372 30436 11376 30492
rect 11312 30432 11376 30436
rect 11392 30492 11456 30496
rect 11392 30436 11396 30492
rect 11396 30436 11452 30492
rect 11452 30436 11456 30492
rect 11392 30432 11456 30436
rect 11472 30492 11536 30496
rect 11472 30436 11476 30492
rect 11476 30436 11532 30492
rect 11532 30436 11536 30492
rect 11472 30432 11536 30436
rect 14659 30492 14723 30496
rect 14659 30436 14663 30492
rect 14663 30436 14719 30492
rect 14719 30436 14723 30492
rect 14659 30432 14723 30436
rect 14739 30492 14803 30496
rect 14739 30436 14743 30492
rect 14743 30436 14799 30492
rect 14799 30436 14803 30492
rect 14739 30432 14803 30436
rect 14819 30492 14883 30496
rect 14819 30436 14823 30492
rect 14823 30436 14879 30492
rect 14879 30436 14883 30492
rect 14819 30432 14883 30436
rect 14899 30492 14963 30496
rect 14899 30436 14903 30492
rect 14903 30436 14959 30492
rect 14959 30436 14963 30492
rect 14899 30432 14963 30436
rect 2665 29948 2729 29952
rect 2665 29892 2669 29948
rect 2669 29892 2725 29948
rect 2725 29892 2729 29948
rect 2665 29888 2729 29892
rect 2745 29948 2809 29952
rect 2745 29892 2749 29948
rect 2749 29892 2805 29948
rect 2805 29892 2809 29948
rect 2745 29888 2809 29892
rect 2825 29948 2889 29952
rect 2825 29892 2829 29948
rect 2829 29892 2885 29948
rect 2885 29892 2889 29948
rect 2825 29888 2889 29892
rect 2905 29948 2969 29952
rect 2905 29892 2909 29948
rect 2909 29892 2965 29948
rect 2965 29892 2969 29948
rect 2905 29888 2969 29892
rect 6092 29948 6156 29952
rect 6092 29892 6096 29948
rect 6096 29892 6152 29948
rect 6152 29892 6156 29948
rect 6092 29888 6156 29892
rect 6172 29948 6236 29952
rect 6172 29892 6176 29948
rect 6176 29892 6232 29948
rect 6232 29892 6236 29948
rect 6172 29888 6236 29892
rect 6252 29948 6316 29952
rect 6252 29892 6256 29948
rect 6256 29892 6312 29948
rect 6312 29892 6316 29948
rect 6252 29888 6316 29892
rect 6332 29948 6396 29952
rect 6332 29892 6336 29948
rect 6336 29892 6392 29948
rect 6392 29892 6396 29948
rect 6332 29888 6396 29892
rect 9519 29948 9583 29952
rect 9519 29892 9523 29948
rect 9523 29892 9579 29948
rect 9579 29892 9583 29948
rect 9519 29888 9583 29892
rect 9599 29948 9663 29952
rect 9599 29892 9603 29948
rect 9603 29892 9659 29948
rect 9659 29892 9663 29948
rect 9599 29888 9663 29892
rect 9679 29948 9743 29952
rect 9679 29892 9683 29948
rect 9683 29892 9739 29948
rect 9739 29892 9743 29948
rect 9679 29888 9743 29892
rect 9759 29948 9823 29952
rect 9759 29892 9763 29948
rect 9763 29892 9819 29948
rect 9819 29892 9823 29948
rect 9759 29888 9823 29892
rect 12946 29948 13010 29952
rect 12946 29892 12950 29948
rect 12950 29892 13006 29948
rect 13006 29892 13010 29948
rect 12946 29888 13010 29892
rect 13026 29948 13090 29952
rect 13026 29892 13030 29948
rect 13030 29892 13086 29948
rect 13086 29892 13090 29948
rect 13026 29888 13090 29892
rect 13106 29948 13170 29952
rect 13106 29892 13110 29948
rect 13110 29892 13166 29948
rect 13166 29892 13170 29948
rect 13106 29888 13170 29892
rect 13186 29948 13250 29952
rect 13186 29892 13190 29948
rect 13190 29892 13246 29948
rect 13246 29892 13250 29948
rect 13186 29888 13250 29892
rect 4378 29404 4442 29408
rect 4378 29348 4382 29404
rect 4382 29348 4438 29404
rect 4438 29348 4442 29404
rect 4378 29344 4442 29348
rect 4458 29404 4522 29408
rect 4458 29348 4462 29404
rect 4462 29348 4518 29404
rect 4518 29348 4522 29404
rect 4458 29344 4522 29348
rect 4538 29404 4602 29408
rect 4538 29348 4542 29404
rect 4542 29348 4598 29404
rect 4598 29348 4602 29404
rect 4538 29344 4602 29348
rect 4618 29404 4682 29408
rect 4618 29348 4622 29404
rect 4622 29348 4678 29404
rect 4678 29348 4682 29404
rect 4618 29344 4682 29348
rect 7805 29404 7869 29408
rect 7805 29348 7809 29404
rect 7809 29348 7865 29404
rect 7865 29348 7869 29404
rect 7805 29344 7869 29348
rect 7885 29404 7949 29408
rect 7885 29348 7889 29404
rect 7889 29348 7945 29404
rect 7945 29348 7949 29404
rect 7885 29344 7949 29348
rect 7965 29404 8029 29408
rect 7965 29348 7969 29404
rect 7969 29348 8025 29404
rect 8025 29348 8029 29404
rect 7965 29344 8029 29348
rect 8045 29404 8109 29408
rect 8045 29348 8049 29404
rect 8049 29348 8105 29404
rect 8105 29348 8109 29404
rect 8045 29344 8109 29348
rect 11232 29404 11296 29408
rect 11232 29348 11236 29404
rect 11236 29348 11292 29404
rect 11292 29348 11296 29404
rect 11232 29344 11296 29348
rect 11312 29404 11376 29408
rect 11312 29348 11316 29404
rect 11316 29348 11372 29404
rect 11372 29348 11376 29404
rect 11312 29344 11376 29348
rect 11392 29404 11456 29408
rect 11392 29348 11396 29404
rect 11396 29348 11452 29404
rect 11452 29348 11456 29404
rect 11392 29344 11456 29348
rect 11472 29404 11536 29408
rect 11472 29348 11476 29404
rect 11476 29348 11532 29404
rect 11532 29348 11536 29404
rect 11472 29344 11536 29348
rect 14659 29404 14723 29408
rect 14659 29348 14663 29404
rect 14663 29348 14719 29404
rect 14719 29348 14723 29404
rect 14659 29344 14723 29348
rect 14739 29404 14803 29408
rect 14739 29348 14743 29404
rect 14743 29348 14799 29404
rect 14799 29348 14803 29404
rect 14739 29344 14803 29348
rect 14819 29404 14883 29408
rect 14819 29348 14823 29404
rect 14823 29348 14879 29404
rect 14879 29348 14883 29404
rect 14819 29344 14883 29348
rect 14899 29404 14963 29408
rect 14899 29348 14903 29404
rect 14903 29348 14959 29404
rect 14959 29348 14963 29404
rect 14899 29344 14963 29348
rect 9076 29004 9140 29068
rect 9260 29064 9324 29068
rect 9260 29008 9274 29064
rect 9274 29008 9324 29064
rect 9260 29004 9324 29008
rect 12020 28928 12084 28932
rect 12020 28872 12034 28928
rect 12034 28872 12084 28928
rect 12020 28868 12084 28872
rect 2665 28860 2729 28864
rect 2665 28804 2669 28860
rect 2669 28804 2725 28860
rect 2725 28804 2729 28860
rect 2665 28800 2729 28804
rect 2745 28860 2809 28864
rect 2745 28804 2749 28860
rect 2749 28804 2805 28860
rect 2805 28804 2809 28860
rect 2745 28800 2809 28804
rect 2825 28860 2889 28864
rect 2825 28804 2829 28860
rect 2829 28804 2885 28860
rect 2885 28804 2889 28860
rect 2825 28800 2889 28804
rect 2905 28860 2969 28864
rect 2905 28804 2909 28860
rect 2909 28804 2965 28860
rect 2965 28804 2969 28860
rect 2905 28800 2969 28804
rect 6092 28860 6156 28864
rect 6092 28804 6096 28860
rect 6096 28804 6152 28860
rect 6152 28804 6156 28860
rect 6092 28800 6156 28804
rect 6172 28860 6236 28864
rect 6172 28804 6176 28860
rect 6176 28804 6232 28860
rect 6232 28804 6236 28860
rect 6172 28800 6236 28804
rect 6252 28860 6316 28864
rect 6252 28804 6256 28860
rect 6256 28804 6312 28860
rect 6312 28804 6316 28860
rect 6252 28800 6316 28804
rect 6332 28860 6396 28864
rect 6332 28804 6336 28860
rect 6336 28804 6392 28860
rect 6392 28804 6396 28860
rect 6332 28800 6396 28804
rect 9519 28860 9583 28864
rect 9519 28804 9523 28860
rect 9523 28804 9579 28860
rect 9579 28804 9583 28860
rect 9519 28800 9583 28804
rect 9599 28860 9663 28864
rect 9599 28804 9603 28860
rect 9603 28804 9659 28860
rect 9659 28804 9663 28860
rect 9599 28800 9663 28804
rect 9679 28860 9743 28864
rect 9679 28804 9683 28860
rect 9683 28804 9739 28860
rect 9739 28804 9743 28860
rect 9679 28800 9743 28804
rect 9759 28860 9823 28864
rect 9759 28804 9763 28860
rect 9763 28804 9819 28860
rect 9819 28804 9823 28860
rect 9759 28800 9823 28804
rect 12946 28860 13010 28864
rect 12946 28804 12950 28860
rect 12950 28804 13006 28860
rect 13006 28804 13010 28860
rect 12946 28800 13010 28804
rect 13026 28860 13090 28864
rect 13026 28804 13030 28860
rect 13030 28804 13086 28860
rect 13086 28804 13090 28860
rect 13026 28800 13090 28804
rect 13106 28860 13170 28864
rect 13106 28804 13110 28860
rect 13110 28804 13166 28860
rect 13166 28804 13170 28860
rect 13106 28800 13170 28804
rect 13186 28860 13250 28864
rect 13186 28804 13190 28860
rect 13190 28804 13246 28860
rect 13246 28804 13250 28860
rect 13186 28800 13250 28804
rect 4378 28316 4442 28320
rect 4378 28260 4382 28316
rect 4382 28260 4438 28316
rect 4438 28260 4442 28316
rect 4378 28256 4442 28260
rect 4458 28316 4522 28320
rect 4458 28260 4462 28316
rect 4462 28260 4518 28316
rect 4518 28260 4522 28316
rect 4458 28256 4522 28260
rect 4538 28316 4602 28320
rect 4538 28260 4542 28316
rect 4542 28260 4598 28316
rect 4598 28260 4602 28316
rect 4538 28256 4602 28260
rect 4618 28316 4682 28320
rect 4618 28260 4622 28316
rect 4622 28260 4678 28316
rect 4678 28260 4682 28316
rect 4618 28256 4682 28260
rect 7805 28316 7869 28320
rect 7805 28260 7809 28316
rect 7809 28260 7865 28316
rect 7865 28260 7869 28316
rect 7805 28256 7869 28260
rect 7885 28316 7949 28320
rect 7885 28260 7889 28316
rect 7889 28260 7945 28316
rect 7945 28260 7949 28316
rect 7885 28256 7949 28260
rect 7965 28316 8029 28320
rect 7965 28260 7969 28316
rect 7969 28260 8025 28316
rect 8025 28260 8029 28316
rect 7965 28256 8029 28260
rect 8045 28316 8109 28320
rect 8045 28260 8049 28316
rect 8049 28260 8105 28316
rect 8105 28260 8109 28316
rect 8045 28256 8109 28260
rect 11232 28316 11296 28320
rect 11232 28260 11236 28316
rect 11236 28260 11292 28316
rect 11292 28260 11296 28316
rect 11232 28256 11296 28260
rect 11312 28316 11376 28320
rect 11312 28260 11316 28316
rect 11316 28260 11372 28316
rect 11372 28260 11376 28316
rect 11312 28256 11376 28260
rect 11392 28316 11456 28320
rect 11392 28260 11396 28316
rect 11396 28260 11452 28316
rect 11452 28260 11456 28316
rect 11392 28256 11456 28260
rect 11472 28316 11536 28320
rect 11472 28260 11476 28316
rect 11476 28260 11532 28316
rect 11532 28260 11536 28316
rect 11472 28256 11536 28260
rect 14659 28316 14723 28320
rect 14659 28260 14663 28316
rect 14663 28260 14719 28316
rect 14719 28260 14723 28316
rect 14659 28256 14723 28260
rect 14739 28316 14803 28320
rect 14739 28260 14743 28316
rect 14743 28260 14799 28316
rect 14799 28260 14803 28316
rect 14739 28256 14803 28260
rect 14819 28316 14883 28320
rect 14819 28260 14823 28316
rect 14823 28260 14879 28316
rect 14879 28260 14883 28316
rect 14819 28256 14883 28260
rect 14899 28316 14963 28320
rect 14899 28260 14903 28316
rect 14903 28260 14959 28316
rect 14959 28260 14963 28316
rect 14899 28256 14963 28260
rect 2665 27772 2729 27776
rect 2665 27716 2669 27772
rect 2669 27716 2725 27772
rect 2725 27716 2729 27772
rect 2665 27712 2729 27716
rect 2745 27772 2809 27776
rect 2745 27716 2749 27772
rect 2749 27716 2805 27772
rect 2805 27716 2809 27772
rect 2745 27712 2809 27716
rect 2825 27772 2889 27776
rect 2825 27716 2829 27772
rect 2829 27716 2885 27772
rect 2885 27716 2889 27772
rect 2825 27712 2889 27716
rect 2905 27772 2969 27776
rect 2905 27716 2909 27772
rect 2909 27716 2965 27772
rect 2965 27716 2969 27772
rect 2905 27712 2969 27716
rect 6092 27772 6156 27776
rect 6092 27716 6096 27772
rect 6096 27716 6152 27772
rect 6152 27716 6156 27772
rect 6092 27712 6156 27716
rect 6172 27772 6236 27776
rect 6172 27716 6176 27772
rect 6176 27716 6232 27772
rect 6232 27716 6236 27772
rect 6172 27712 6236 27716
rect 6252 27772 6316 27776
rect 6252 27716 6256 27772
rect 6256 27716 6312 27772
rect 6312 27716 6316 27772
rect 6252 27712 6316 27716
rect 6332 27772 6396 27776
rect 6332 27716 6336 27772
rect 6336 27716 6392 27772
rect 6392 27716 6396 27772
rect 6332 27712 6396 27716
rect 9519 27772 9583 27776
rect 9519 27716 9523 27772
rect 9523 27716 9579 27772
rect 9579 27716 9583 27772
rect 9519 27712 9583 27716
rect 9599 27772 9663 27776
rect 9599 27716 9603 27772
rect 9603 27716 9659 27772
rect 9659 27716 9663 27772
rect 9599 27712 9663 27716
rect 9679 27772 9743 27776
rect 9679 27716 9683 27772
rect 9683 27716 9739 27772
rect 9739 27716 9743 27772
rect 9679 27712 9743 27716
rect 9759 27772 9823 27776
rect 9759 27716 9763 27772
rect 9763 27716 9819 27772
rect 9819 27716 9823 27772
rect 9759 27712 9823 27716
rect 1716 27704 1780 27708
rect 1716 27648 1730 27704
rect 1730 27648 1780 27704
rect 1716 27644 1780 27648
rect 12946 27772 13010 27776
rect 12946 27716 12950 27772
rect 12950 27716 13006 27772
rect 13006 27716 13010 27772
rect 12946 27712 13010 27716
rect 13026 27772 13090 27776
rect 13026 27716 13030 27772
rect 13030 27716 13086 27772
rect 13086 27716 13090 27772
rect 13026 27712 13090 27716
rect 13106 27772 13170 27776
rect 13106 27716 13110 27772
rect 13110 27716 13166 27772
rect 13166 27716 13170 27772
rect 13106 27712 13170 27716
rect 13186 27772 13250 27776
rect 13186 27716 13190 27772
rect 13190 27716 13246 27772
rect 13246 27716 13250 27772
rect 13186 27712 13250 27716
rect 4378 27228 4442 27232
rect 4378 27172 4382 27228
rect 4382 27172 4438 27228
rect 4438 27172 4442 27228
rect 4378 27168 4442 27172
rect 4458 27228 4522 27232
rect 4458 27172 4462 27228
rect 4462 27172 4518 27228
rect 4518 27172 4522 27228
rect 4458 27168 4522 27172
rect 4538 27228 4602 27232
rect 4538 27172 4542 27228
rect 4542 27172 4598 27228
rect 4598 27172 4602 27228
rect 4538 27168 4602 27172
rect 4618 27228 4682 27232
rect 4618 27172 4622 27228
rect 4622 27172 4678 27228
rect 4678 27172 4682 27228
rect 4618 27168 4682 27172
rect 7805 27228 7869 27232
rect 7805 27172 7809 27228
rect 7809 27172 7865 27228
rect 7865 27172 7869 27228
rect 7805 27168 7869 27172
rect 7885 27228 7949 27232
rect 7885 27172 7889 27228
rect 7889 27172 7945 27228
rect 7945 27172 7949 27228
rect 7885 27168 7949 27172
rect 7965 27228 8029 27232
rect 7965 27172 7969 27228
rect 7969 27172 8025 27228
rect 8025 27172 8029 27228
rect 7965 27168 8029 27172
rect 8045 27228 8109 27232
rect 8045 27172 8049 27228
rect 8049 27172 8105 27228
rect 8105 27172 8109 27228
rect 8045 27168 8109 27172
rect 11232 27228 11296 27232
rect 11232 27172 11236 27228
rect 11236 27172 11292 27228
rect 11292 27172 11296 27228
rect 11232 27168 11296 27172
rect 11312 27228 11376 27232
rect 11312 27172 11316 27228
rect 11316 27172 11372 27228
rect 11372 27172 11376 27228
rect 11312 27168 11376 27172
rect 11392 27228 11456 27232
rect 11392 27172 11396 27228
rect 11396 27172 11452 27228
rect 11452 27172 11456 27228
rect 11392 27168 11456 27172
rect 11472 27228 11536 27232
rect 11472 27172 11476 27228
rect 11476 27172 11532 27228
rect 11532 27172 11536 27228
rect 11472 27168 11536 27172
rect 14659 27228 14723 27232
rect 14659 27172 14663 27228
rect 14663 27172 14719 27228
rect 14719 27172 14723 27228
rect 14659 27168 14723 27172
rect 14739 27228 14803 27232
rect 14739 27172 14743 27228
rect 14743 27172 14799 27228
rect 14799 27172 14803 27228
rect 14739 27168 14803 27172
rect 14819 27228 14883 27232
rect 14819 27172 14823 27228
rect 14823 27172 14879 27228
rect 14879 27172 14883 27228
rect 14819 27168 14883 27172
rect 14899 27228 14963 27232
rect 14899 27172 14903 27228
rect 14903 27172 14959 27228
rect 14959 27172 14963 27228
rect 14899 27168 14963 27172
rect 2665 26684 2729 26688
rect 2665 26628 2669 26684
rect 2669 26628 2725 26684
rect 2725 26628 2729 26684
rect 2665 26624 2729 26628
rect 2745 26684 2809 26688
rect 2745 26628 2749 26684
rect 2749 26628 2805 26684
rect 2805 26628 2809 26684
rect 2745 26624 2809 26628
rect 2825 26684 2889 26688
rect 2825 26628 2829 26684
rect 2829 26628 2885 26684
rect 2885 26628 2889 26684
rect 2825 26624 2889 26628
rect 2905 26684 2969 26688
rect 2905 26628 2909 26684
rect 2909 26628 2965 26684
rect 2965 26628 2969 26684
rect 2905 26624 2969 26628
rect 6092 26684 6156 26688
rect 6092 26628 6096 26684
rect 6096 26628 6152 26684
rect 6152 26628 6156 26684
rect 6092 26624 6156 26628
rect 6172 26684 6236 26688
rect 6172 26628 6176 26684
rect 6176 26628 6232 26684
rect 6232 26628 6236 26684
rect 6172 26624 6236 26628
rect 6252 26684 6316 26688
rect 6252 26628 6256 26684
rect 6256 26628 6312 26684
rect 6312 26628 6316 26684
rect 6252 26624 6316 26628
rect 6332 26684 6396 26688
rect 6332 26628 6336 26684
rect 6336 26628 6392 26684
rect 6392 26628 6396 26684
rect 6332 26624 6396 26628
rect 9519 26684 9583 26688
rect 9519 26628 9523 26684
rect 9523 26628 9579 26684
rect 9579 26628 9583 26684
rect 9519 26624 9583 26628
rect 9599 26684 9663 26688
rect 9599 26628 9603 26684
rect 9603 26628 9659 26684
rect 9659 26628 9663 26684
rect 9599 26624 9663 26628
rect 9679 26684 9743 26688
rect 9679 26628 9683 26684
rect 9683 26628 9739 26684
rect 9739 26628 9743 26684
rect 9679 26624 9743 26628
rect 9759 26684 9823 26688
rect 9759 26628 9763 26684
rect 9763 26628 9819 26684
rect 9819 26628 9823 26684
rect 9759 26624 9823 26628
rect 12946 26684 13010 26688
rect 12946 26628 12950 26684
rect 12950 26628 13006 26684
rect 13006 26628 13010 26684
rect 12946 26624 13010 26628
rect 13026 26684 13090 26688
rect 13026 26628 13030 26684
rect 13030 26628 13086 26684
rect 13086 26628 13090 26684
rect 13026 26624 13090 26628
rect 13106 26684 13170 26688
rect 13106 26628 13110 26684
rect 13110 26628 13166 26684
rect 13166 26628 13170 26684
rect 13106 26624 13170 26628
rect 13186 26684 13250 26688
rect 13186 26628 13190 26684
rect 13190 26628 13246 26684
rect 13246 26628 13250 26684
rect 13186 26624 13250 26628
rect 5212 26420 5276 26484
rect 8892 26284 8956 26348
rect 4378 26140 4442 26144
rect 4378 26084 4382 26140
rect 4382 26084 4438 26140
rect 4438 26084 4442 26140
rect 4378 26080 4442 26084
rect 4458 26140 4522 26144
rect 4458 26084 4462 26140
rect 4462 26084 4518 26140
rect 4518 26084 4522 26140
rect 4458 26080 4522 26084
rect 4538 26140 4602 26144
rect 4538 26084 4542 26140
rect 4542 26084 4598 26140
rect 4598 26084 4602 26140
rect 4538 26080 4602 26084
rect 4618 26140 4682 26144
rect 4618 26084 4622 26140
rect 4622 26084 4678 26140
rect 4678 26084 4682 26140
rect 4618 26080 4682 26084
rect 7805 26140 7869 26144
rect 7805 26084 7809 26140
rect 7809 26084 7865 26140
rect 7865 26084 7869 26140
rect 7805 26080 7869 26084
rect 7885 26140 7949 26144
rect 7885 26084 7889 26140
rect 7889 26084 7945 26140
rect 7945 26084 7949 26140
rect 7885 26080 7949 26084
rect 7965 26140 8029 26144
rect 7965 26084 7969 26140
rect 7969 26084 8025 26140
rect 8025 26084 8029 26140
rect 7965 26080 8029 26084
rect 8045 26140 8109 26144
rect 8045 26084 8049 26140
rect 8049 26084 8105 26140
rect 8105 26084 8109 26140
rect 8045 26080 8109 26084
rect 11232 26140 11296 26144
rect 11232 26084 11236 26140
rect 11236 26084 11292 26140
rect 11292 26084 11296 26140
rect 11232 26080 11296 26084
rect 11312 26140 11376 26144
rect 11312 26084 11316 26140
rect 11316 26084 11372 26140
rect 11372 26084 11376 26140
rect 11312 26080 11376 26084
rect 11392 26140 11456 26144
rect 11392 26084 11396 26140
rect 11396 26084 11452 26140
rect 11452 26084 11456 26140
rect 11392 26080 11456 26084
rect 11472 26140 11536 26144
rect 11472 26084 11476 26140
rect 11476 26084 11532 26140
rect 11532 26084 11536 26140
rect 11472 26080 11536 26084
rect 14659 26140 14723 26144
rect 14659 26084 14663 26140
rect 14663 26084 14719 26140
rect 14719 26084 14723 26140
rect 14659 26080 14723 26084
rect 14739 26140 14803 26144
rect 14739 26084 14743 26140
rect 14743 26084 14799 26140
rect 14799 26084 14803 26140
rect 14739 26080 14803 26084
rect 14819 26140 14883 26144
rect 14819 26084 14823 26140
rect 14823 26084 14879 26140
rect 14879 26084 14883 26140
rect 14819 26080 14883 26084
rect 14899 26140 14963 26144
rect 14899 26084 14903 26140
rect 14903 26084 14959 26140
rect 14959 26084 14963 26140
rect 14899 26080 14963 26084
rect 2665 25596 2729 25600
rect 2665 25540 2669 25596
rect 2669 25540 2725 25596
rect 2725 25540 2729 25596
rect 2665 25536 2729 25540
rect 2745 25596 2809 25600
rect 2745 25540 2749 25596
rect 2749 25540 2805 25596
rect 2805 25540 2809 25596
rect 2745 25536 2809 25540
rect 2825 25596 2889 25600
rect 2825 25540 2829 25596
rect 2829 25540 2885 25596
rect 2885 25540 2889 25596
rect 2825 25536 2889 25540
rect 2905 25596 2969 25600
rect 2905 25540 2909 25596
rect 2909 25540 2965 25596
rect 2965 25540 2969 25596
rect 2905 25536 2969 25540
rect 6092 25596 6156 25600
rect 6092 25540 6096 25596
rect 6096 25540 6152 25596
rect 6152 25540 6156 25596
rect 6092 25536 6156 25540
rect 6172 25596 6236 25600
rect 6172 25540 6176 25596
rect 6176 25540 6232 25596
rect 6232 25540 6236 25596
rect 6172 25536 6236 25540
rect 6252 25596 6316 25600
rect 6252 25540 6256 25596
rect 6256 25540 6312 25596
rect 6312 25540 6316 25596
rect 6252 25536 6316 25540
rect 6332 25596 6396 25600
rect 6332 25540 6336 25596
rect 6336 25540 6392 25596
rect 6392 25540 6396 25596
rect 6332 25536 6396 25540
rect 9519 25596 9583 25600
rect 9519 25540 9523 25596
rect 9523 25540 9579 25596
rect 9579 25540 9583 25596
rect 9519 25536 9583 25540
rect 9599 25596 9663 25600
rect 9599 25540 9603 25596
rect 9603 25540 9659 25596
rect 9659 25540 9663 25596
rect 9599 25536 9663 25540
rect 9679 25596 9743 25600
rect 9679 25540 9683 25596
rect 9683 25540 9739 25596
rect 9739 25540 9743 25596
rect 9679 25536 9743 25540
rect 9759 25596 9823 25600
rect 9759 25540 9763 25596
rect 9763 25540 9819 25596
rect 9819 25540 9823 25596
rect 9759 25536 9823 25540
rect 12946 25596 13010 25600
rect 12946 25540 12950 25596
rect 12950 25540 13006 25596
rect 13006 25540 13010 25596
rect 12946 25536 13010 25540
rect 13026 25596 13090 25600
rect 13026 25540 13030 25596
rect 13030 25540 13086 25596
rect 13086 25540 13090 25596
rect 13026 25536 13090 25540
rect 13106 25596 13170 25600
rect 13106 25540 13110 25596
rect 13110 25540 13166 25596
rect 13166 25540 13170 25596
rect 13106 25536 13170 25540
rect 13186 25596 13250 25600
rect 13186 25540 13190 25596
rect 13190 25540 13246 25596
rect 13246 25540 13250 25596
rect 13186 25536 13250 25540
rect 4378 25052 4442 25056
rect 4378 24996 4382 25052
rect 4382 24996 4438 25052
rect 4438 24996 4442 25052
rect 4378 24992 4442 24996
rect 4458 25052 4522 25056
rect 4458 24996 4462 25052
rect 4462 24996 4518 25052
rect 4518 24996 4522 25052
rect 4458 24992 4522 24996
rect 4538 25052 4602 25056
rect 4538 24996 4542 25052
rect 4542 24996 4598 25052
rect 4598 24996 4602 25052
rect 4538 24992 4602 24996
rect 4618 25052 4682 25056
rect 4618 24996 4622 25052
rect 4622 24996 4678 25052
rect 4678 24996 4682 25052
rect 4618 24992 4682 24996
rect 7805 25052 7869 25056
rect 7805 24996 7809 25052
rect 7809 24996 7865 25052
rect 7865 24996 7869 25052
rect 7805 24992 7869 24996
rect 7885 25052 7949 25056
rect 7885 24996 7889 25052
rect 7889 24996 7945 25052
rect 7945 24996 7949 25052
rect 7885 24992 7949 24996
rect 7965 25052 8029 25056
rect 7965 24996 7969 25052
rect 7969 24996 8025 25052
rect 8025 24996 8029 25052
rect 7965 24992 8029 24996
rect 8045 25052 8109 25056
rect 8045 24996 8049 25052
rect 8049 24996 8105 25052
rect 8105 24996 8109 25052
rect 8045 24992 8109 24996
rect 11232 25052 11296 25056
rect 11232 24996 11236 25052
rect 11236 24996 11292 25052
rect 11292 24996 11296 25052
rect 11232 24992 11296 24996
rect 11312 25052 11376 25056
rect 11312 24996 11316 25052
rect 11316 24996 11372 25052
rect 11372 24996 11376 25052
rect 11312 24992 11376 24996
rect 11392 25052 11456 25056
rect 11392 24996 11396 25052
rect 11396 24996 11452 25052
rect 11452 24996 11456 25052
rect 11392 24992 11456 24996
rect 11472 25052 11536 25056
rect 11472 24996 11476 25052
rect 11476 24996 11532 25052
rect 11532 24996 11536 25052
rect 11472 24992 11536 24996
rect 14659 25052 14723 25056
rect 14659 24996 14663 25052
rect 14663 24996 14719 25052
rect 14719 24996 14723 25052
rect 14659 24992 14723 24996
rect 14739 25052 14803 25056
rect 14739 24996 14743 25052
rect 14743 24996 14799 25052
rect 14799 24996 14803 25052
rect 14739 24992 14803 24996
rect 14819 25052 14883 25056
rect 14819 24996 14823 25052
rect 14823 24996 14879 25052
rect 14879 24996 14883 25052
rect 14819 24992 14883 24996
rect 14899 25052 14963 25056
rect 14899 24996 14903 25052
rect 14903 24996 14959 25052
rect 14959 24996 14963 25052
rect 14899 24992 14963 24996
rect 2665 24508 2729 24512
rect 2665 24452 2669 24508
rect 2669 24452 2725 24508
rect 2725 24452 2729 24508
rect 2665 24448 2729 24452
rect 2745 24508 2809 24512
rect 2745 24452 2749 24508
rect 2749 24452 2805 24508
rect 2805 24452 2809 24508
rect 2745 24448 2809 24452
rect 2825 24508 2889 24512
rect 2825 24452 2829 24508
rect 2829 24452 2885 24508
rect 2885 24452 2889 24508
rect 2825 24448 2889 24452
rect 2905 24508 2969 24512
rect 2905 24452 2909 24508
rect 2909 24452 2965 24508
rect 2965 24452 2969 24508
rect 2905 24448 2969 24452
rect 6092 24508 6156 24512
rect 6092 24452 6096 24508
rect 6096 24452 6152 24508
rect 6152 24452 6156 24508
rect 6092 24448 6156 24452
rect 6172 24508 6236 24512
rect 6172 24452 6176 24508
rect 6176 24452 6232 24508
rect 6232 24452 6236 24508
rect 6172 24448 6236 24452
rect 6252 24508 6316 24512
rect 6252 24452 6256 24508
rect 6256 24452 6312 24508
rect 6312 24452 6316 24508
rect 6252 24448 6316 24452
rect 6332 24508 6396 24512
rect 6332 24452 6336 24508
rect 6336 24452 6392 24508
rect 6392 24452 6396 24508
rect 6332 24448 6396 24452
rect 9519 24508 9583 24512
rect 9519 24452 9523 24508
rect 9523 24452 9579 24508
rect 9579 24452 9583 24508
rect 9519 24448 9583 24452
rect 9599 24508 9663 24512
rect 9599 24452 9603 24508
rect 9603 24452 9659 24508
rect 9659 24452 9663 24508
rect 9599 24448 9663 24452
rect 9679 24508 9743 24512
rect 9679 24452 9683 24508
rect 9683 24452 9739 24508
rect 9739 24452 9743 24508
rect 9679 24448 9743 24452
rect 9759 24508 9823 24512
rect 9759 24452 9763 24508
rect 9763 24452 9819 24508
rect 9819 24452 9823 24508
rect 9759 24448 9823 24452
rect 12946 24508 13010 24512
rect 12946 24452 12950 24508
rect 12950 24452 13006 24508
rect 13006 24452 13010 24508
rect 12946 24448 13010 24452
rect 13026 24508 13090 24512
rect 13026 24452 13030 24508
rect 13030 24452 13086 24508
rect 13086 24452 13090 24508
rect 13026 24448 13090 24452
rect 13106 24508 13170 24512
rect 13106 24452 13110 24508
rect 13110 24452 13166 24508
rect 13166 24452 13170 24508
rect 13106 24448 13170 24452
rect 13186 24508 13250 24512
rect 13186 24452 13190 24508
rect 13190 24452 13246 24508
rect 13246 24452 13250 24508
rect 13186 24448 13250 24452
rect 4378 23964 4442 23968
rect 4378 23908 4382 23964
rect 4382 23908 4438 23964
rect 4438 23908 4442 23964
rect 4378 23904 4442 23908
rect 4458 23964 4522 23968
rect 4458 23908 4462 23964
rect 4462 23908 4518 23964
rect 4518 23908 4522 23964
rect 4458 23904 4522 23908
rect 4538 23964 4602 23968
rect 4538 23908 4542 23964
rect 4542 23908 4598 23964
rect 4598 23908 4602 23964
rect 4538 23904 4602 23908
rect 4618 23964 4682 23968
rect 4618 23908 4622 23964
rect 4622 23908 4678 23964
rect 4678 23908 4682 23964
rect 4618 23904 4682 23908
rect 7805 23964 7869 23968
rect 7805 23908 7809 23964
rect 7809 23908 7865 23964
rect 7865 23908 7869 23964
rect 7805 23904 7869 23908
rect 7885 23964 7949 23968
rect 7885 23908 7889 23964
rect 7889 23908 7945 23964
rect 7945 23908 7949 23964
rect 7885 23904 7949 23908
rect 7965 23964 8029 23968
rect 7965 23908 7969 23964
rect 7969 23908 8025 23964
rect 8025 23908 8029 23964
rect 7965 23904 8029 23908
rect 8045 23964 8109 23968
rect 8045 23908 8049 23964
rect 8049 23908 8105 23964
rect 8105 23908 8109 23964
rect 8045 23904 8109 23908
rect 11232 23964 11296 23968
rect 11232 23908 11236 23964
rect 11236 23908 11292 23964
rect 11292 23908 11296 23964
rect 11232 23904 11296 23908
rect 11312 23964 11376 23968
rect 11312 23908 11316 23964
rect 11316 23908 11372 23964
rect 11372 23908 11376 23964
rect 11312 23904 11376 23908
rect 11392 23964 11456 23968
rect 11392 23908 11396 23964
rect 11396 23908 11452 23964
rect 11452 23908 11456 23964
rect 11392 23904 11456 23908
rect 11472 23964 11536 23968
rect 11472 23908 11476 23964
rect 11476 23908 11532 23964
rect 11532 23908 11536 23964
rect 11472 23904 11536 23908
rect 14659 23964 14723 23968
rect 14659 23908 14663 23964
rect 14663 23908 14719 23964
rect 14719 23908 14723 23964
rect 14659 23904 14723 23908
rect 14739 23964 14803 23968
rect 14739 23908 14743 23964
rect 14743 23908 14799 23964
rect 14799 23908 14803 23964
rect 14739 23904 14803 23908
rect 14819 23964 14883 23968
rect 14819 23908 14823 23964
rect 14823 23908 14879 23964
rect 14879 23908 14883 23964
rect 14819 23904 14883 23908
rect 14899 23964 14963 23968
rect 14899 23908 14903 23964
rect 14903 23908 14959 23964
rect 14959 23908 14963 23964
rect 14899 23904 14963 23908
rect 13492 23836 13556 23900
rect 2665 23420 2729 23424
rect 2665 23364 2669 23420
rect 2669 23364 2725 23420
rect 2725 23364 2729 23420
rect 2665 23360 2729 23364
rect 2745 23420 2809 23424
rect 2745 23364 2749 23420
rect 2749 23364 2805 23420
rect 2805 23364 2809 23420
rect 2745 23360 2809 23364
rect 2825 23420 2889 23424
rect 2825 23364 2829 23420
rect 2829 23364 2885 23420
rect 2885 23364 2889 23420
rect 2825 23360 2889 23364
rect 2905 23420 2969 23424
rect 2905 23364 2909 23420
rect 2909 23364 2965 23420
rect 2965 23364 2969 23420
rect 2905 23360 2969 23364
rect 6092 23420 6156 23424
rect 6092 23364 6096 23420
rect 6096 23364 6152 23420
rect 6152 23364 6156 23420
rect 6092 23360 6156 23364
rect 6172 23420 6236 23424
rect 6172 23364 6176 23420
rect 6176 23364 6232 23420
rect 6232 23364 6236 23420
rect 6172 23360 6236 23364
rect 6252 23420 6316 23424
rect 6252 23364 6256 23420
rect 6256 23364 6312 23420
rect 6312 23364 6316 23420
rect 6252 23360 6316 23364
rect 6332 23420 6396 23424
rect 6332 23364 6336 23420
rect 6336 23364 6392 23420
rect 6392 23364 6396 23420
rect 6332 23360 6396 23364
rect 9519 23420 9583 23424
rect 9519 23364 9523 23420
rect 9523 23364 9579 23420
rect 9579 23364 9583 23420
rect 9519 23360 9583 23364
rect 9599 23420 9663 23424
rect 9599 23364 9603 23420
rect 9603 23364 9659 23420
rect 9659 23364 9663 23420
rect 9599 23360 9663 23364
rect 9679 23420 9743 23424
rect 9679 23364 9683 23420
rect 9683 23364 9739 23420
rect 9739 23364 9743 23420
rect 9679 23360 9743 23364
rect 9759 23420 9823 23424
rect 9759 23364 9763 23420
rect 9763 23364 9819 23420
rect 9819 23364 9823 23420
rect 9759 23360 9823 23364
rect 12946 23420 13010 23424
rect 12946 23364 12950 23420
rect 12950 23364 13006 23420
rect 13006 23364 13010 23420
rect 12946 23360 13010 23364
rect 13026 23420 13090 23424
rect 13026 23364 13030 23420
rect 13030 23364 13086 23420
rect 13086 23364 13090 23420
rect 13026 23360 13090 23364
rect 13106 23420 13170 23424
rect 13106 23364 13110 23420
rect 13110 23364 13166 23420
rect 13166 23364 13170 23420
rect 13106 23360 13170 23364
rect 13186 23420 13250 23424
rect 13186 23364 13190 23420
rect 13190 23364 13246 23420
rect 13246 23364 13250 23420
rect 13186 23360 13250 23364
rect 4378 22876 4442 22880
rect 4378 22820 4382 22876
rect 4382 22820 4438 22876
rect 4438 22820 4442 22876
rect 4378 22816 4442 22820
rect 4458 22876 4522 22880
rect 4458 22820 4462 22876
rect 4462 22820 4518 22876
rect 4518 22820 4522 22876
rect 4458 22816 4522 22820
rect 4538 22876 4602 22880
rect 4538 22820 4542 22876
rect 4542 22820 4598 22876
rect 4598 22820 4602 22876
rect 4538 22816 4602 22820
rect 4618 22876 4682 22880
rect 4618 22820 4622 22876
rect 4622 22820 4678 22876
rect 4678 22820 4682 22876
rect 4618 22816 4682 22820
rect 7805 22876 7869 22880
rect 7805 22820 7809 22876
rect 7809 22820 7865 22876
rect 7865 22820 7869 22876
rect 7805 22816 7869 22820
rect 7885 22876 7949 22880
rect 7885 22820 7889 22876
rect 7889 22820 7945 22876
rect 7945 22820 7949 22876
rect 7885 22816 7949 22820
rect 7965 22876 8029 22880
rect 7965 22820 7969 22876
rect 7969 22820 8025 22876
rect 8025 22820 8029 22876
rect 7965 22816 8029 22820
rect 8045 22876 8109 22880
rect 8045 22820 8049 22876
rect 8049 22820 8105 22876
rect 8105 22820 8109 22876
rect 8045 22816 8109 22820
rect 11232 22876 11296 22880
rect 11232 22820 11236 22876
rect 11236 22820 11292 22876
rect 11292 22820 11296 22876
rect 11232 22816 11296 22820
rect 11312 22876 11376 22880
rect 11312 22820 11316 22876
rect 11316 22820 11372 22876
rect 11372 22820 11376 22876
rect 11312 22816 11376 22820
rect 11392 22876 11456 22880
rect 11392 22820 11396 22876
rect 11396 22820 11452 22876
rect 11452 22820 11456 22876
rect 11392 22816 11456 22820
rect 11472 22876 11536 22880
rect 11472 22820 11476 22876
rect 11476 22820 11532 22876
rect 11532 22820 11536 22876
rect 11472 22816 11536 22820
rect 14659 22876 14723 22880
rect 14659 22820 14663 22876
rect 14663 22820 14719 22876
rect 14719 22820 14723 22876
rect 14659 22816 14723 22820
rect 14739 22876 14803 22880
rect 14739 22820 14743 22876
rect 14743 22820 14799 22876
rect 14799 22820 14803 22876
rect 14739 22816 14803 22820
rect 14819 22876 14883 22880
rect 14819 22820 14823 22876
rect 14823 22820 14879 22876
rect 14879 22820 14883 22876
rect 14819 22816 14883 22820
rect 14899 22876 14963 22880
rect 14899 22820 14903 22876
rect 14903 22820 14959 22876
rect 14959 22820 14963 22876
rect 14899 22816 14963 22820
rect 13860 22340 13924 22404
rect 2665 22332 2729 22336
rect 2665 22276 2669 22332
rect 2669 22276 2725 22332
rect 2725 22276 2729 22332
rect 2665 22272 2729 22276
rect 2745 22332 2809 22336
rect 2745 22276 2749 22332
rect 2749 22276 2805 22332
rect 2805 22276 2809 22332
rect 2745 22272 2809 22276
rect 2825 22332 2889 22336
rect 2825 22276 2829 22332
rect 2829 22276 2885 22332
rect 2885 22276 2889 22332
rect 2825 22272 2889 22276
rect 2905 22332 2969 22336
rect 2905 22276 2909 22332
rect 2909 22276 2965 22332
rect 2965 22276 2969 22332
rect 2905 22272 2969 22276
rect 6092 22332 6156 22336
rect 6092 22276 6096 22332
rect 6096 22276 6152 22332
rect 6152 22276 6156 22332
rect 6092 22272 6156 22276
rect 6172 22332 6236 22336
rect 6172 22276 6176 22332
rect 6176 22276 6232 22332
rect 6232 22276 6236 22332
rect 6172 22272 6236 22276
rect 6252 22332 6316 22336
rect 6252 22276 6256 22332
rect 6256 22276 6312 22332
rect 6312 22276 6316 22332
rect 6252 22272 6316 22276
rect 6332 22332 6396 22336
rect 6332 22276 6336 22332
rect 6336 22276 6392 22332
rect 6392 22276 6396 22332
rect 6332 22272 6396 22276
rect 9519 22332 9583 22336
rect 9519 22276 9523 22332
rect 9523 22276 9579 22332
rect 9579 22276 9583 22332
rect 9519 22272 9583 22276
rect 9599 22332 9663 22336
rect 9599 22276 9603 22332
rect 9603 22276 9659 22332
rect 9659 22276 9663 22332
rect 9599 22272 9663 22276
rect 9679 22332 9743 22336
rect 9679 22276 9683 22332
rect 9683 22276 9739 22332
rect 9739 22276 9743 22332
rect 9679 22272 9743 22276
rect 9759 22332 9823 22336
rect 9759 22276 9763 22332
rect 9763 22276 9819 22332
rect 9819 22276 9823 22332
rect 9759 22272 9823 22276
rect 12946 22332 13010 22336
rect 12946 22276 12950 22332
rect 12950 22276 13006 22332
rect 13006 22276 13010 22332
rect 12946 22272 13010 22276
rect 13026 22332 13090 22336
rect 13026 22276 13030 22332
rect 13030 22276 13086 22332
rect 13086 22276 13090 22332
rect 13026 22272 13090 22276
rect 13106 22332 13170 22336
rect 13106 22276 13110 22332
rect 13110 22276 13166 22332
rect 13166 22276 13170 22332
rect 13106 22272 13170 22276
rect 13186 22332 13250 22336
rect 13186 22276 13190 22332
rect 13190 22276 13246 22332
rect 13246 22276 13250 22332
rect 13186 22272 13250 22276
rect 11836 21932 11900 21996
rect 12572 21932 12636 21996
rect 15332 21992 15396 21996
rect 15332 21936 15382 21992
rect 15382 21936 15396 21992
rect 15332 21932 15396 21936
rect 4378 21788 4442 21792
rect 4378 21732 4382 21788
rect 4382 21732 4438 21788
rect 4438 21732 4442 21788
rect 4378 21728 4442 21732
rect 4458 21788 4522 21792
rect 4458 21732 4462 21788
rect 4462 21732 4518 21788
rect 4518 21732 4522 21788
rect 4458 21728 4522 21732
rect 4538 21788 4602 21792
rect 4538 21732 4542 21788
rect 4542 21732 4598 21788
rect 4598 21732 4602 21788
rect 4538 21728 4602 21732
rect 4618 21788 4682 21792
rect 4618 21732 4622 21788
rect 4622 21732 4678 21788
rect 4678 21732 4682 21788
rect 4618 21728 4682 21732
rect 7805 21788 7869 21792
rect 7805 21732 7809 21788
rect 7809 21732 7865 21788
rect 7865 21732 7869 21788
rect 7805 21728 7869 21732
rect 7885 21788 7949 21792
rect 7885 21732 7889 21788
rect 7889 21732 7945 21788
rect 7945 21732 7949 21788
rect 7885 21728 7949 21732
rect 7965 21788 8029 21792
rect 7965 21732 7969 21788
rect 7969 21732 8025 21788
rect 8025 21732 8029 21788
rect 7965 21728 8029 21732
rect 8045 21788 8109 21792
rect 8045 21732 8049 21788
rect 8049 21732 8105 21788
rect 8105 21732 8109 21788
rect 8045 21728 8109 21732
rect 11232 21788 11296 21792
rect 11232 21732 11236 21788
rect 11236 21732 11292 21788
rect 11292 21732 11296 21788
rect 11232 21728 11296 21732
rect 11312 21788 11376 21792
rect 11312 21732 11316 21788
rect 11316 21732 11372 21788
rect 11372 21732 11376 21788
rect 11312 21728 11376 21732
rect 11392 21788 11456 21792
rect 11392 21732 11396 21788
rect 11396 21732 11452 21788
rect 11452 21732 11456 21788
rect 11392 21728 11456 21732
rect 11472 21788 11536 21792
rect 11472 21732 11476 21788
rect 11476 21732 11532 21788
rect 11532 21732 11536 21788
rect 11472 21728 11536 21732
rect 14659 21788 14723 21792
rect 14659 21732 14663 21788
rect 14663 21732 14719 21788
rect 14719 21732 14723 21788
rect 14659 21728 14723 21732
rect 14739 21788 14803 21792
rect 14739 21732 14743 21788
rect 14743 21732 14799 21788
rect 14799 21732 14803 21788
rect 14739 21728 14803 21732
rect 14819 21788 14883 21792
rect 14819 21732 14823 21788
rect 14823 21732 14879 21788
rect 14879 21732 14883 21788
rect 14819 21728 14883 21732
rect 14899 21788 14963 21792
rect 14899 21732 14903 21788
rect 14903 21732 14959 21788
rect 14959 21732 14963 21788
rect 14899 21728 14963 21732
rect 2665 21244 2729 21248
rect 2665 21188 2669 21244
rect 2669 21188 2725 21244
rect 2725 21188 2729 21244
rect 2665 21184 2729 21188
rect 2745 21244 2809 21248
rect 2745 21188 2749 21244
rect 2749 21188 2805 21244
rect 2805 21188 2809 21244
rect 2745 21184 2809 21188
rect 2825 21244 2889 21248
rect 2825 21188 2829 21244
rect 2829 21188 2885 21244
rect 2885 21188 2889 21244
rect 2825 21184 2889 21188
rect 2905 21244 2969 21248
rect 2905 21188 2909 21244
rect 2909 21188 2965 21244
rect 2965 21188 2969 21244
rect 2905 21184 2969 21188
rect 6092 21244 6156 21248
rect 6092 21188 6096 21244
rect 6096 21188 6152 21244
rect 6152 21188 6156 21244
rect 6092 21184 6156 21188
rect 6172 21244 6236 21248
rect 6172 21188 6176 21244
rect 6176 21188 6232 21244
rect 6232 21188 6236 21244
rect 6172 21184 6236 21188
rect 6252 21244 6316 21248
rect 6252 21188 6256 21244
rect 6256 21188 6312 21244
rect 6312 21188 6316 21244
rect 6252 21184 6316 21188
rect 6332 21244 6396 21248
rect 6332 21188 6336 21244
rect 6336 21188 6392 21244
rect 6392 21188 6396 21244
rect 6332 21184 6396 21188
rect 9519 21244 9583 21248
rect 9519 21188 9523 21244
rect 9523 21188 9579 21244
rect 9579 21188 9583 21244
rect 9519 21184 9583 21188
rect 9599 21244 9663 21248
rect 9599 21188 9603 21244
rect 9603 21188 9659 21244
rect 9659 21188 9663 21244
rect 9599 21184 9663 21188
rect 9679 21244 9743 21248
rect 9679 21188 9683 21244
rect 9683 21188 9739 21244
rect 9739 21188 9743 21244
rect 9679 21184 9743 21188
rect 9759 21244 9823 21248
rect 9759 21188 9763 21244
rect 9763 21188 9819 21244
rect 9819 21188 9823 21244
rect 9759 21184 9823 21188
rect 12946 21244 13010 21248
rect 12946 21188 12950 21244
rect 12950 21188 13006 21244
rect 13006 21188 13010 21244
rect 12946 21184 13010 21188
rect 13026 21244 13090 21248
rect 13026 21188 13030 21244
rect 13030 21188 13086 21244
rect 13086 21188 13090 21244
rect 13026 21184 13090 21188
rect 13106 21244 13170 21248
rect 13106 21188 13110 21244
rect 13110 21188 13166 21244
rect 13166 21188 13170 21244
rect 13106 21184 13170 21188
rect 13186 21244 13250 21248
rect 13186 21188 13190 21244
rect 13190 21188 13246 21244
rect 13246 21188 13250 21244
rect 13186 21184 13250 21188
rect 13492 21176 13556 21180
rect 13492 21120 13542 21176
rect 13542 21120 13556 21176
rect 13492 21116 13556 21120
rect 4378 20700 4442 20704
rect 4378 20644 4382 20700
rect 4382 20644 4438 20700
rect 4438 20644 4442 20700
rect 4378 20640 4442 20644
rect 4458 20700 4522 20704
rect 4458 20644 4462 20700
rect 4462 20644 4518 20700
rect 4518 20644 4522 20700
rect 4458 20640 4522 20644
rect 4538 20700 4602 20704
rect 4538 20644 4542 20700
rect 4542 20644 4598 20700
rect 4598 20644 4602 20700
rect 4538 20640 4602 20644
rect 4618 20700 4682 20704
rect 4618 20644 4622 20700
rect 4622 20644 4678 20700
rect 4678 20644 4682 20700
rect 4618 20640 4682 20644
rect 7805 20700 7869 20704
rect 7805 20644 7809 20700
rect 7809 20644 7865 20700
rect 7865 20644 7869 20700
rect 7805 20640 7869 20644
rect 7885 20700 7949 20704
rect 7885 20644 7889 20700
rect 7889 20644 7945 20700
rect 7945 20644 7949 20700
rect 7885 20640 7949 20644
rect 7965 20700 8029 20704
rect 7965 20644 7969 20700
rect 7969 20644 8025 20700
rect 8025 20644 8029 20700
rect 7965 20640 8029 20644
rect 8045 20700 8109 20704
rect 8045 20644 8049 20700
rect 8049 20644 8105 20700
rect 8105 20644 8109 20700
rect 8045 20640 8109 20644
rect 12756 20708 12820 20772
rect 11232 20700 11296 20704
rect 11232 20644 11236 20700
rect 11236 20644 11292 20700
rect 11292 20644 11296 20700
rect 11232 20640 11296 20644
rect 11312 20700 11376 20704
rect 11312 20644 11316 20700
rect 11316 20644 11372 20700
rect 11372 20644 11376 20700
rect 11312 20640 11376 20644
rect 11392 20700 11456 20704
rect 11392 20644 11396 20700
rect 11396 20644 11452 20700
rect 11452 20644 11456 20700
rect 11392 20640 11456 20644
rect 11472 20700 11536 20704
rect 11472 20644 11476 20700
rect 11476 20644 11532 20700
rect 11532 20644 11536 20700
rect 11472 20640 11536 20644
rect 14659 20700 14723 20704
rect 14659 20644 14663 20700
rect 14663 20644 14719 20700
rect 14719 20644 14723 20700
rect 14659 20640 14723 20644
rect 14739 20700 14803 20704
rect 14739 20644 14743 20700
rect 14743 20644 14799 20700
rect 14799 20644 14803 20700
rect 14739 20640 14803 20644
rect 14819 20700 14883 20704
rect 14819 20644 14823 20700
rect 14823 20644 14879 20700
rect 14879 20644 14883 20700
rect 14819 20640 14883 20644
rect 14899 20700 14963 20704
rect 14899 20644 14903 20700
rect 14903 20644 14959 20700
rect 14959 20644 14963 20700
rect 14899 20640 14963 20644
rect 8708 20436 8772 20500
rect 7236 20360 7300 20364
rect 7236 20304 7286 20360
rect 7286 20304 7300 20360
rect 7236 20300 7300 20304
rect 2665 20156 2729 20160
rect 2665 20100 2669 20156
rect 2669 20100 2725 20156
rect 2725 20100 2729 20156
rect 2665 20096 2729 20100
rect 2745 20156 2809 20160
rect 2745 20100 2749 20156
rect 2749 20100 2805 20156
rect 2805 20100 2809 20156
rect 2745 20096 2809 20100
rect 2825 20156 2889 20160
rect 2825 20100 2829 20156
rect 2829 20100 2885 20156
rect 2885 20100 2889 20156
rect 2825 20096 2889 20100
rect 2905 20156 2969 20160
rect 2905 20100 2909 20156
rect 2909 20100 2965 20156
rect 2965 20100 2969 20156
rect 2905 20096 2969 20100
rect 6092 20156 6156 20160
rect 6092 20100 6096 20156
rect 6096 20100 6152 20156
rect 6152 20100 6156 20156
rect 6092 20096 6156 20100
rect 6172 20156 6236 20160
rect 6172 20100 6176 20156
rect 6176 20100 6232 20156
rect 6232 20100 6236 20156
rect 6172 20096 6236 20100
rect 6252 20156 6316 20160
rect 6252 20100 6256 20156
rect 6256 20100 6312 20156
rect 6312 20100 6316 20156
rect 6252 20096 6316 20100
rect 6332 20156 6396 20160
rect 6332 20100 6336 20156
rect 6336 20100 6392 20156
rect 6392 20100 6396 20156
rect 6332 20096 6396 20100
rect 9519 20156 9583 20160
rect 9519 20100 9523 20156
rect 9523 20100 9579 20156
rect 9579 20100 9583 20156
rect 9519 20096 9583 20100
rect 9599 20156 9663 20160
rect 9599 20100 9603 20156
rect 9603 20100 9659 20156
rect 9659 20100 9663 20156
rect 9599 20096 9663 20100
rect 9679 20156 9743 20160
rect 9679 20100 9683 20156
rect 9683 20100 9739 20156
rect 9739 20100 9743 20156
rect 9679 20096 9743 20100
rect 9759 20156 9823 20160
rect 9759 20100 9763 20156
rect 9763 20100 9819 20156
rect 9819 20100 9823 20156
rect 9759 20096 9823 20100
rect 12946 20156 13010 20160
rect 12946 20100 12950 20156
rect 12950 20100 13006 20156
rect 13006 20100 13010 20156
rect 12946 20096 13010 20100
rect 13026 20156 13090 20160
rect 13026 20100 13030 20156
rect 13030 20100 13086 20156
rect 13086 20100 13090 20156
rect 13026 20096 13090 20100
rect 13106 20156 13170 20160
rect 13106 20100 13110 20156
rect 13110 20100 13166 20156
rect 13166 20100 13170 20156
rect 13106 20096 13170 20100
rect 13186 20156 13250 20160
rect 13186 20100 13190 20156
rect 13190 20100 13246 20156
rect 13246 20100 13250 20156
rect 13186 20096 13250 20100
rect 9076 20028 9140 20092
rect 9260 19892 9324 19956
rect 8708 19756 8772 19820
rect 9076 19680 9140 19684
rect 9076 19624 9126 19680
rect 9126 19624 9140 19680
rect 9076 19620 9140 19624
rect 4378 19612 4442 19616
rect 4378 19556 4382 19612
rect 4382 19556 4438 19612
rect 4438 19556 4442 19612
rect 4378 19552 4442 19556
rect 4458 19612 4522 19616
rect 4458 19556 4462 19612
rect 4462 19556 4518 19612
rect 4518 19556 4522 19612
rect 4458 19552 4522 19556
rect 4538 19612 4602 19616
rect 4538 19556 4542 19612
rect 4542 19556 4598 19612
rect 4598 19556 4602 19612
rect 4538 19552 4602 19556
rect 4618 19612 4682 19616
rect 4618 19556 4622 19612
rect 4622 19556 4678 19612
rect 4678 19556 4682 19612
rect 4618 19552 4682 19556
rect 7805 19612 7869 19616
rect 7805 19556 7809 19612
rect 7809 19556 7865 19612
rect 7865 19556 7869 19612
rect 7805 19552 7869 19556
rect 7885 19612 7949 19616
rect 7885 19556 7889 19612
rect 7889 19556 7945 19612
rect 7945 19556 7949 19612
rect 7885 19552 7949 19556
rect 7965 19612 8029 19616
rect 7965 19556 7969 19612
rect 7969 19556 8025 19612
rect 8025 19556 8029 19612
rect 7965 19552 8029 19556
rect 8045 19612 8109 19616
rect 8045 19556 8049 19612
rect 8049 19556 8105 19612
rect 8105 19556 8109 19612
rect 8045 19552 8109 19556
rect 11232 19612 11296 19616
rect 11232 19556 11236 19612
rect 11236 19556 11292 19612
rect 11292 19556 11296 19612
rect 11232 19552 11296 19556
rect 11312 19612 11376 19616
rect 11312 19556 11316 19612
rect 11316 19556 11372 19612
rect 11372 19556 11376 19612
rect 11312 19552 11376 19556
rect 11392 19612 11456 19616
rect 11392 19556 11396 19612
rect 11396 19556 11452 19612
rect 11452 19556 11456 19612
rect 11392 19552 11456 19556
rect 11472 19612 11536 19616
rect 11472 19556 11476 19612
rect 11476 19556 11532 19612
rect 11532 19556 11536 19612
rect 11472 19552 11536 19556
rect 14659 19612 14723 19616
rect 14659 19556 14663 19612
rect 14663 19556 14719 19612
rect 14719 19556 14723 19612
rect 14659 19552 14723 19556
rect 14739 19612 14803 19616
rect 14739 19556 14743 19612
rect 14743 19556 14799 19612
rect 14799 19556 14803 19612
rect 14739 19552 14803 19556
rect 14819 19612 14883 19616
rect 14819 19556 14823 19612
rect 14823 19556 14879 19612
rect 14879 19556 14883 19612
rect 14819 19552 14883 19556
rect 14899 19612 14963 19616
rect 14899 19556 14903 19612
rect 14903 19556 14959 19612
rect 14959 19556 14963 19612
rect 14899 19552 14963 19556
rect 10548 19272 10612 19276
rect 10548 19216 10562 19272
rect 10562 19216 10612 19272
rect 10548 19212 10612 19216
rect 2665 19068 2729 19072
rect 2665 19012 2669 19068
rect 2669 19012 2725 19068
rect 2725 19012 2729 19068
rect 2665 19008 2729 19012
rect 2745 19068 2809 19072
rect 2745 19012 2749 19068
rect 2749 19012 2805 19068
rect 2805 19012 2809 19068
rect 2745 19008 2809 19012
rect 2825 19068 2889 19072
rect 2825 19012 2829 19068
rect 2829 19012 2885 19068
rect 2885 19012 2889 19068
rect 2825 19008 2889 19012
rect 2905 19068 2969 19072
rect 2905 19012 2909 19068
rect 2909 19012 2965 19068
rect 2965 19012 2969 19068
rect 2905 19008 2969 19012
rect 6092 19068 6156 19072
rect 6092 19012 6096 19068
rect 6096 19012 6152 19068
rect 6152 19012 6156 19068
rect 6092 19008 6156 19012
rect 6172 19068 6236 19072
rect 6172 19012 6176 19068
rect 6176 19012 6232 19068
rect 6232 19012 6236 19068
rect 6172 19008 6236 19012
rect 6252 19068 6316 19072
rect 6252 19012 6256 19068
rect 6256 19012 6312 19068
rect 6312 19012 6316 19068
rect 6252 19008 6316 19012
rect 6332 19068 6396 19072
rect 6332 19012 6336 19068
rect 6336 19012 6392 19068
rect 6392 19012 6396 19068
rect 6332 19008 6396 19012
rect 9519 19068 9583 19072
rect 9519 19012 9523 19068
rect 9523 19012 9579 19068
rect 9579 19012 9583 19068
rect 9519 19008 9583 19012
rect 9599 19068 9663 19072
rect 9599 19012 9603 19068
rect 9603 19012 9659 19068
rect 9659 19012 9663 19068
rect 9599 19008 9663 19012
rect 9679 19068 9743 19072
rect 9679 19012 9683 19068
rect 9683 19012 9739 19068
rect 9739 19012 9743 19068
rect 9679 19008 9743 19012
rect 9759 19068 9823 19072
rect 9759 19012 9763 19068
rect 9763 19012 9819 19068
rect 9819 19012 9823 19068
rect 9759 19008 9823 19012
rect 12946 19068 13010 19072
rect 12946 19012 12950 19068
rect 12950 19012 13006 19068
rect 13006 19012 13010 19068
rect 12946 19008 13010 19012
rect 13026 19068 13090 19072
rect 13026 19012 13030 19068
rect 13030 19012 13086 19068
rect 13086 19012 13090 19068
rect 13026 19008 13090 19012
rect 13106 19068 13170 19072
rect 13106 19012 13110 19068
rect 13110 19012 13166 19068
rect 13166 19012 13170 19068
rect 13106 19008 13170 19012
rect 13186 19068 13250 19072
rect 13186 19012 13190 19068
rect 13190 19012 13246 19068
rect 13246 19012 13250 19068
rect 13186 19008 13250 19012
rect 4378 18524 4442 18528
rect 4378 18468 4382 18524
rect 4382 18468 4438 18524
rect 4438 18468 4442 18524
rect 4378 18464 4442 18468
rect 4458 18524 4522 18528
rect 4458 18468 4462 18524
rect 4462 18468 4518 18524
rect 4518 18468 4522 18524
rect 4458 18464 4522 18468
rect 4538 18524 4602 18528
rect 4538 18468 4542 18524
rect 4542 18468 4598 18524
rect 4598 18468 4602 18524
rect 4538 18464 4602 18468
rect 4618 18524 4682 18528
rect 4618 18468 4622 18524
rect 4622 18468 4678 18524
rect 4678 18468 4682 18524
rect 4618 18464 4682 18468
rect 7805 18524 7869 18528
rect 7805 18468 7809 18524
rect 7809 18468 7865 18524
rect 7865 18468 7869 18524
rect 7805 18464 7869 18468
rect 7885 18524 7949 18528
rect 7885 18468 7889 18524
rect 7889 18468 7945 18524
rect 7945 18468 7949 18524
rect 7885 18464 7949 18468
rect 7965 18524 8029 18528
rect 7965 18468 7969 18524
rect 7969 18468 8025 18524
rect 8025 18468 8029 18524
rect 7965 18464 8029 18468
rect 8045 18524 8109 18528
rect 8045 18468 8049 18524
rect 8049 18468 8105 18524
rect 8105 18468 8109 18524
rect 8045 18464 8109 18468
rect 11232 18524 11296 18528
rect 11232 18468 11236 18524
rect 11236 18468 11292 18524
rect 11292 18468 11296 18524
rect 11232 18464 11296 18468
rect 11312 18524 11376 18528
rect 11312 18468 11316 18524
rect 11316 18468 11372 18524
rect 11372 18468 11376 18524
rect 11312 18464 11376 18468
rect 11392 18524 11456 18528
rect 11392 18468 11396 18524
rect 11396 18468 11452 18524
rect 11452 18468 11456 18524
rect 11392 18464 11456 18468
rect 11472 18524 11536 18528
rect 11472 18468 11476 18524
rect 11476 18468 11532 18524
rect 11532 18468 11536 18524
rect 11472 18464 11536 18468
rect 14659 18524 14723 18528
rect 14659 18468 14663 18524
rect 14663 18468 14719 18524
rect 14719 18468 14723 18524
rect 14659 18464 14723 18468
rect 14739 18524 14803 18528
rect 14739 18468 14743 18524
rect 14743 18468 14799 18524
rect 14799 18468 14803 18524
rect 14739 18464 14803 18468
rect 14819 18524 14883 18528
rect 14819 18468 14823 18524
rect 14823 18468 14879 18524
rect 14879 18468 14883 18524
rect 14819 18464 14883 18468
rect 14899 18524 14963 18528
rect 14899 18468 14903 18524
rect 14903 18468 14959 18524
rect 14959 18468 14963 18524
rect 14899 18464 14963 18468
rect 10364 18124 10428 18188
rect 13492 18124 13556 18188
rect 2665 17980 2729 17984
rect 2665 17924 2669 17980
rect 2669 17924 2725 17980
rect 2725 17924 2729 17980
rect 2665 17920 2729 17924
rect 2745 17980 2809 17984
rect 2745 17924 2749 17980
rect 2749 17924 2805 17980
rect 2805 17924 2809 17980
rect 2745 17920 2809 17924
rect 2825 17980 2889 17984
rect 2825 17924 2829 17980
rect 2829 17924 2885 17980
rect 2885 17924 2889 17980
rect 2825 17920 2889 17924
rect 2905 17980 2969 17984
rect 2905 17924 2909 17980
rect 2909 17924 2965 17980
rect 2965 17924 2969 17980
rect 2905 17920 2969 17924
rect 6092 17980 6156 17984
rect 6092 17924 6096 17980
rect 6096 17924 6152 17980
rect 6152 17924 6156 17980
rect 6092 17920 6156 17924
rect 6172 17980 6236 17984
rect 6172 17924 6176 17980
rect 6176 17924 6232 17980
rect 6232 17924 6236 17980
rect 6172 17920 6236 17924
rect 6252 17980 6316 17984
rect 6252 17924 6256 17980
rect 6256 17924 6312 17980
rect 6312 17924 6316 17980
rect 6252 17920 6316 17924
rect 6332 17980 6396 17984
rect 6332 17924 6336 17980
rect 6336 17924 6392 17980
rect 6392 17924 6396 17980
rect 6332 17920 6396 17924
rect 9519 17980 9583 17984
rect 9519 17924 9523 17980
rect 9523 17924 9579 17980
rect 9579 17924 9583 17980
rect 9519 17920 9583 17924
rect 9599 17980 9663 17984
rect 9599 17924 9603 17980
rect 9603 17924 9659 17980
rect 9659 17924 9663 17980
rect 9599 17920 9663 17924
rect 9679 17980 9743 17984
rect 9679 17924 9683 17980
rect 9683 17924 9739 17980
rect 9739 17924 9743 17980
rect 9679 17920 9743 17924
rect 9759 17980 9823 17984
rect 9759 17924 9763 17980
rect 9763 17924 9819 17980
rect 9819 17924 9823 17980
rect 9759 17920 9823 17924
rect 12946 17980 13010 17984
rect 12946 17924 12950 17980
rect 12950 17924 13006 17980
rect 13006 17924 13010 17980
rect 12946 17920 13010 17924
rect 13026 17980 13090 17984
rect 13026 17924 13030 17980
rect 13030 17924 13086 17980
rect 13086 17924 13090 17980
rect 13026 17920 13090 17924
rect 13106 17980 13170 17984
rect 13106 17924 13110 17980
rect 13110 17924 13166 17980
rect 13166 17924 13170 17980
rect 13106 17920 13170 17924
rect 13186 17980 13250 17984
rect 13186 17924 13190 17980
rect 13190 17924 13246 17980
rect 13246 17924 13250 17980
rect 13186 17920 13250 17924
rect 11836 17852 11900 17916
rect 4378 17436 4442 17440
rect 4378 17380 4382 17436
rect 4382 17380 4438 17436
rect 4438 17380 4442 17436
rect 4378 17376 4442 17380
rect 4458 17436 4522 17440
rect 4458 17380 4462 17436
rect 4462 17380 4518 17436
rect 4518 17380 4522 17436
rect 4458 17376 4522 17380
rect 4538 17436 4602 17440
rect 4538 17380 4542 17436
rect 4542 17380 4598 17436
rect 4598 17380 4602 17436
rect 4538 17376 4602 17380
rect 4618 17436 4682 17440
rect 4618 17380 4622 17436
rect 4622 17380 4678 17436
rect 4678 17380 4682 17436
rect 4618 17376 4682 17380
rect 7805 17436 7869 17440
rect 7805 17380 7809 17436
rect 7809 17380 7865 17436
rect 7865 17380 7869 17436
rect 7805 17376 7869 17380
rect 7885 17436 7949 17440
rect 7885 17380 7889 17436
rect 7889 17380 7945 17436
rect 7945 17380 7949 17436
rect 7885 17376 7949 17380
rect 7965 17436 8029 17440
rect 7965 17380 7969 17436
rect 7969 17380 8025 17436
rect 8025 17380 8029 17436
rect 7965 17376 8029 17380
rect 8045 17436 8109 17440
rect 8045 17380 8049 17436
rect 8049 17380 8105 17436
rect 8105 17380 8109 17436
rect 8045 17376 8109 17380
rect 11232 17436 11296 17440
rect 11232 17380 11236 17436
rect 11236 17380 11292 17436
rect 11292 17380 11296 17436
rect 11232 17376 11296 17380
rect 11312 17436 11376 17440
rect 11312 17380 11316 17436
rect 11316 17380 11372 17436
rect 11372 17380 11376 17436
rect 11312 17376 11376 17380
rect 11392 17436 11456 17440
rect 11392 17380 11396 17436
rect 11396 17380 11452 17436
rect 11452 17380 11456 17436
rect 11392 17376 11456 17380
rect 11472 17436 11536 17440
rect 11472 17380 11476 17436
rect 11476 17380 11532 17436
rect 11532 17380 11536 17436
rect 11472 17376 11536 17380
rect 14659 17436 14723 17440
rect 14659 17380 14663 17436
rect 14663 17380 14719 17436
rect 14719 17380 14723 17436
rect 14659 17376 14723 17380
rect 14739 17436 14803 17440
rect 14739 17380 14743 17436
rect 14743 17380 14799 17436
rect 14799 17380 14803 17436
rect 14739 17376 14803 17380
rect 14819 17436 14883 17440
rect 14819 17380 14823 17436
rect 14823 17380 14879 17436
rect 14879 17380 14883 17436
rect 14819 17376 14883 17380
rect 14899 17436 14963 17440
rect 14899 17380 14903 17436
rect 14903 17380 14959 17436
rect 14959 17380 14963 17436
rect 14899 17376 14963 17380
rect 13860 17172 13924 17236
rect 2665 16892 2729 16896
rect 2665 16836 2669 16892
rect 2669 16836 2725 16892
rect 2725 16836 2729 16892
rect 2665 16832 2729 16836
rect 2745 16892 2809 16896
rect 2745 16836 2749 16892
rect 2749 16836 2805 16892
rect 2805 16836 2809 16892
rect 2745 16832 2809 16836
rect 2825 16892 2889 16896
rect 2825 16836 2829 16892
rect 2829 16836 2885 16892
rect 2885 16836 2889 16892
rect 2825 16832 2889 16836
rect 2905 16892 2969 16896
rect 2905 16836 2909 16892
rect 2909 16836 2965 16892
rect 2965 16836 2969 16892
rect 2905 16832 2969 16836
rect 6092 16892 6156 16896
rect 6092 16836 6096 16892
rect 6096 16836 6152 16892
rect 6152 16836 6156 16892
rect 6092 16832 6156 16836
rect 6172 16892 6236 16896
rect 6172 16836 6176 16892
rect 6176 16836 6232 16892
rect 6232 16836 6236 16892
rect 6172 16832 6236 16836
rect 6252 16892 6316 16896
rect 6252 16836 6256 16892
rect 6256 16836 6312 16892
rect 6312 16836 6316 16892
rect 6252 16832 6316 16836
rect 6332 16892 6396 16896
rect 6332 16836 6336 16892
rect 6336 16836 6392 16892
rect 6392 16836 6396 16892
rect 6332 16832 6396 16836
rect 9519 16892 9583 16896
rect 9519 16836 9523 16892
rect 9523 16836 9579 16892
rect 9579 16836 9583 16892
rect 9519 16832 9583 16836
rect 9599 16892 9663 16896
rect 9599 16836 9603 16892
rect 9603 16836 9659 16892
rect 9659 16836 9663 16892
rect 9599 16832 9663 16836
rect 9679 16892 9743 16896
rect 9679 16836 9683 16892
rect 9683 16836 9739 16892
rect 9739 16836 9743 16892
rect 9679 16832 9743 16836
rect 9759 16892 9823 16896
rect 9759 16836 9763 16892
rect 9763 16836 9819 16892
rect 9819 16836 9823 16892
rect 9759 16832 9823 16836
rect 12946 16892 13010 16896
rect 12946 16836 12950 16892
rect 12950 16836 13006 16892
rect 13006 16836 13010 16892
rect 12946 16832 13010 16836
rect 13026 16892 13090 16896
rect 13026 16836 13030 16892
rect 13030 16836 13086 16892
rect 13086 16836 13090 16892
rect 13026 16832 13090 16836
rect 13106 16892 13170 16896
rect 13106 16836 13110 16892
rect 13110 16836 13166 16892
rect 13166 16836 13170 16892
rect 13106 16832 13170 16836
rect 13186 16892 13250 16896
rect 13186 16836 13190 16892
rect 13190 16836 13246 16892
rect 13246 16836 13250 16892
rect 13186 16832 13250 16836
rect 10548 16492 10612 16556
rect 4378 16348 4442 16352
rect 4378 16292 4382 16348
rect 4382 16292 4438 16348
rect 4438 16292 4442 16348
rect 4378 16288 4442 16292
rect 4458 16348 4522 16352
rect 4458 16292 4462 16348
rect 4462 16292 4518 16348
rect 4518 16292 4522 16348
rect 4458 16288 4522 16292
rect 4538 16348 4602 16352
rect 4538 16292 4542 16348
rect 4542 16292 4598 16348
rect 4598 16292 4602 16348
rect 4538 16288 4602 16292
rect 4618 16348 4682 16352
rect 4618 16292 4622 16348
rect 4622 16292 4678 16348
rect 4678 16292 4682 16348
rect 4618 16288 4682 16292
rect 7805 16348 7869 16352
rect 7805 16292 7809 16348
rect 7809 16292 7865 16348
rect 7865 16292 7869 16348
rect 7805 16288 7869 16292
rect 7885 16348 7949 16352
rect 7885 16292 7889 16348
rect 7889 16292 7945 16348
rect 7945 16292 7949 16348
rect 7885 16288 7949 16292
rect 7965 16348 8029 16352
rect 7965 16292 7969 16348
rect 7969 16292 8025 16348
rect 8025 16292 8029 16348
rect 7965 16288 8029 16292
rect 8045 16348 8109 16352
rect 8045 16292 8049 16348
rect 8049 16292 8105 16348
rect 8105 16292 8109 16348
rect 8045 16288 8109 16292
rect 11232 16348 11296 16352
rect 11232 16292 11236 16348
rect 11236 16292 11292 16348
rect 11292 16292 11296 16348
rect 11232 16288 11296 16292
rect 11312 16348 11376 16352
rect 11312 16292 11316 16348
rect 11316 16292 11372 16348
rect 11372 16292 11376 16348
rect 11312 16288 11376 16292
rect 11392 16348 11456 16352
rect 11392 16292 11396 16348
rect 11396 16292 11452 16348
rect 11452 16292 11456 16348
rect 11392 16288 11456 16292
rect 11472 16348 11536 16352
rect 11472 16292 11476 16348
rect 11476 16292 11532 16348
rect 11532 16292 11536 16348
rect 11472 16288 11536 16292
rect 14659 16348 14723 16352
rect 14659 16292 14663 16348
rect 14663 16292 14719 16348
rect 14719 16292 14723 16348
rect 14659 16288 14723 16292
rect 14739 16348 14803 16352
rect 14739 16292 14743 16348
rect 14743 16292 14799 16348
rect 14799 16292 14803 16348
rect 14739 16288 14803 16292
rect 14819 16348 14883 16352
rect 14819 16292 14823 16348
rect 14823 16292 14879 16348
rect 14879 16292 14883 16348
rect 14819 16288 14883 16292
rect 14899 16348 14963 16352
rect 14899 16292 14903 16348
rect 14903 16292 14959 16348
rect 14959 16292 14963 16348
rect 14899 16288 14963 16292
rect 13492 16220 13556 16284
rect 13860 16280 13924 16284
rect 13860 16224 13874 16280
rect 13874 16224 13924 16280
rect 13860 16220 13924 16224
rect 8892 16084 8956 16148
rect 12756 16144 12820 16148
rect 12756 16088 12770 16144
rect 12770 16088 12820 16144
rect 12756 16084 12820 16088
rect 12572 15812 12636 15876
rect 2665 15804 2729 15808
rect 2665 15748 2669 15804
rect 2669 15748 2725 15804
rect 2725 15748 2729 15804
rect 2665 15744 2729 15748
rect 2745 15804 2809 15808
rect 2745 15748 2749 15804
rect 2749 15748 2805 15804
rect 2805 15748 2809 15804
rect 2745 15744 2809 15748
rect 2825 15804 2889 15808
rect 2825 15748 2829 15804
rect 2829 15748 2885 15804
rect 2885 15748 2889 15804
rect 2825 15744 2889 15748
rect 2905 15804 2969 15808
rect 2905 15748 2909 15804
rect 2909 15748 2965 15804
rect 2965 15748 2969 15804
rect 2905 15744 2969 15748
rect 6092 15804 6156 15808
rect 6092 15748 6096 15804
rect 6096 15748 6152 15804
rect 6152 15748 6156 15804
rect 6092 15744 6156 15748
rect 6172 15804 6236 15808
rect 6172 15748 6176 15804
rect 6176 15748 6232 15804
rect 6232 15748 6236 15804
rect 6172 15744 6236 15748
rect 6252 15804 6316 15808
rect 6252 15748 6256 15804
rect 6256 15748 6312 15804
rect 6312 15748 6316 15804
rect 6252 15744 6316 15748
rect 6332 15804 6396 15808
rect 6332 15748 6336 15804
rect 6336 15748 6392 15804
rect 6392 15748 6396 15804
rect 6332 15744 6396 15748
rect 9519 15804 9583 15808
rect 9519 15748 9523 15804
rect 9523 15748 9579 15804
rect 9579 15748 9583 15804
rect 9519 15744 9583 15748
rect 9599 15804 9663 15808
rect 9599 15748 9603 15804
rect 9603 15748 9659 15804
rect 9659 15748 9663 15804
rect 9599 15744 9663 15748
rect 9679 15804 9743 15808
rect 9679 15748 9683 15804
rect 9683 15748 9739 15804
rect 9739 15748 9743 15804
rect 9679 15744 9743 15748
rect 9759 15804 9823 15808
rect 9759 15748 9763 15804
rect 9763 15748 9819 15804
rect 9819 15748 9823 15804
rect 9759 15744 9823 15748
rect 12946 15804 13010 15808
rect 12946 15748 12950 15804
rect 12950 15748 13006 15804
rect 13006 15748 13010 15804
rect 12946 15744 13010 15748
rect 13026 15804 13090 15808
rect 13026 15748 13030 15804
rect 13030 15748 13086 15804
rect 13086 15748 13090 15804
rect 13026 15744 13090 15748
rect 13106 15804 13170 15808
rect 13106 15748 13110 15804
rect 13110 15748 13166 15804
rect 13166 15748 13170 15804
rect 13106 15744 13170 15748
rect 13186 15804 13250 15808
rect 13186 15748 13190 15804
rect 13190 15748 13246 15804
rect 13246 15748 13250 15804
rect 13186 15744 13250 15748
rect 11652 15540 11716 15604
rect 4378 15260 4442 15264
rect 4378 15204 4382 15260
rect 4382 15204 4438 15260
rect 4438 15204 4442 15260
rect 4378 15200 4442 15204
rect 4458 15260 4522 15264
rect 4458 15204 4462 15260
rect 4462 15204 4518 15260
rect 4518 15204 4522 15260
rect 4458 15200 4522 15204
rect 4538 15260 4602 15264
rect 4538 15204 4542 15260
rect 4542 15204 4598 15260
rect 4598 15204 4602 15260
rect 4538 15200 4602 15204
rect 4618 15260 4682 15264
rect 4618 15204 4622 15260
rect 4622 15204 4678 15260
rect 4678 15204 4682 15260
rect 4618 15200 4682 15204
rect 7805 15260 7869 15264
rect 7805 15204 7809 15260
rect 7809 15204 7865 15260
rect 7865 15204 7869 15260
rect 7805 15200 7869 15204
rect 7885 15260 7949 15264
rect 7885 15204 7889 15260
rect 7889 15204 7945 15260
rect 7945 15204 7949 15260
rect 7885 15200 7949 15204
rect 7965 15260 8029 15264
rect 7965 15204 7969 15260
rect 7969 15204 8025 15260
rect 8025 15204 8029 15260
rect 7965 15200 8029 15204
rect 8045 15260 8109 15264
rect 8045 15204 8049 15260
rect 8049 15204 8105 15260
rect 8105 15204 8109 15260
rect 8045 15200 8109 15204
rect 11232 15260 11296 15264
rect 11232 15204 11236 15260
rect 11236 15204 11292 15260
rect 11292 15204 11296 15260
rect 11232 15200 11296 15204
rect 11312 15260 11376 15264
rect 11312 15204 11316 15260
rect 11316 15204 11372 15260
rect 11372 15204 11376 15260
rect 11312 15200 11376 15204
rect 11392 15260 11456 15264
rect 11392 15204 11396 15260
rect 11396 15204 11452 15260
rect 11452 15204 11456 15260
rect 11392 15200 11456 15204
rect 11472 15260 11536 15264
rect 11472 15204 11476 15260
rect 11476 15204 11532 15260
rect 11532 15204 11536 15260
rect 11472 15200 11536 15204
rect 14659 15260 14723 15264
rect 14659 15204 14663 15260
rect 14663 15204 14719 15260
rect 14719 15204 14723 15260
rect 14659 15200 14723 15204
rect 14739 15260 14803 15264
rect 14739 15204 14743 15260
rect 14743 15204 14799 15260
rect 14799 15204 14803 15260
rect 14739 15200 14803 15204
rect 14819 15260 14883 15264
rect 14819 15204 14823 15260
rect 14823 15204 14879 15260
rect 14879 15204 14883 15260
rect 14819 15200 14883 15204
rect 14899 15260 14963 15264
rect 14899 15204 14903 15260
rect 14903 15204 14959 15260
rect 14959 15204 14963 15260
rect 14899 15200 14963 15204
rect 2665 14716 2729 14720
rect 2665 14660 2669 14716
rect 2669 14660 2725 14716
rect 2725 14660 2729 14716
rect 2665 14656 2729 14660
rect 2745 14716 2809 14720
rect 2745 14660 2749 14716
rect 2749 14660 2805 14716
rect 2805 14660 2809 14716
rect 2745 14656 2809 14660
rect 2825 14716 2889 14720
rect 2825 14660 2829 14716
rect 2829 14660 2885 14716
rect 2885 14660 2889 14716
rect 2825 14656 2889 14660
rect 2905 14716 2969 14720
rect 2905 14660 2909 14716
rect 2909 14660 2965 14716
rect 2965 14660 2969 14716
rect 2905 14656 2969 14660
rect 6092 14716 6156 14720
rect 6092 14660 6096 14716
rect 6096 14660 6152 14716
rect 6152 14660 6156 14716
rect 6092 14656 6156 14660
rect 6172 14716 6236 14720
rect 6172 14660 6176 14716
rect 6176 14660 6232 14716
rect 6232 14660 6236 14716
rect 6172 14656 6236 14660
rect 6252 14716 6316 14720
rect 6252 14660 6256 14716
rect 6256 14660 6312 14716
rect 6312 14660 6316 14716
rect 6252 14656 6316 14660
rect 6332 14716 6396 14720
rect 6332 14660 6336 14716
rect 6336 14660 6392 14716
rect 6392 14660 6396 14716
rect 6332 14656 6396 14660
rect 9519 14716 9583 14720
rect 9519 14660 9523 14716
rect 9523 14660 9579 14716
rect 9579 14660 9583 14716
rect 9519 14656 9583 14660
rect 9599 14716 9663 14720
rect 9599 14660 9603 14716
rect 9603 14660 9659 14716
rect 9659 14660 9663 14716
rect 9599 14656 9663 14660
rect 9679 14716 9743 14720
rect 9679 14660 9683 14716
rect 9683 14660 9739 14716
rect 9739 14660 9743 14716
rect 9679 14656 9743 14660
rect 9759 14716 9823 14720
rect 9759 14660 9763 14716
rect 9763 14660 9819 14716
rect 9819 14660 9823 14716
rect 9759 14656 9823 14660
rect 12946 14716 13010 14720
rect 12946 14660 12950 14716
rect 12950 14660 13006 14716
rect 13006 14660 13010 14716
rect 12946 14656 13010 14660
rect 13026 14716 13090 14720
rect 13026 14660 13030 14716
rect 13030 14660 13086 14716
rect 13086 14660 13090 14716
rect 13026 14656 13090 14660
rect 13106 14716 13170 14720
rect 13106 14660 13110 14716
rect 13110 14660 13166 14716
rect 13166 14660 13170 14716
rect 13106 14656 13170 14660
rect 13186 14716 13250 14720
rect 13186 14660 13190 14716
rect 13190 14660 13246 14716
rect 13246 14660 13250 14716
rect 13186 14656 13250 14660
rect 10364 14452 10428 14516
rect 4378 14172 4442 14176
rect 4378 14116 4382 14172
rect 4382 14116 4438 14172
rect 4438 14116 4442 14172
rect 4378 14112 4442 14116
rect 4458 14172 4522 14176
rect 4458 14116 4462 14172
rect 4462 14116 4518 14172
rect 4518 14116 4522 14172
rect 4458 14112 4522 14116
rect 4538 14172 4602 14176
rect 4538 14116 4542 14172
rect 4542 14116 4598 14172
rect 4598 14116 4602 14172
rect 4538 14112 4602 14116
rect 4618 14172 4682 14176
rect 4618 14116 4622 14172
rect 4622 14116 4678 14172
rect 4678 14116 4682 14172
rect 4618 14112 4682 14116
rect 7805 14172 7869 14176
rect 7805 14116 7809 14172
rect 7809 14116 7865 14172
rect 7865 14116 7869 14172
rect 7805 14112 7869 14116
rect 7885 14172 7949 14176
rect 7885 14116 7889 14172
rect 7889 14116 7945 14172
rect 7945 14116 7949 14172
rect 7885 14112 7949 14116
rect 7965 14172 8029 14176
rect 7965 14116 7969 14172
rect 7969 14116 8025 14172
rect 8025 14116 8029 14172
rect 7965 14112 8029 14116
rect 8045 14172 8109 14176
rect 8045 14116 8049 14172
rect 8049 14116 8105 14172
rect 8105 14116 8109 14172
rect 8045 14112 8109 14116
rect 11232 14172 11296 14176
rect 11232 14116 11236 14172
rect 11236 14116 11292 14172
rect 11292 14116 11296 14172
rect 11232 14112 11296 14116
rect 11312 14172 11376 14176
rect 11312 14116 11316 14172
rect 11316 14116 11372 14172
rect 11372 14116 11376 14172
rect 11312 14112 11376 14116
rect 11392 14172 11456 14176
rect 11392 14116 11396 14172
rect 11396 14116 11452 14172
rect 11452 14116 11456 14172
rect 11392 14112 11456 14116
rect 11472 14172 11536 14176
rect 11472 14116 11476 14172
rect 11476 14116 11532 14172
rect 11532 14116 11536 14172
rect 11472 14112 11536 14116
rect 14659 14172 14723 14176
rect 14659 14116 14663 14172
rect 14663 14116 14719 14172
rect 14719 14116 14723 14172
rect 14659 14112 14723 14116
rect 14739 14172 14803 14176
rect 14739 14116 14743 14172
rect 14743 14116 14799 14172
rect 14799 14116 14803 14172
rect 14739 14112 14803 14116
rect 14819 14172 14883 14176
rect 14819 14116 14823 14172
rect 14823 14116 14879 14172
rect 14879 14116 14883 14172
rect 14819 14112 14883 14116
rect 14899 14172 14963 14176
rect 14899 14116 14903 14172
rect 14903 14116 14959 14172
rect 14959 14116 14963 14172
rect 14899 14112 14963 14116
rect 1716 14104 1780 14108
rect 1716 14048 1730 14104
rect 1730 14048 1780 14104
rect 1716 14044 1780 14048
rect 13676 13832 13740 13836
rect 13676 13776 13726 13832
rect 13726 13776 13740 13832
rect 13676 13772 13740 13776
rect 2665 13628 2729 13632
rect 2665 13572 2669 13628
rect 2669 13572 2725 13628
rect 2725 13572 2729 13628
rect 2665 13568 2729 13572
rect 2745 13628 2809 13632
rect 2745 13572 2749 13628
rect 2749 13572 2805 13628
rect 2805 13572 2809 13628
rect 2745 13568 2809 13572
rect 2825 13628 2889 13632
rect 2825 13572 2829 13628
rect 2829 13572 2885 13628
rect 2885 13572 2889 13628
rect 2825 13568 2889 13572
rect 2905 13628 2969 13632
rect 2905 13572 2909 13628
rect 2909 13572 2965 13628
rect 2965 13572 2969 13628
rect 2905 13568 2969 13572
rect 6092 13628 6156 13632
rect 6092 13572 6096 13628
rect 6096 13572 6152 13628
rect 6152 13572 6156 13628
rect 6092 13568 6156 13572
rect 6172 13628 6236 13632
rect 6172 13572 6176 13628
rect 6176 13572 6232 13628
rect 6232 13572 6236 13628
rect 6172 13568 6236 13572
rect 6252 13628 6316 13632
rect 6252 13572 6256 13628
rect 6256 13572 6312 13628
rect 6312 13572 6316 13628
rect 6252 13568 6316 13572
rect 6332 13628 6396 13632
rect 6332 13572 6336 13628
rect 6336 13572 6392 13628
rect 6392 13572 6396 13628
rect 6332 13568 6396 13572
rect 9519 13628 9583 13632
rect 9519 13572 9523 13628
rect 9523 13572 9579 13628
rect 9579 13572 9583 13628
rect 9519 13568 9583 13572
rect 9599 13628 9663 13632
rect 9599 13572 9603 13628
rect 9603 13572 9659 13628
rect 9659 13572 9663 13628
rect 9599 13568 9663 13572
rect 9679 13628 9743 13632
rect 9679 13572 9683 13628
rect 9683 13572 9739 13628
rect 9739 13572 9743 13628
rect 9679 13568 9743 13572
rect 9759 13628 9823 13632
rect 9759 13572 9763 13628
rect 9763 13572 9819 13628
rect 9819 13572 9823 13628
rect 9759 13568 9823 13572
rect 12946 13628 13010 13632
rect 12946 13572 12950 13628
rect 12950 13572 13006 13628
rect 13006 13572 13010 13628
rect 12946 13568 13010 13572
rect 13026 13628 13090 13632
rect 13026 13572 13030 13628
rect 13030 13572 13086 13628
rect 13086 13572 13090 13628
rect 13026 13568 13090 13572
rect 13106 13628 13170 13632
rect 13106 13572 13110 13628
rect 13110 13572 13166 13628
rect 13166 13572 13170 13628
rect 13106 13568 13170 13572
rect 13186 13628 13250 13632
rect 13186 13572 13190 13628
rect 13190 13572 13246 13628
rect 13246 13572 13250 13628
rect 13186 13568 13250 13572
rect 10732 13500 10796 13564
rect 11836 13500 11900 13564
rect 4378 13084 4442 13088
rect 4378 13028 4382 13084
rect 4382 13028 4438 13084
rect 4438 13028 4442 13084
rect 4378 13024 4442 13028
rect 4458 13084 4522 13088
rect 4458 13028 4462 13084
rect 4462 13028 4518 13084
rect 4518 13028 4522 13084
rect 4458 13024 4522 13028
rect 4538 13084 4602 13088
rect 4538 13028 4542 13084
rect 4542 13028 4598 13084
rect 4598 13028 4602 13084
rect 4538 13024 4602 13028
rect 4618 13084 4682 13088
rect 4618 13028 4622 13084
rect 4622 13028 4678 13084
rect 4678 13028 4682 13084
rect 4618 13024 4682 13028
rect 7805 13084 7869 13088
rect 7805 13028 7809 13084
rect 7809 13028 7865 13084
rect 7865 13028 7869 13084
rect 7805 13024 7869 13028
rect 7885 13084 7949 13088
rect 7885 13028 7889 13084
rect 7889 13028 7945 13084
rect 7945 13028 7949 13084
rect 7885 13024 7949 13028
rect 7965 13084 8029 13088
rect 7965 13028 7969 13084
rect 7969 13028 8025 13084
rect 8025 13028 8029 13084
rect 7965 13024 8029 13028
rect 8045 13084 8109 13088
rect 8045 13028 8049 13084
rect 8049 13028 8105 13084
rect 8105 13028 8109 13084
rect 8045 13024 8109 13028
rect 3924 12820 3988 12884
rect 15332 13500 15396 13564
rect 11232 13084 11296 13088
rect 11232 13028 11236 13084
rect 11236 13028 11292 13084
rect 11292 13028 11296 13084
rect 11232 13024 11296 13028
rect 11312 13084 11376 13088
rect 11312 13028 11316 13084
rect 11316 13028 11372 13084
rect 11372 13028 11376 13084
rect 11312 13024 11376 13028
rect 11392 13084 11456 13088
rect 11392 13028 11396 13084
rect 11396 13028 11452 13084
rect 11452 13028 11456 13084
rect 11392 13024 11456 13028
rect 11472 13084 11536 13088
rect 11472 13028 11476 13084
rect 11476 13028 11532 13084
rect 11532 13028 11536 13084
rect 11472 13024 11536 13028
rect 14659 13084 14723 13088
rect 14659 13028 14663 13084
rect 14663 13028 14719 13084
rect 14719 13028 14723 13084
rect 14659 13024 14723 13028
rect 14739 13084 14803 13088
rect 14739 13028 14743 13084
rect 14743 13028 14799 13084
rect 14799 13028 14803 13084
rect 14739 13024 14803 13028
rect 14819 13084 14883 13088
rect 14819 13028 14823 13084
rect 14823 13028 14879 13084
rect 14879 13028 14883 13084
rect 14819 13024 14883 13028
rect 14899 13084 14963 13088
rect 14899 13028 14903 13084
rect 14903 13028 14959 13084
rect 14959 13028 14963 13084
rect 14899 13024 14963 13028
rect 12572 12548 12636 12612
rect 2665 12540 2729 12544
rect 2665 12484 2669 12540
rect 2669 12484 2725 12540
rect 2725 12484 2729 12540
rect 2665 12480 2729 12484
rect 2745 12540 2809 12544
rect 2745 12484 2749 12540
rect 2749 12484 2805 12540
rect 2805 12484 2809 12540
rect 2745 12480 2809 12484
rect 2825 12540 2889 12544
rect 2825 12484 2829 12540
rect 2829 12484 2885 12540
rect 2885 12484 2889 12540
rect 2825 12480 2889 12484
rect 2905 12540 2969 12544
rect 2905 12484 2909 12540
rect 2909 12484 2965 12540
rect 2965 12484 2969 12540
rect 2905 12480 2969 12484
rect 6092 12540 6156 12544
rect 6092 12484 6096 12540
rect 6096 12484 6152 12540
rect 6152 12484 6156 12540
rect 6092 12480 6156 12484
rect 6172 12540 6236 12544
rect 6172 12484 6176 12540
rect 6176 12484 6232 12540
rect 6232 12484 6236 12540
rect 6172 12480 6236 12484
rect 6252 12540 6316 12544
rect 6252 12484 6256 12540
rect 6256 12484 6312 12540
rect 6312 12484 6316 12540
rect 6252 12480 6316 12484
rect 6332 12540 6396 12544
rect 6332 12484 6336 12540
rect 6336 12484 6392 12540
rect 6392 12484 6396 12540
rect 6332 12480 6396 12484
rect 9519 12540 9583 12544
rect 9519 12484 9523 12540
rect 9523 12484 9579 12540
rect 9579 12484 9583 12540
rect 9519 12480 9583 12484
rect 9599 12540 9663 12544
rect 9599 12484 9603 12540
rect 9603 12484 9659 12540
rect 9659 12484 9663 12540
rect 9599 12480 9663 12484
rect 9679 12540 9743 12544
rect 9679 12484 9683 12540
rect 9683 12484 9739 12540
rect 9739 12484 9743 12540
rect 9679 12480 9743 12484
rect 9759 12540 9823 12544
rect 9759 12484 9763 12540
rect 9763 12484 9819 12540
rect 9819 12484 9823 12540
rect 9759 12480 9823 12484
rect 12946 12540 13010 12544
rect 12946 12484 12950 12540
rect 12950 12484 13006 12540
rect 13006 12484 13010 12540
rect 12946 12480 13010 12484
rect 13026 12540 13090 12544
rect 13026 12484 13030 12540
rect 13030 12484 13086 12540
rect 13086 12484 13090 12540
rect 13026 12480 13090 12484
rect 13106 12540 13170 12544
rect 13106 12484 13110 12540
rect 13110 12484 13166 12540
rect 13166 12484 13170 12540
rect 13106 12480 13170 12484
rect 13186 12540 13250 12544
rect 13186 12484 13190 12540
rect 13190 12484 13246 12540
rect 13246 12484 13250 12540
rect 13186 12480 13250 12484
rect 12756 12412 12820 12476
rect 13860 12412 13924 12476
rect 11652 12336 11716 12340
rect 11652 12280 11666 12336
rect 11666 12280 11716 12336
rect 11652 12276 11716 12280
rect 4378 11996 4442 12000
rect 4378 11940 4382 11996
rect 4382 11940 4438 11996
rect 4438 11940 4442 11996
rect 4378 11936 4442 11940
rect 4458 11996 4522 12000
rect 4458 11940 4462 11996
rect 4462 11940 4518 11996
rect 4518 11940 4522 11996
rect 4458 11936 4522 11940
rect 4538 11996 4602 12000
rect 4538 11940 4542 11996
rect 4542 11940 4598 11996
rect 4598 11940 4602 11996
rect 4538 11936 4602 11940
rect 4618 11996 4682 12000
rect 4618 11940 4622 11996
rect 4622 11940 4678 11996
rect 4678 11940 4682 11996
rect 4618 11936 4682 11940
rect 7805 11996 7869 12000
rect 7805 11940 7809 11996
rect 7809 11940 7865 11996
rect 7865 11940 7869 11996
rect 7805 11936 7869 11940
rect 7885 11996 7949 12000
rect 7885 11940 7889 11996
rect 7889 11940 7945 11996
rect 7945 11940 7949 11996
rect 7885 11936 7949 11940
rect 7965 11996 8029 12000
rect 7965 11940 7969 11996
rect 7969 11940 8025 11996
rect 8025 11940 8029 11996
rect 7965 11936 8029 11940
rect 8045 11996 8109 12000
rect 8045 11940 8049 11996
rect 8049 11940 8105 11996
rect 8105 11940 8109 11996
rect 8045 11936 8109 11940
rect 11232 11996 11296 12000
rect 11232 11940 11236 11996
rect 11236 11940 11292 11996
rect 11292 11940 11296 11996
rect 11232 11936 11296 11940
rect 11312 11996 11376 12000
rect 11312 11940 11316 11996
rect 11316 11940 11372 11996
rect 11372 11940 11376 11996
rect 11312 11936 11376 11940
rect 11392 11996 11456 12000
rect 11392 11940 11396 11996
rect 11396 11940 11452 11996
rect 11452 11940 11456 11996
rect 11392 11936 11456 11940
rect 11472 11996 11536 12000
rect 11472 11940 11476 11996
rect 11476 11940 11532 11996
rect 11532 11940 11536 11996
rect 11472 11936 11536 11940
rect 14659 11996 14723 12000
rect 14659 11940 14663 11996
rect 14663 11940 14719 11996
rect 14719 11940 14723 11996
rect 14659 11936 14723 11940
rect 14739 11996 14803 12000
rect 14739 11940 14743 11996
rect 14743 11940 14799 11996
rect 14799 11940 14803 11996
rect 14739 11936 14803 11940
rect 14819 11996 14883 12000
rect 14819 11940 14823 11996
rect 14823 11940 14879 11996
rect 14879 11940 14883 11996
rect 14819 11936 14883 11940
rect 14899 11996 14963 12000
rect 14899 11940 14903 11996
rect 14903 11940 14959 11996
rect 14959 11940 14963 11996
rect 14899 11936 14963 11940
rect 7236 11732 7300 11796
rect 2665 11452 2729 11456
rect 2665 11396 2669 11452
rect 2669 11396 2725 11452
rect 2725 11396 2729 11452
rect 2665 11392 2729 11396
rect 2745 11452 2809 11456
rect 2745 11396 2749 11452
rect 2749 11396 2805 11452
rect 2805 11396 2809 11452
rect 2745 11392 2809 11396
rect 2825 11452 2889 11456
rect 2825 11396 2829 11452
rect 2829 11396 2885 11452
rect 2885 11396 2889 11452
rect 2825 11392 2889 11396
rect 2905 11452 2969 11456
rect 2905 11396 2909 11452
rect 2909 11396 2965 11452
rect 2965 11396 2969 11452
rect 2905 11392 2969 11396
rect 6092 11452 6156 11456
rect 6092 11396 6096 11452
rect 6096 11396 6152 11452
rect 6152 11396 6156 11452
rect 6092 11392 6156 11396
rect 6172 11452 6236 11456
rect 6172 11396 6176 11452
rect 6176 11396 6232 11452
rect 6232 11396 6236 11452
rect 6172 11392 6236 11396
rect 6252 11452 6316 11456
rect 6252 11396 6256 11452
rect 6256 11396 6312 11452
rect 6312 11396 6316 11452
rect 6252 11392 6316 11396
rect 6332 11452 6396 11456
rect 6332 11396 6336 11452
rect 6336 11396 6392 11452
rect 6392 11396 6396 11452
rect 6332 11392 6396 11396
rect 9519 11452 9583 11456
rect 9519 11396 9523 11452
rect 9523 11396 9579 11452
rect 9579 11396 9583 11452
rect 9519 11392 9583 11396
rect 9599 11452 9663 11456
rect 9599 11396 9603 11452
rect 9603 11396 9659 11452
rect 9659 11396 9663 11452
rect 9599 11392 9663 11396
rect 9679 11452 9743 11456
rect 9679 11396 9683 11452
rect 9683 11396 9739 11452
rect 9739 11396 9743 11452
rect 9679 11392 9743 11396
rect 9759 11452 9823 11456
rect 9759 11396 9763 11452
rect 9763 11396 9819 11452
rect 9819 11396 9823 11452
rect 9759 11392 9823 11396
rect 12946 11452 13010 11456
rect 12946 11396 12950 11452
rect 12950 11396 13006 11452
rect 13006 11396 13010 11452
rect 12946 11392 13010 11396
rect 13026 11452 13090 11456
rect 13026 11396 13030 11452
rect 13030 11396 13086 11452
rect 13086 11396 13090 11452
rect 13026 11392 13090 11396
rect 13106 11452 13170 11456
rect 13106 11396 13110 11452
rect 13110 11396 13166 11452
rect 13166 11396 13170 11452
rect 13106 11392 13170 11396
rect 13186 11452 13250 11456
rect 13186 11396 13190 11452
rect 13190 11396 13246 11452
rect 13246 11396 13250 11452
rect 13186 11392 13250 11396
rect 4378 10908 4442 10912
rect 4378 10852 4382 10908
rect 4382 10852 4438 10908
rect 4438 10852 4442 10908
rect 4378 10848 4442 10852
rect 4458 10908 4522 10912
rect 4458 10852 4462 10908
rect 4462 10852 4518 10908
rect 4518 10852 4522 10908
rect 4458 10848 4522 10852
rect 4538 10908 4602 10912
rect 4538 10852 4542 10908
rect 4542 10852 4598 10908
rect 4598 10852 4602 10908
rect 4538 10848 4602 10852
rect 4618 10908 4682 10912
rect 4618 10852 4622 10908
rect 4622 10852 4678 10908
rect 4678 10852 4682 10908
rect 4618 10848 4682 10852
rect 7805 10908 7869 10912
rect 7805 10852 7809 10908
rect 7809 10852 7865 10908
rect 7865 10852 7869 10908
rect 7805 10848 7869 10852
rect 7885 10908 7949 10912
rect 7885 10852 7889 10908
rect 7889 10852 7945 10908
rect 7945 10852 7949 10908
rect 7885 10848 7949 10852
rect 7965 10908 8029 10912
rect 7965 10852 7969 10908
rect 7969 10852 8025 10908
rect 8025 10852 8029 10908
rect 7965 10848 8029 10852
rect 8045 10908 8109 10912
rect 8045 10852 8049 10908
rect 8049 10852 8105 10908
rect 8105 10852 8109 10908
rect 8045 10848 8109 10852
rect 11232 10908 11296 10912
rect 11232 10852 11236 10908
rect 11236 10852 11292 10908
rect 11292 10852 11296 10908
rect 11232 10848 11296 10852
rect 11312 10908 11376 10912
rect 11312 10852 11316 10908
rect 11316 10852 11372 10908
rect 11372 10852 11376 10908
rect 11312 10848 11376 10852
rect 11392 10908 11456 10912
rect 11392 10852 11396 10908
rect 11396 10852 11452 10908
rect 11452 10852 11456 10908
rect 11392 10848 11456 10852
rect 11472 10908 11536 10912
rect 11472 10852 11476 10908
rect 11476 10852 11532 10908
rect 11532 10852 11536 10908
rect 11472 10848 11536 10852
rect 14659 10908 14723 10912
rect 14659 10852 14663 10908
rect 14663 10852 14719 10908
rect 14719 10852 14723 10908
rect 14659 10848 14723 10852
rect 14739 10908 14803 10912
rect 14739 10852 14743 10908
rect 14743 10852 14799 10908
rect 14799 10852 14803 10908
rect 14739 10848 14803 10852
rect 14819 10908 14883 10912
rect 14819 10852 14823 10908
rect 14823 10852 14879 10908
rect 14879 10852 14883 10908
rect 14819 10848 14883 10852
rect 14899 10908 14963 10912
rect 14899 10852 14903 10908
rect 14903 10852 14959 10908
rect 14959 10852 14963 10908
rect 14899 10848 14963 10852
rect 12204 10372 12268 10436
rect 2665 10364 2729 10368
rect 2665 10308 2669 10364
rect 2669 10308 2725 10364
rect 2725 10308 2729 10364
rect 2665 10304 2729 10308
rect 2745 10364 2809 10368
rect 2745 10308 2749 10364
rect 2749 10308 2805 10364
rect 2805 10308 2809 10364
rect 2745 10304 2809 10308
rect 2825 10364 2889 10368
rect 2825 10308 2829 10364
rect 2829 10308 2885 10364
rect 2885 10308 2889 10364
rect 2825 10304 2889 10308
rect 2905 10364 2969 10368
rect 2905 10308 2909 10364
rect 2909 10308 2965 10364
rect 2965 10308 2969 10364
rect 2905 10304 2969 10308
rect 6092 10364 6156 10368
rect 6092 10308 6096 10364
rect 6096 10308 6152 10364
rect 6152 10308 6156 10364
rect 6092 10304 6156 10308
rect 6172 10364 6236 10368
rect 6172 10308 6176 10364
rect 6176 10308 6232 10364
rect 6232 10308 6236 10364
rect 6172 10304 6236 10308
rect 6252 10364 6316 10368
rect 6252 10308 6256 10364
rect 6256 10308 6312 10364
rect 6312 10308 6316 10364
rect 6252 10304 6316 10308
rect 6332 10364 6396 10368
rect 6332 10308 6336 10364
rect 6336 10308 6392 10364
rect 6392 10308 6396 10364
rect 6332 10304 6396 10308
rect 9519 10364 9583 10368
rect 9519 10308 9523 10364
rect 9523 10308 9579 10364
rect 9579 10308 9583 10364
rect 9519 10304 9583 10308
rect 9599 10364 9663 10368
rect 9599 10308 9603 10364
rect 9603 10308 9659 10364
rect 9659 10308 9663 10364
rect 9599 10304 9663 10308
rect 9679 10364 9743 10368
rect 9679 10308 9683 10364
rect 9683 10308 9739 10364
rect 9739 10308 9743 10364
rect 9679 10304 9743 10308
rect 9759 10364 9823 10368
rect 9759 10308 9763 10364
rect 9763 10308 9819 10364
rect 9819 10308 9823 10364
rect 9759 10304 9823 10308
rect 12946 10364 13010 10368
rect 12946 10308 12950 10364
rect 12950 10308 13006 10364
rect 13006 10308 13010 10364
rect 12946 10304 13010 10308
rect 13026 10364 13090 10368
rect 13026 10308 13030 10364
rect 13030 10308 13086 10364
rect 13086 10308 13090 10364
rect 13026 10304 13090 10308
rect 13106 10364 13170 10368
rect 13106 10308 13110 10364
rect 13110 10308 13166 10364
rect 13166 10308 13170 10364
rect 13106 10304 13170 10308
rect 13186 10364 13250 10368
rect 13186 10308 13190 10364
rect 13190 10308 13246 10364
rect 13246 10308 13250 10364
rect 13186 10304 13250 10308
rect 10732 9828 10796 9892
rect 4378 9820 4442 9824
rect 4378 9764 4382 9820
rect 4382 9764 4438 9820
rect 4438 9764 4442 9820
rect 4378 9760 4442 9764
rect 4458 9820 4522 9824
rect 4458 9764 4462 9820
rect 4462 9764 4518 9820
rect 4518 9764 4522 9820
rect 4458 9760 4522 9764
rect 4538 9820 4602 9824
rect 4538 9764 4542 9820
rect 4542 9764 4598 9820
rect 4598 9764 4602 9820
rect 4538 9760 4602 9764
rect 4618 9820 4682 9824
rect 4618 9764 4622 9820
rect 4622 9764 4678 9820
rect 4678 9764 4682 9820
rect 4618 9760 4682 9764
rect 7805 9820 7869 9824
rect 7805 9764 7809 9820
rect 7809 9764 7865 9820
rect 7865 9764 7869 9820
rect 7805 9760 7869 9764
rect 7885 9820 7949 9824
rect 7885 9764 7889 9820
rect 7889 9764 7945 9820
rect 7945 9764 7949 9820
rect 7885 9760 7949 9764
rect 7965 9820 8029 9824
rect 7965 9764 7969 9820
rect 7969 9764 8025 9820
rect 8025 9764 8029 9820
rect 7965 9760 8029 9764
rect 8045 9820 8109 9824
rect 8045 9764 8049 9820
rect 8049 9764 8105 9820
rect 8105 9764 8109 9820
rect 8045 9760 8109 9764
rect 11232 9820 11296 9824
rect 11232 9764 11236 9820
rect 11236 9764 11292 9820
rect 11292 9764 11296 9820
rect 11232 9760 11296 9764
rect 11312 9820 11376 9824
rect 11312 9764 11316 9820
rect 11316 9764 11372 9820
rect 11372 9764 11376 9820
rect 11312 9760 11376 9764
rect 11392 9820 11456 9824
rect 11392 9764 11396 9820
rect 11396 9764 11452 9820
rect 11452 9764 11456 9820
rect 11392 9760 11456 9764
rect 11472 9820 11536 9824
rect 11472 9764 11476 9820
rect 11476 9764 11532 9820
rect 11532 9764 11536 9820
rect 11472 9760 11536 9764
rect 14659 9820 14723 9824
rect 14659 9764 14663 9820
rect 14663 9764 14719 9820
rect 14719 9764 14723 9820
rect 14659 9760 14723 9764
rect 14739 9820 14803 9824
rect 14739 9764 14743 9820
rect 14743 9764 14799 9820
rect 14799 9764 14803 9820
rect 14739 9760 14803 9764
rect 14819 9820 14883 9824
rect 14819 9764 14823 9820
rect 14823 9764 14879 9820
rect 14879 9764 14883 9820
rect 14819 9760 14883 9764
rect 14899 9820 14963 9824
rect 14899 9764 14903 9820
rect 14903 9764 14959 9820
rect 14959 9764 14963 9820
rect 14899 9760 14963 9764
rect 2665 9276 2729 9280
rect 2665 9220 2669 9276
rect 2669 9220 2725 9276
rect 2725 9220 2729 9276
rect 2665 9216 2729 9220
rect 2745 9276 2809 9280
rect 2745 9220 2749 9276
rect 2749 9220 2805 9276
rect 2805 9220 2809 9276
rect 2745 9216 2809 9220
rect 2825 9276 2889 9280
rect 2825 9220 2829 9276
rect 2829 9220 2885 9276
rect 2885 9220 2889 9276
rect 2825 9216 2889 9220
rect 2905 9276 2969 9280
rect 2905 9220 2909 9276
rect 2909 9220 2965 9276
rect 2965 9220 2969 9276
rect 2905 9216 2969 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 6332 9276 6396 9280
rect 6332 9220 6336 9276
rect 6336 9220 6392 9276
rect 6392 9220 6396 9276
rect 6332 9216 6396 9220
rect 9519 9276 9583 9280
rect 9519 9220 9523 9276
rect 9523 9220 9579 9276
rect 9579 9220 9583 9276
rect 9519 9216 9583 9220
rect 9599 9276 9663 9280
rect 9599 9220 9603 9276
rect 9603 9220 9659 9276
rect 9659 9220 9663 9276
rect 9599 9216 9663 9220
rect 9679 9276 9743 9280
rect 9679 9220 9683 9276
rect 9683 9220 9739 9276
rect 9739 9220 9743 9276
rect 9679 9216 9743 9220
rect 9759 9276 9823 9280
rect 9759 9220 9763 9276
rect 9763 9220 9819 9276
rect 9819 9220 9823 9276
rect 9759 9216 9823 9220
rect 10548 9148 10612 9212
rect 11652 9284 11716 9348
rect 12204 9480 12268 9484
rect 12204 9424 12254 9480
rect 12254 9424 12268 9480
rect 12204 9420 12268 9424
rect 12204 9284 12268 9348
rect 12946 9276 13010 9280
rect 12946 9220 12950 9276
rect 12950 9220 13006 9276
rect 13006 9220 13010 9276
rect 12946 9216 13010 9220
rect 13026 9276 13090 9280
rect 13026 9220 13030 9276
rect 13030 9220 13086 9276
rect 13086 9220 13090 9276
rect 13026 9216 13090 9220
rect 13106 9276 13170 9280
rect 13106 9220 13110 9276
rect 13110 9220 13166 9276
rect 13166 9220 13170 9276
rect 13106 9216 13170 9220
rect 13186 9276 13250 9280
rect 13186 9220 13190 9276
rect 13190 9220 13246 9276
rect 13246 9220 13250 9276
rect 13186 9216 13250 9220
rect 12756 9148 12820 9212
rect 11836 8740 11900 8804
rect 4378 8732 4442 8736
rect 4378 8676 4382 8732
rect 4382 8676 4438 8732
rect 4438 8676 4442 8732
rect 4378 8672 4442 8676
rect 4458 8732 4522 8736
rect 4458 8676 4462 8732
rect 4462 8676 4518 8732
rect 4518 8676 4522 8732
rect 4458 8672 4522 8676
rect 4538 8732 4602 8736
rect 4538 8676 4542 8732
rect 4542 8676 4598 8732
rect 4598 8676 4602 8732
rect 4538 8672 4602 8676
rect 4618 8732 4682 8736
rect 4618 8676 4622 8732
rect 4622 8676 4678 8732
rect 4678 8676 4682 8732
rect 4618 8672 4682 8676
rect 7805 8732 7869 8736
rect 7805 8676 7809 8732
rect 7809 8676 7865 8732
rect 7865 8676 7869 8732
rect 7805 8672 7869 8676
rect 7885 8732 7949 8736
rect 7885 8676 7889 8732
rect 7889 8676 7945 8732
rect 7945 8676 7949 8732
rect 7885 8672 7949 8676
rect 7965 8732 8029 8736
rect 7965 8676 7969 8732
rect 7969 8676 8025 8732
rect 8025 8676 8029 8732
rect 7965 8672 8029 8676
rect 8045 8732 8109 8736
rect 8045 8676 8049 8732
rect 8049 8676 8105 8732
rect 8105 8676 8109 8732
rect 8045 8672 8109 8676
rect 11232 8732 11296 8736
rect 11232 8676 11236 8732
rect 11236 8676 11292 8732
rect 11292 8676 11296 8732
rect 11232 8672 11296 8676
rect 11312 8732 11376 8736
rect 11312 8676 11316 8732
rect 11316 8676 11372 8732
rect 11372 8676 11376 8732
rect 11312 8672 11376 8676
rect 11392 8732 11456 8736
rect 11392 8676 11396 8732
rect 11396 8676 11452 8732
rect 11452 8676 11456 8732
rect 11392 8672 11456 8676
rect 11472 8732 11536 8736
rect 11472 8676 11476 8732
rect 11476 8676 11532 8732
rect 11532 8676 11536 8732
rect 11472 8672 11536 8676
rect 14659 8732 14723 8736
rect 14659 8676 14663 8732
rect 14663 8676 14719 8732
rect 14719 8676 14723 8732
rect 14659 8672 14723 8676
rect 14739 8732 14803 8736
rect 14739 8676 14743 8732
rect 14743 8676 14799 8732
rect 14799 8676 14803 8732
rect 14739 8672 14803 8676
rect 14819 8732 14883 8736
rect 14819 8676 14823 8732
rect 14823 8676 14879 8732
rect 14879 8676 14883 8732
rect 14819 8672 14883 8676
rect 14899 8732 14963 8736
rect 14899 8676 14903 8732
rect 14903 8676 14959 8732
rect 14959 8676 14963 8732
rect 14899 8672 14963 8676
rect 12204 8604 12268 8668
rect 13676 8256 13740 8260
rect 13676 8200 13726 8256
rect 13726 8200 13740 8256
rect 13676 8196 13740 8200
rect 2665 8188 2729 8192
rect 2665 8132 2669 8188
rect 2669 8132 2725 8188
rect 2725 8132 2729 8188
rect 2665 8128 2729 8132
rect 2745 8188 2809 8192
rect 2745 8132 2749 8188
rect 2749 8132 2805 8188
rect 2805 8132 2809 8188
rect 2745 8128 2809 8132
rect 2825 8188 2889 8192
rect 2825 8132 2829 8188
rect 2829 8132 2885 8188
rect 2885 8132 2889 8188
rect 2825 8128 2889 8132
rect 2905 8188 2969 8192
rect 2905 8132 2909 8188
rect 2909 8132 2965 8188
rect 2965 8132 2969 8188
rect 2905 8128 2969 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 6332 8188 6396 8192
rect 6332 8132 6336 8188
rect 6336 8132 6392 8188
rect 6392 8132 6396 8188
rect 6332 8128 6396 8132
rect 9519 8188 9583 8192
rect 9519 8132 9523 8188
rect 9523 8132 9579 8188
rect 9579 8132 9583 8188
rect 9519 8128 9583 8132
rect 9599 8188 9663 8192
rect 9599 8132 9603 8188
rect 9603 8132 9659 8188
rect 9659 8132 9663 8188
rect 9599 8128 9663 8132
rect 9679 8188 9743 8192
rect 9679 8132 9683 8188
rect 9683 8132 9739 8188
rect 9739 8132 9743 8188
rect 9679 8128 9743 8132
rect 9759 8188 9823 8192
rect 9759 8132 9763 8188
rect 9763 8132 9819 8188
rect 9819 8132 9823 8188
rect 9759 8128 9823 8132
rect 12946 8188 13010 8192
rect 12946 8132 12950 8188
rect 12950 8132 13006 8188
rect 13006 8132 13010 8188
rect 12946 8128 13010 8132
rect 13026 8188 13090 8192
rect 13026 8132 13030 8188
rect 13030 8132 13086 8188
rect 13086 8132 13090 8188
rect 13026 8128 13090 8132
rect 13106 8188 13170 8192
rect 13106 8132 13110 8188
rect 13110 8132 13166 8188
rect 13166 8132 13170 8188
rect 13106 8128 13170 8132
rect 13186 8188 13250 8192
rect 13186 8132 13190 8188
rect 13190 8132 13246 8188
rect 13246 8132 13250 8188
rect 13186 8128 13250 8132
rect 10548 7848 10612 7852
rect 10548 7792 10598 7848
rect 10598 7792 10612 7848
rect 10548 7788 10612 7792
rect 12572 7788 12636 7852
rect 4378 7644 4442 7648
rect 4378 7588 4382 7644
rect 4382 7588 4438 7644
rect 4438 7588 4442 7644
rect 4378 7584 4442 7588
rect 4458 7644 4522 7648
rect 4458 7588 4462 7644
rect 4462 7588 4518 7644
rect 4518 7588 4522 7644
rect 4458 7584 4522 7588
rect 4538 7644 4602 7648
rect 4538 7588 4542 7644
rect 4542 7588 4598 7644
rect 4598 7588 4602 7644
rect 4538 7584 4602 7588
rect 4618 7644 4682 7648
rect 4618 7588 4622 7644
rect 4622 7588 4678 7644
rect 4678 7588 4682 7644
rect 4618 7584 4682 7588
rect 7805 7644 7869 7648
rect 7805 7588 7809 7644
rect 7809 7588 7865 7644
rect 7865 7588 7869 7644
rect 7805 7584 7869 7588
rect 7885 7644 7949 7648
rect 7885 7588 7889 7644
rect 7889 7588 7945 7644
rect 7945 7588 7949 7644
rect 7885 7584 7949 7588
rect 7965 7644 8029 7648
rect 7965 7588 7969 7644
rect 7969 7588 8025 7644
rect 8025 7588 8029 7644
rect 7965 7584 8029 7588
rect 8045 7644 8109 7648
rect 8045 7588 8049 7644
rect 8049 7588 8105 7644
rect 8105 7588 8109 7644
rect 8045 7584 8109 7588
rect 11232 7644 11296 7648
rect 11232 7588 11236 7644
rect 11236 7588 11292 7644
rect 11292 7588 11296 7644
rect 11232 7584 11296 7588
rect 11312 7644 11376 7648
rect 11312 7588 11316 7644
rect 11316 7588 11372 7644
rect 11372 7588 11376 7644
rect 11312 7584 11376 7588
rect 11392 7644 11456 7648
rect 11392 7588 11396 7644
rect 11396 7588 11452 7644
rect 11452 7588 11456 7644
rect 11392 7584 11456 7588
rect 11472 7644 11536 7648
rect 11472 7588 11476 7644
rect 11476 7588 11532 7644
rect 11532 7588 11536 7644
rect 11472 7584 11536 7588
rect 14659 7644 14723 7648
rect 14659 7588 14663 7644
rect 14663 7588 14719 7644
rect 14719 7588 14723 7644
rect 14659 7584 14723 7588
rect 14739 7644 14803 7648
rect 14739 7588 14743 7644
rect 14743 7588 14799 7644
rect 14799 7588 14803 7644
rect 14739 7584 14803 7588
rect 14819 7644 14883 7648
rect 14819 7588 14823 7644
rect 14823 7588 14879 7644
rect 14879 7588 14883 7644
rect 14819 7584 14883 7588
rect 14899 7644 14963 7648
rect 14899 7588 14903 7644
rect 14903 7588 14959 7644
rect 14959 7588 14963 7644
rect 14899 7584 14963 7588
rect 2665 7100 2729 7104
rect 2665 7044 2669 7100
rect 2669 7044 2725 7100
rect 2725 7044 2729 7100
rect 2665 7040 2729 7044
rect 2745 7100 2809 7104
rect 2745 7044 2749 7100
rect 2749 7044 2805 7100
rect 2805 7044 2809 7100
rect 2745 7040 2809 7044
rect 2825 7100 2889 7104
rect 2825 7044 2829 7100
rect 2829 7044 2885 7100
rect 2885 7044 2889 7100
rect 2825 7040 2889 7044
rect 2905 7100 2969 7104
rect 2905 7044 2909 7100
rect 2909 7044 2965 7100
rect 2965 7044 2969 7100
rect 2905 7040 2969 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 6332 7100 6396 7104
rect 6332 7044 6336 7100
rect 6336 7044 6392 7100
rect 6392 7044 6396 7100
rect 6332 7040 6396 7044
rect 9519 7100 9583 7104
rect 9519 7044 9523 7100
rect 9523 7044 9579 7100
rect 9579 7044 9583 7100
rect 9519 7040 9583 7044
rect 9599 7100 9663 7104
rect 9599 7044 9603 7100
rect 9603 7044 9659 7100
rect 9659 7044 9663 7100
rect 9599 7040 9663 7044
rect 9679 7100 9743 7104
rect 9679 7044 9683 7100
rect 9683 7044 9739 7100
rect 9739 7044 9743 7100
rect 9679 7040 9743 7044
rect 9759 7100 9823 7104
rect 9759 7044 9763 7100
rect 9763 7044 9819 7100
rect 9819 7044 9823 7100
rect 9759 7040 9823 7044
rect 12946 7100 13010 7104
rect 12946 7044 12950 7100
rect 12950 7044 13006 7100
rect 13006 7044 13010 7100
rect 12946 7040 13010 7044
rect 13026 7100 13090 7104
rect 13026 7044 13030 7100
rect 13030 7044 13086 7100
rect 13086 7044 13090 7100
rect 13026 7040 13090 7044
rect 13106 7100 13170 7104
rect 13106 7044 13110 7100
rect 13110 7044 13166 7100
rect 13166 7044 13170 7100
rect 13106 7040 13170 7044
rect 13186 7100 13250 7104
rect 13186 7044 13190 7100
rect 13190 7044 13246 7100
rect 13246 7044 13250 7100
rect 13186 7040 13250 7044
rect 5212 6836 5276 6900
rect 4378 6556 4442 6560
rect 4378 6500 4382 6556
rect 4382 6500 4438 6556
rect 4438 6500 4442 6556
rect 4378 6496 4442 6500
rect 4458 6556 4522 6560
rect 4458 6500 4462 6556
rect 4462 6500 4518 6556
rect 4518 6500 4522 6556
rect 4458 6496 4522 6500
rect 4538 6556 4602 6560
rect 4538 6500 4542 6556
rect 4542 6500 4598 6556
rect 4598 6500 4602 6556
rect 4538 6496 4602 6500
rect 4618 6556 4682 6560
rect 4618 6500 4622 6556
rect 4622 6500 4678 6556
rect 4678 6500 4682 6556
rect 4618 6496 4682 6500
rect 7805 6556 7869 6560
rect 7805 6500 7809 6556
rect 7809 6500 7865 6556
rect 7865 6500 7869 6556
rect 7805 6496 7869 6500
rect 7885 6556 7949 6560
rect 7885 6500 7889 6556
rect 7889 6500 7945 6556
rect 7945 6500 7949 6556
rect 7885 6496 7949 6500
rect 7965 6556 8029 6560
rect 7965 6500 7969 6556
rect 7969 6500 8025 6556
rect 8025 6500 8029 6556
rect 7965 6496 8029 6500
rect 8045 6556 8109 6560
rect 8045 6500 8049 6556
rect 8049 6500 8105 6556
rect 8105 6500 8109 6556
rect 8045 6496 8109 6500
rect 11232 6556 11296 6560
rect 11232 6500 11236 6556
rect 11236 6500 11292 6556
rect 11292 6500 11296 6556
rect 11232 6496 11296 6500
rect 11312 6556 11376 6560
rect 11312 6500 11316 6556
rect 11316 6500 11372 6556
rect 11372 6500 11376 6556
rect 11312 6496 11376 6500
rect 11392 6556 11456 6560
rect 11392 6500 11396 6556
rect 11396 6500 11452 6556
rect 11452 6500 11456 6556
rect 11392 6496 11456 6500
rect 11472 6556 11536 6560
rect 11472 6500 11476 6556
rect 11476 6500 11532 6556
rect 11532 6500 11536 6556
rect 11472 6496 11536 6500
rect 14659 6556 14723 6560
rect 14659 6500 14663 6556
rect 14663 6500 14719 6556
rect 14719 6500 14723 6556
rect 14659 6496 14723 6500
rect 14739 6556 14803 6560
rect 14739 6500 14743 6556
rect 14743 6500 14799 6556
rect 14799 6500 14803 6556
rect 14739 6496 14803 6500
rect 14819 6556 14883 6560
rect 14819 6500 14823 6556
rect 14823 6500 14879 6556
rect 14879 6500 14883 6556
rect 14819 6496 14883 6500
rect 14899 6556 14963 6560
rect 14899 6500 14903 6556
rect 14903 6500 14959 6556
rect 14959 6500 14963 6556
rect 14899 6496 14963 6500
rect 2665 6012 2729 6016
rect 2665 5956 2669 6012
rect 2669 5956 2725 6012
rect 2725 5956 2729 6012
rect 2665 5952 2729 5956
rect 2745 6012 2809 6016
rect 2745 5956 2749 6012
rect 2749 5956 2805 6012
rect 2805 5956 2809 6012
rect 2745 5952 2809 5956
rect 2825 6012 2889 6016
rect 2825 5956 2829 6012
rect 2829 5956 2885 6012
rect 2885 5956 2889 6012
rect 2825 5952 2889 5956
rect 2905 6012 2969 6016
rect 2905 5956 2909 6012
rect 2909 5956 2965 6012
rect 2965 5956 2969 6012
rect 2905 5952 2969 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 6332 6012 6396 6016
rect 6332 5956 6336 6012
rect 6336 5956 6392 6012
rect 6392 5956 6396 6012
rect 6332 5952 6396 5956
rect 9519 6012 9583 6016
rect 9519 5956 9523 6012
rect 9523 5956 9579 6012
rect 9579 5956 9583 6012
rect 9519 5952 9583 5956
rect 9599 6012 9663 6016
rect 9599 5956 9603 6012
rect 9603 5956 9659 6012
rect 9659 5956 9663 6012
rect 9599 5952 9663 5956
rect 9679 6012 9743 6016
rect 9679 5956 9683 6012
rect 9683 5956 9739 6012
rect 9739 5956 9743 6012
rect 9679 5952 9743 5956
rect 9759 6012 9823 6016
rect 9759 5956 9763 6012
rect 9763 5956 9819 6012
rect 9819 5956 9823 6012
rect 9759 5952 9823 5956
rect 11652 5884 11716 5948
rect 12572 6020 12636 6084
rect 12946 6012 13010 6016
rect 12946 5956 12950 6012
rect 12950 5956 13006 6012
rect 13006 5956 13010 6012
rect 12946 5952 13010 5956
rect 13026 6012 13090 6016
rect 13026 5956 13030 6012
rect 13030 5956 13086 6012
rect 13086 5956 13090 6012
rect 13026 5952 13090 5956
rect 13106 6012 13170 6016
rect 13106 5956 13110 6012
rect 13110 5956 13166 6012
rect 13166 5956 13170 6012
rect 13106 5952 13170 5956
rect 13186 6012 13250 6016
rect 13186 5956 13190 6012
rect 13190 5956 13246 6012
rect 13246 5956 13250 6012
rect 13186 5952 13250 5956
rect 4378 5468 4442 5472
rect 4378 5412 4382 5468
rect 4382 5412 4438 5468
rect 4438 5412 4442 5468
rect 4378 5408 4442 5412
rect 4458 5468 4522 5472
rect 4458 5412 4462 5468
rect 4462 5412 4518 5468
rect 4518 5412 4522 5468
rect 4458 5408 4522 5412
rect 4538 5468 4602 5472
rect 4538 5412 4542 5468
rect 4542 5412 4598 5468
rect 4598 5412 4602 5468
rect 4538 5408 4602 5412
rect 4618 5468 4682 5472
rect 4618 5412 4622 5468
rect 4622 5412 4678 5468
rect 4678 5412 4682 5468
rect 4618 5408 4682 5412
rect 7805 5468 7869 5472
rect 7805 5412 7809 5468
rect 7809 5412 7865 5468
rect 7865 5412 7869 5468
rect 7805 5408 7869 5412
rect 7885 5468 7949 5472
rect 7885 5412 7889 5468
rect 7889 5412 7945 5468
rect 7945 5412 7949 5468
rect 7885 5408 7949 5412
rect 7965 5468 8029 5472
rect 7965 5412 7969 5468
rect 7969 5412 8025 5468
rect 8025 5412 8029 5468
rect 7965 5408 8029 5412
rect 8045 5468 8109 5472
rect 8045 5412 8049 5468
rect 8049 5412 8105 5468
rect 8105 5412 8109 5468
rect 8045 5408 8109 5412
rect 11232 5468 11296 5472
rect 11232 5412 11236 5468
rect 11236 5412 11292 5468
rect 11292 5412 11296 5468
rect 11232 5408 11296 5412
rect 11312 5468 11376 5472
rect 11312 5412 11316 5468
rect 11316 5412 11372 5468
rect 11372 5412 11376 5468
rect 11312 5408 11376 5412
rect 11392 5468 11456 5472
rect 11392 5412 11396 5468
rect 11396 5412 11452 5468
rect 11452 5412 11456 5468
rect 11392 5408 11456 5412
rect 11472 5468 11536 5472
rect 11472 5412 11476 5468
rect 11476 5412 11532 5468
rect 11532 5412 11536 5468
rect 11472 5408 11536 5412
rect 10732 5204 10796 5268
rect 14659 5468 14723 5472
rect 14659 5412 14663 5468
rect 14663 5412 14719 5468
rect 14719 5412 14723 5468
rect 14659 5408 14723 5412
rect 14739 5468 14803 5472
rect 14739 5412 14743 5468
rect 14743 5412 14799 5468
rect 14799 5412 14803 5468
rect 14739 5408 14803 5412
rect 14819 5468 14883 5472
rect 14819 5412 14823 5468
rect 14823 5412 14879 5468
rect 14879 5412 14883 5468
rect 14819 5408 14883 5412
rect 14899 5468 14963 5472
rect 14899 5412 14903 5468
rect 14903 5412 14959 5468
rect 14959 5412 14963 5468
rect 14899 5408 14963 5412
rect 2665 4924 2729 4928
rect 2665 4868 2669 4924
rect 2669 4868 2725 4924
rect 2725 4868 2729 4924
rect 2665 4864 2729 4868
rect 2745 4924 2809 4928
rect 2745 4868 2749 4924
rect 2749 4868 2805 4924
rect 2805 4868 2809 4924
rect 2745 4864 2809 4868
rect 2825 4924 2889 4928
rect 2825 4868 2829 4924
rect 2829 4868 2885 4924
rect 2885 4868 2889 4924
rect 2825 4864 2889 4868
rect 2905 4924 2969 4928
rect 2905 4868 2909 4924
rect 2909 4868 2965 4924
rect 2965 4868 2969 4924
rect 2905 4864 2969 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 6332 4924 6396 4928
rect 6332 4868 6336 4924
rect 6336 4868 6392 4924
rect 6392 4868 6396 4924
rect 6332 4864 6396 4868
rect 9519 4924 9583 4928
rect 9519 4868 9523 4924
rect 9523 4868 9579 4924
rect 9579 4868 9583 4924
rect 9519 4864 9583 4868
rect 9599 4924 9663 4928
rect 9599 4868 9603 4924
rect 9603 4868 9659 4924
rect 9659 4868 9663 4924
rect 9599 4864 9663 4868
rect 9679 4924 9743 4928
rect 9679 4868 9683 4924
rect 9683 4868 9739 4924
rect 9739 4868 9743 4924
rect 9679 4864 9743 4868
rect 9759 4924 9823 4928
rect 9759 4868 9763 4924
rect 9763 4868 9819 4924
rect 9819 4868 9823 4924
rect 9759 4864 9823 4868
rect 12946 4924 13010 4928
rect 12946 4868 12950 4924
rect 12950 4868 13006 4924
rect 13006 4868 13010 4924
rect 12946 4864 13010 4868
rect 13026 4924 13090 4928
rect 13026 4868 13030 4924
rect 13030 4868 13086 4924
rect 13086 4868 13090 4924
rect 13026 4864 13090 4868
rect 13106 4924 13170 4928
rect 13106 4868 13110 4924
rect 13110 4868 13166 4924
rect 13166 4868 13170 4924
rect 13106 4864 13170 4868
rect 13186 4924 13250 4928
rect 13186 4868 13190 4924
rect 13190 4868 13246 4924
rect 13246 4868 13250 4924
rect 13186 4864 13250 4868
rect 4378 4380 4442 4384
rect 4378 4324 4382 4380
rect 4382 4324 4438 4380
rect 4438 4324 4442 4380
rect 4378 4320 4442 4324
rect 4458 4380 4522 4384
rect 4458 4324 4462 4380
rect 4462 4324 4518 4380
rect 4518 4324 4522 4380
rect 4458 4320 4522 4324
rect 4538 4380 4602 4384
rect 4538 4324 4542 4380
rect 4542 4324 4598 4380
rect 4598 4324 4602 4380
rect 4538 4320 4602 4324
rect 4618 4380 4682 4384
rect 4618 4324 4622 4380
rect 4622 4324 4678 4380
rect 4678 4324 4682 4380
rect 4618 4320 4682 4324
rect 7805 4380 7869 4384
rect 7805 4324 7809 4380
rect 7809 4324 7865 4380
rect 7865 4324 7869 4380
rect 7805 4320 7869 4324
rect 7885 4380 7949 4384
rect 7885 4324 7889 4380
rect 7889 4324 7945 4380
rect 7945 4324 7949 4380
rect 7885 4320 7949 4324
rect 7965 4380 8029 4384
rect 7965 4324 7969 4380
rect 7969 4324 8025 4380
rect 8025 4324 8029 4380
rect 7965 4320 8029 4324
rect 8045 4380 8109 4384
rect 8045 4324 8049 4380
rect 8049 4324 8105 4380
rect 8105 4324 8109 4380
rect 8045 4320 8109 4324
rect 11232 4380 11296 4384
rect 11232 4324 11236 4380
rect 11236 4324 11292 4380
rect 11292 4324 11296 4380
rect 11232 4320 11296 4324
rect 11312 4380 11376 4384
rect 11312 4324 11316 4380
rect 11316 4324 11372 4380
rect 11372 4324 11376 4380
rect 11312 4320 11376 4324
rect 11392 4380 11456 4384
rect 11392 4324 11396 4380
rect 11396 4324 11452 4380
rect 11452 4324 11456 4380
rect 11392 4320 11456 4324
rect 11472 4380 11536 4384
rect 11472 4324 11476 4380
rect 11476 4324 11532 4380
rect 11532 4324 11536 4380
rect 11472 4320 11536 4324
rect 14659 4380 14723 4384
rect 14659 4324 14663 4380
rect 14663 4324 14719 4380
rect 14719 4324 14723 4380
rect 14659 4320 14723 4324
rect 14739 4380 14803 4384
rect 14739 4324 14743 4380
rect 14743 4324 14799 4380
rect 14799 4324 14803 4380
rect 14739 4320 14803 4324
rect 14819 4380 14883 4384
rect 14819 4324 14823 4380
rect 14823 4324 14879 4380
rect 14879 4324 14883 4380
rect 14819 4320 14883 4324
rect 14899 4380 14963 4384
rect 14899 4324 14903 4380
rect 14903 4324 14959 4380
rect 14959 4324 14963 4380
rect 14899 4320 14963 4324
rect 8708 3980 8772 4044
rect 2665 3836 2729 3840
rect 2665 3780 2669 3836
rect 2669 3780 2725 3836
rect 2725 3780 2729 3836
rect 2665 3776 2729 3780
rect 2745 3836 2809 3840
rect 2745 3780 2749 3836
rect 2749 3780 2805 3836
rect 2805 3780 2809 3836
rect 2745 3776 2809 3780
rect 2825 3836 2889 3840
rect 2825 3780 2829 3836
rect 2829 3780 2885 3836
rect 2885 3780 2889 3836
rect 2825 3776 2889 3780
rect 2905 3836 2969 3840
rect 2905 3780 2909 3836
rect 2909 3780 2965 3836
rect 2965 3780 2969 3836
rect 2905 3776 2969 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 6332 3836 6396 3840
rect 6332 3780 6336 3836
rect 6336 3780 6392 3836
rect 6392 3780 6396 3836
rect 6332 3776 6396 3780
rect 9519 3836 9583 3840
rect 9519 3780 9523 3836
rect 9523 3780 9579 3836
rect 9579 3780 9583 3836
rect 9519 3776 9583 3780
rect 9599 3836 9663 3840
rect 9599 3780 9603 3836
rect 9603 3780 9659 3836
rect 9659 3780 9663 3836
rect 9599 3776 9663 3780
rect 9679 3836 9743 3840
rect 9679 3780 9683 3836
rect 9683 3780 9739 3836
rect 9739 3780 9743 3836
rect 9679 3776 9743 3780
rect 9759 3836 9823 3840
rect 9759 3780 9763 3836
rect 9763 3780 9819 3836
rect 9819 3780 9823 3836
rect 9759 3776 9823 3780
rect 12946 3836 13010 3840
rect 12946 3780 12950 3836
rect 12950 3780 13006 3836
rect 13006 3780 13010 3836
rect 12946 3776 13010 3780
rect 13026 3836 13090 3840
rect 13026 3780 13030 3836
rect 13030 3780 13086 3836
rect 13086 3780 13090 3836
rect 13026 3776 13090 3780
rect 13106 3836 13170 3840
rect 13106 3780 13110 3836
rect 13110 3780 13166 3836
rect 13166 3780 13170 3836
rect 13106 3776 13170 3780
rect 13186 3836 13250 3840
rect 13186 3780 13190 3836
rect 13190 3780 13246 3836
rect 13246 3780 13250 3836
rect 13186 3776 13250 3780
rect 4378 3292 4442 3296
rect 4378 3236 4382 3292
rect 4382 3236 4438 3292
rect 4438 3236 4442 3292
rect 4378 3232 4442 3236
rect 4458 3292 4522 3296
rect 4458 3236 4462 3292
rect 4462 3236 4518 3292
rect 4518 3236 4522 3292
rect 4458 3232 4522 3236
rect 4538 3292 4602 3296
rect 4538 3236 4542 3292
rect 4542 3236 4598 3292
rect 4598 3236 4602 3292
rect 4538 3232 4602 3236
rect 4618 3292 4682 3296
rect 4618 3236 4622 3292
rect 4622 3236 4678 3292
rect 4678 3236 4682 3292
rect 4618 3232 4682 3236
rect 7805 3292 7869 3296
rect 7805 3236 7809 3292
rect 7809 3236 7865 3292
rect 7865 3236 7869 3292
rect 7805 3232 7869 3236
rect 7885 3292 7949 3296
rect 7885 3236 7889 3292
rect 7889 3236 7945 3292
rect 7945 3236 7949 3292
rect 7885 3232 7949 3236
rect 7965 3292 8029 3296
rect 7965 3236 7969 3292
rect 7969 3236 8025 3292
rect 8025 3236 8029 3292
rect 7965 3232 8029 3236
rect 8045 3292 8109 3296
rect 8045 3236 8049 3292
rect 8049 3236 8105 3292
rect 8105 3236 8109 3292
rect 8045 3232 8109 3236
rect 11232 3292 11296 3296
rect 11232 3236 11236 3292
rect 11236 3236 11292 3292
rect 11292 3236 11296 3292
rect 11232 3232 11296 3236
rect 11312 3292 11376 3296
rect 11312 3236 11316 3292
rect 11316 3236 11372 3292
rect 11372 3236 11376 3292
rect 11312 3232 11376 3236
rect 11392 3292 11456 3296
rect 11392 3236 11396 3292
rect 11396 3236 11452 3292
rect 11452 3236 11456 3292
rect 11392 3232 11456 3236
rect 11472 3292 11536 3296
rect 11472 3236 11476 3292
rect 11476 3236 11532 3292
rect 11532 3236 11536 3292
rect 11472 3232 11536 3236
rect 14659 3292 14723 3296
rect 14659 3236 14663 3292
rect 14663 3236 14719 3292
rect 14719 3236 14723 3292
rect 14659 3232 14723 3236
rect 14739 3292 14803 3296
rect 14739 3236 14743 3292
rect 14743 3236 14799 3292
rect 14799 3236 14803 3292
rect 14739 3232 14803 3236
rect 14819 3292 14883 3296
rect 14819 3236 14823 3292
rect 14823 3236 14879 3292
rect 14879 3236 14883 3292
rect 14819 3232 14883 3236
rect 14899 3292 14963 3296
rect 14899 3236 14903 3292
rect 14903 3236 14959 3292
rect 14959 3236 14963 3292
rect 14899 3232 14963 3236
rect 2665 2748 2729 2752
rect 2665 2692 2669 2748
rect 2669 2692 2725 2748
rect 2725 2692 2729 2748
rect 2665 2688 2729 2692
rect 2745 2748 2809 2752
rect 2745 2692 2749 2748
rect 2749 2692 2805 2748
rect 2805 2692 2809 2748
rect 2745 2688 2809 2692
rect 2825 2748 2889 2752
rect 2825 2692 2829 2748
rect 2829 2692 2885 2748
rect 2885 2692 2889 2748
rect 2825 2688 2889 2692
rect 2905 2748 2969 2752
rect 2905 2692 2909 2748
rect 2909 2692 2965 2748
rect 2965 2692 2969 2748
rect 2905 2688 2969 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 6332 2748 6396 2752
rect 6332 2692 6336 2748
rect 6336 2692 6392 2748
rect 6392 2692 6396 2748
rect 6332 2688 6396 2692
rect 9519 2748 9583 2752
rect 9519 2692 9523 2748
rect 9523 2692 9579 2748
rect 9579 2692 9583 2748
rect 9519 2688 9583 2692
rect 9599 2748 9663 2752
rect 9599 2692 9603 2748
rect 9603 2692 9659 2748
rect 9659 2692 9663 2748
rect 9599 2688 9663 2692
rect 9679 2748 9743 2752
rect 9679 2692 9683 2748
rect 9683 2692 9739 2748
rect 9739 2692 9743 2748
rect 9679 2688 9743 2692
rect 9759 2748 9823 2752
rect 9759 2692 9763 2748
rect 9763 2692 9819 2748
rect 9819 2692 9823 2748
rect 9759 2688 9823 2692
rect 12946 2748 13010 2752
rect 12946 2692 12950 2748
rect 12950 2692 13006 2748
rect 13006 2692 13010 2748
rect 12946 2688 13010 2692
rect 13026 2748 13090 2752
rect 13026 2692 13030 2748
rect 13030 2692 13086 2748
rect 13086 2692 13090 2748
rect 13026 2688 13090 2692
rect 13106 2748 13170 2752
rect 13106 2692 13110 2748
rect 13110 2692 13166 2748
rect 13166 2692 13170 2748
rect 13106 2688 13170 2692
rect 13186 2748 13250 2752
rect 13186 2692 13190 2748
rect 13190 2692 13246 2748
rect 13246 2692 13250 2748
rect 13186 2688 13250 2692
rect 5764 2680 5828 2684
rect 5764 2624 5814 2680
rect 5814 2624 5828 2680
rect 5764 2620 5828 2624
rect 6684 2680 6748 2684
rect 6684 2624 6698 2680
rect 6698 2624 6748 2680
rect 6684 2620 6748 2624
rect 7420 2620 7484 2684
rect 10916 2680 10980 2684
rect 10916 2624 10930 2680
rect 10930 2624 10980 2680
rect 10916 2620 10980 2624
rect 4378 2204 4442 2208
rect 4378 2148 4382 2204
rect 4382 2148 4438 2204
rect 4438 2148 4442 2204
rect 4378 2144 4442 2148
rect 4458 2204 4522 2208
rect 4458 2148 4462 2204
rect 4462 2148 4518 2204
rect 4518 2148 4522 2204
rect 4458 2144 4522 2148
rect 4538 2204 4602 2208
rect 4538 2148 4542 2204
rect 4542 2148 4598 2204
rect 4598 2148 4602 2204
rect 4538 2144 4602 2148
rect 4618 2204 4682 2208
rect 4618 2148 4622 2204
rect 4622 2148 4678 2204
rect 4678 2148 4682 2204
rect 4618 2144 4682 2148
rect 7805 2204 7869 2208
rect 7805 2148 7809 2204
rect 7809 2148 7865 2204
rect 7865 2148 7869 2204
rect 7805 2144 7869 2148
rect 7885 2204 7949 2208
rect 7885 2148 7889 2204
rect 7889 2148 7945 2204
rect 7945 2148 7949 2204
rect 7885 2144 7949 2148
rect 7965 2204 8029 2208
rect 7965 2148 7969 2204
rect 7969 2148 8025 2204
rect 8025 2148 8029 2204
rect 7965 2144 8029 2148
rect 8045 2204 8109 2208
rect 8045 2148 8049 2204
rect 8049 2148 8105 2204
rect 8105 2148 8109 2204
rect 8045 2144 8109 2148
rect 11232 2204 11296 2208
rect 11232 2148 11236 2204
rect 11236 2148 11292 2204
rect 11292 2148 11296 2204
rect 11232 2144 11296 2148
rect 11312 2204 11376 2208
rect 11312 2148 11316 2204
rect 11316 2148 11372 2204
rect 11372 2148 11376 2204
rect 11312 2144 11376 2148
rect 11392 2204 11456 2208
rect 11392 2148 11396 2204
rect 11396 2148 11452 2204
rect 11452 2148 11456 2204
rect 11392 2144 11456 2148
rect 11472 2204 11536 2208
rect 11472 2148 11476 2204
rect 11476 2148 11532 2204
rect 11532 2148 11536 2204
rect 11472 2144 11536 2148
rect 14659 2204 14723 2208
rect 14659 2148 14663 2204
rect 14663 2148 14719 2204
rect 14719 2148 14723 2204
rect 14659 2144 14723 2148
rect 14739 2204 14803 2208
rect 14739 2148 14743 2204
rect 14743 2148 14799 2204
rect 14799 2148 14803 2204
rect 14739 2144 14803 2148
rect 14819 2204 14883 2208
rect 14819 2148 14823 2204
rect 14823 2148 14879 2204
rect 14879 2148 14883 2204
rect 14819 2144 14883 2148
rect 14899 2204 14963 2208
rect 14899 2148 14903 2204
rect 14903 2148 14959 2204
rect 14959 2148 14963 2204
rect 14899 2144 14963 2148
rect 5396 1804 5460 1868
rect 2665 1660 2729 1664
rect 2665 1604 2669 1660
rect 2669 1604 2725 1660
rect 2725 1604 2729 1660
rect 2665 1600 2729 1604
rect 2745 1660 2809 1664
rect 2745 1604 2749 1660
rect 2749 1604 2805 1660
rect 2805 1604 2809 1660
rect 2745 1600 2809 1604
rect 2825 1660 2889 1664
rect 2825 1604 2829 1660
rect 2829 1604 2885 1660
rect 2885 1604 2889 1660
rect 2825 1600 2889 1604
rect 2905 1660 2969 1664
rect 2905 1604 2909 1660
rect 2909 1604 2965 1660
rect 2965 1604 2969 1660
rect 2905 1600 2969 1604
rect 6092 1660 6156 1664
rect 6092 1604 6096 1660
rect 6096 1604 6152 1660
rect 6152 1604 6156 1660
rect 6092 1600 6156 1604
rect 6172 1660 6236 1664
rect 6172 1604 6176 1660
rect 6176 1604 6232 1660
rect 6232 1604 6236 1660
rect 6172 1600 6236 1604
rect 6252 1660 6316 1664
rect 6252 1604 6256 1660
rect 6256 1604 6312 1660
rect 6312 1604 6316 1660
rect 6252 1600 6316 1604
rect 6332 1660 6396 1664
rect 6332 1604 6336 1660
rect 6336 1604 6392 1660
rect 6392 1604 6396 1660
rect 6332 1600 6396 1604
rect 9519 1660 9583 1664
rect 9519 1604 9523 1660
rect 9523 1604 9579 1660
rect 9579 1604 9583 1660
rect 9519 1600 9583 1604
rect 9599 1660 9663 1664
rect 9599 1604 9603 1660
rect 9603 1604 9659 1660
rect 9659 1604 9663 1660
rect 9599 1600 9663 1604
rect 9679 1660 9743 1664
rect 9679 1604 9683 1660
rect 9683 1604 9739 1660
rect 9739 1604 9743 1660
rect 9679 1600 9743 1604
rect 9759 1660 9823 1664
rect 9759 1604 9763 1660
rect 9763 1604 9819 1660
rect 9819 1604 9823 1660
rect 9759 1600 9823 1604
rect 12946 1660 13010 1664
rect 12946 1604 12950 1660
rect 12950 1604 13006 1660
rect 13006 1604 13010 1660
rect 12946 1600 13010 1604
rect 13026 1660 13090 1664
rect 13026 1604 13030 1660
rect 13030 1604 13086 1660
rect 13086 1604 13090 1660
rect 13026 1600 13090 1604
rect 13106 1660 13170 1664
rect 13106 1604 13110 1660
rect 13110 1604 13166 1660
rect 13166 1604 13170 1660
rect 13106 1600 13170 1604
rect 13186 1660 13250 1664
rect 13186 1604 13190 1660
rect 13190 1604 13246 1660
rect 13246 1604 13250 1660
rect 13186 1600 13250 1604
rect 4378 1116 4442 1120
rect 4378 1060 4382 1116
rect 4382 1060 4438 1116
rect 4438 1060 4442 1116
rect 4378 1056 4442 1060
rect 4458 1116 4522 1120
rect 4458 1060 4462 1116
rect 4462 1060 4518 1116
rect 4518 1060 4522 1116
rect 4458 1056 4522 1060
rect 4538 1116 4602 1120
rect 4538 1060 4542 1116
rect 4542 1060 4598 1116
rect 4598 1060 4602 1116
rect 4538 1056 4602 1060
rect 4618 1116 4682 1120
rect 4618 1060 4622 1116
rect 4622 1060 4678 1116
rect 4678 1060 4682 1116
rect 4618 1056 4682 1060
rect 7805 1116 7869 1120
rect 7805 1060 7809 1116
rect 7809 1060 7865 1116
rect 7865 1060 7869 1116
rect 7805 1056 7869 1060
rect 7885 1116 7949 1120
rect 7885 1060 7889 1116
rect 7889 1060 7945 1116
rect 7945 1060 7949 1116
rect 7885 1056 7949 1060
rect 7965 1116 8029 1120
rect 7965 1060 7969 1116
rect 7969 1060 8025 1116
rect 8025 1060 8029 1116
rect 7965 1056 8029 1060
rect 8045 1116 8109 1120
rect 8045 1060 8049 1116
rect 8049 1060 8105 1116
rect 8105 1060 8109 1116
rect 8045 1056 8109 1060
rect 11232 1116 11296 1120
rect 11232 1060 11236 1116
rect 11236 1060 11292 1116
rect 11292 1060 11296 1116
rect 11232 1056 11296 1060
rect 11312 1116 11376 1120
rect 11312 1060 11316 1116
rect 11316 1060 11372 1116
rect 11372 1060 11376 1116
rect 11312 1056 11376 1060
rect 11392 1116 11456 1120
rect 11392 1060 11396 1116
rect 11396 1060 11452 1116
rect 11452 1060 11456 1116
rect 11392 1056 11456 1060
rect 11472 1116 11536 1120
rect 11472 1060 11476 1116
rect 11476 1060 11532 1116
rect 11532 1060 11536 1116
rect 11472 1056 11536 1060
rect 14659 1116 14723 1120
rect 14659 1060 14663 1116
rect 14663 1060 14719 1116
rect 14719 1060 14723 1116
rect 14659 1056 14723 1060
rect 14739 1116 14803 1120
rect 14739 1060 14743 1116
rect 14743 1060 14799 1116
rect 14799 1060 14803 1116
rect 14739 1056 14803 1060
rect 14819 1116 14883 1120
rect 14819 1060 14823 1116
rect 14823 1060 14879 1116
rect 14879 1060 14883 1116
rect 14819 1056 14883 1060
rect 14899 1116 14963 1120
rect 14899 1060 14903 1116
rect 14903 1060 14959 1116
rect 14959 1060 14963 1116
rect 14899 1056 14963 1060
<< metal4 >>
rect 2657 43008 2977 43568
rect 2657 42944 2665 43008
rect 2729 42944 2745 43008
rect 2809 42944 2825 43008
rect 2889 42944 2905 43008
rect 2969 42944 2977 43008
rect 2657 41920 2977 42944
rect 2657 41856 2665 41920
rect 2729 41856 2745 41920
rect 2809 41856 2825 41920
rect 2889 41856 2905 41920
rect 2969 41856 2977 41920
rect 2657 40832 2977 41856
rect 4370 43552 4690 43568
rect 4370 43488 4378 43552
rect 4442 43488 4458 43552
rect 4522 43488 4538 43552
rect 4602 43488 4618 43552
rect 4682 43488 4690 43552
rect 4370 42464 4690 43488
rect 4370 42400 4378 42464
rect 4442 42400 4458 42464
rect 4522 42400 4538 42464
rect 4602 42400 4618 42464
rect 4682 42400 4690 42464
rect 3923 41580 3989 41581
rect 3923 41516 3924 41580
rect 3988 41516 3989 41580
rect 3923 41515 3989 41516
rect 2657 40768 2665 40832
rect 2729 40768 2745 40832
rect 2809 40768 2825 40832
rect 2889 40768 2905 40832
rect 2969 40768 2977 40832
rect 2657 39744 2977 40768
rect 2657 39680 2665 39744
rect 2729 39680 2745 39744
rect 2809 39680 2825 39744
rect 2889 39680 2905 39744
rect 2969 39680 2977 39744
rect 2657 38656 2977 39680
rect 2657 38592 2665 38656
rect 2729 38592 2745 38656
rect 2809 38592 2825 38656
rect 2889 38592 2905 38656
rect 2969 38592 2977 38656
rect 2657 37568 2977 38592
rect 2657 37504 2665 37568
rect 2729 37504 2745 37568
rect 2809 37504 2825 37568
rect 2889 37504 2905 37568
rect 2969 37504 2977 37568
rect 2657 36480 2977 37504
rect 2657 36416 2665 36480
rect 2729 36416 2745 36480
rect 2809 36416 2825 36480
rect 2889 36416 2905 36480
rect 2969 36416 2977 36480
rect 2657 35392 2977 36416
rect 2657 35328 2665 35392
rect 2729 35328 2745 35392
rect 2809 35328 2825 35392
rect 2889 35328 2905 35392
rect 2969 35328 2977 35392
rect 2657 34304 2977 35328
rect 2657 34240 2665 34304
rect 2729 34240 2745 34304
rect 2809 34240 2825 34304
rect 2889 34240 2905 34304
rect 2969 34240 2977 34304
rect 2657 33216 2977 34240
rect 2657 33152 2665 33216
rect 2729 33152 2745 33216
rect 2809 33152 2825 33216
rect 2889 33152 2905 33216
rect 2969 33152 2977 33216
rect 2657 32128 2977 33152
rect 2657 32064 2665 32128
rect 2729 32064 2745 32128
rect 2809 32064 2825 32128
rect 2889 32064 2905 32128
rect 2969 32064 2977 32128
rect 2657 31040 2977 32064
rect 2657 30976 2665 31040
rect 2729 30976 2745 31040
rect 2809 30976 2825 31040
rect 2889 30976 2905 31040
rect 2969 30976 2977 31040
rect 2657 29952 2977 30976
rect 2657 29888 2665 29952
rect 2729 29888 2745 29952
rect 2809 29888 2825 29952
rect 2889 29888 2905 29952
rect 2969 29888 2977 29952
rect 2657 28864 2977 29888
rect 2657 28800 2665 28864
rect 2729 28800 2745 28864
rect 2809 28800 2825 28864
rect 2889 28800 2905 28864
rect 2969 28800 2977 28864
rect 2657 27776 2977 28800
rect 2657 27712 2665 27776
rect 2729 27712 2745 27776
rect 2809 27712 2825 27776
rect 2889 27712 2905 27776
rect 2969 27712 2977 27776
rect 1715 27708 1781 27709
rect 1715 27644 1716 27708
rect 1780 27644 1781 27708
rect 1715 27643 1781 27644
rect 1718 14109 1778 27643
rect 2657 26688 2977 27712
rect 2657 26624 2665 26688
rect 2729 26624 2745 26688
rect 2809 26624 2825 26688
rect 2889 26624 2905 26688
rect 2969 26624 2977 26688
rect 2657 25600 2977 26624
rect 2657 25536 2665 25600
rect 2729 25536 2745 25600
rect 2809 25536 2825 25600
rect 2889 25536 2905 25600
rect 2969 25536 2977 25600
rect 2657 24512 2977 25536
rect 2657 24448 2665 24512
rect 2729 24448 2745 24512
rect 2809 24448 2825 24512
rect 2889 24448 2905 24512
rect 2969 24448 2977 24512
rect 2657 23424 2977 24448
rect 2657 23360 2665 23424
rect 2729 23360 2745 23424
rect 2809 23360 2825 23424
rect 2889 23360 2905 23424
rect 2969 23360 2977 23424
rect 2657 22336 2977 23360
rect 2657 22272 2665 22336
rect 2729 22272 2745 22336
rect 2809 22272 2825 22336
rect 2889 22272 2905 22336
rect 2969 22272 2977 22336
rect 2657 21248 2977 22272
rect 2657 21184 2665 21248
rect 2729 21184 2745 21248
rect 2809 21184 2825 21248
rect 2889 21184 2905 21248
rect 2969 21184 2977 21248
rect 2657 20160 2977 21184
rect 2657 20096 2665 20160
rect 2729 20096 2745 20160
rect 2809 20096 2825 20160
rect 2889 20096 2905 20160
rect 2969 20096 2977 20160
rect 2657 19072 2977 20096
rect 2657 19008 2665 19072
rect 2729 19008 2745 19072
rect 2809 19008 2825 19072
rect 2889 19008 2905 19072
rect 2969 19008 2977 19072
rect 2657 17984 2977 19008
rect 2657 17920 2665 17984
rect 2729 17920 2745 17984
rect 2809 17920 2825 17984
rect 2889 17920 2905 17984
rect 2969 17920 2977 17984
rect 2657 16896 2977 17920
rect 2657 16832 2665 16896
rect 2729 16832 2745 16896
rect 2809 16832 2825 16896
rect 2889 16832 2905 16896
rect 2969 16832 2977 16896
rect 2657 15808 2977 16832
rect 2657 15744 2665 15808
rect 2729 15744 2745 15808
rect 2809 15744 2825 15808
rect 2889 15744 2905 15808
rect 2969 15744 2977 15808
rect 2657 14720 2977 15744
rect 2657 14656 2665 14720
rect 2729 14656 2745 14720
rect 2809 14656 2825 14720
rect 2889 14656 2905 14720
rect 2969 14656 2977 14720
rect 1715 14108 1781 14109
rect 1715 14044 1716 14108
rect 1780 14044 1781 14108
rect 1715 14043 1781 14044
rect 2657 13632 2977 14656
rect 2657 13568 2665 13632
rect 2729 13568 2745 13632
rect 2809 13568 2825 13632
rect 2889 13568 2905 13632
rect 2969 13568 2977 13632
rect 2657 12544 2977 13568
rect 3926 12885 3986 41515
rect 4370 41376 4690 42400
rect 6084 43008 6404 43568
rect 6084 42944 6092 43008
rect 6156 42944 6172 43008
rect 6236 42944 6252 43008
rect 6316 42944 6332 43008
rect 6396 42944 6404 43008
rect 5395 42124 5461 42125
rect 5395 42060 5396 42124
rect 5460 42060 5461 42124
rect 5395 42059 5461 42060
rect 4370 41312 4378 41376
rect 4442 41312 4458 41376
rect 4522 41312 4538 41376
rect 4602 41312 4618 41376
rect 4682 41312 4690 41376
rect 4370 40288 4690 41312
rect 4370 40224 4378 40288
rect 4442 40224 4458 40288
rect 4522 40224 4538 40288
rect 4602 40224 4618 40288
rect 4682 40224 4690 40288
rect 4370 39200 4690 40224
rect 4370 39136 4378 39200
rect 4442 39136 4458 39200
rect 4522 39136 4538 39200
rect 4602 39136 4618 39200
rect 4682 39136 4690 39200
rect 4370 38112 4690 39136
rect 4370 38048 4378 38112
rect 4442 38048 4458 38112
rect 4522 38048 4538 38112
rect 4602 38048 4618 38112
rect 4682 38048 4690 38112
rect 4370 37024 4690 38048
rect 4370 36960 4378 37024
rect 4442 36960 4458 37024
rect 4522 36960 4538 37024
rect 4602 36960 4618 37024
rect 4682 36960 4690 37024
rect 4370 35936 4690 36960
rect 4370 35872 4378 35936
rect 4442 35872 4458 35936
rect 4522 35872 4538 35936
rect 4602 35872 4618 35936
rect 4682 35872 4690 35936
rect 4370 34848 4690 35872
rect 4370 34784 4378 34848
rect 4442 34784 4458 34848
rect 4522 34784 4538 34848
rect 4602 34784 4618 34848
rect 4682 34784 4690 34848
rect 4370 33760 4690 34784
rect 4370 33696 4378 33760
rect 4442 33696 4458 33760
rect 4522 33696 4538 33760
rect 4602 33696 4618 33760
rect 4682 33696 4690 33760
rect 4370 32672 4690 33696
rect 4370 32608 4378 32672
rect 4442 32608 4458 32672
rect 4522 32608 4538 32672
rect 4602 32608 4618 32672
rect 4682 32608 4690 32672
rect 4370 31584 4690 32608
rect 4370 31520 4378 31584
rect 4442 31520 4458 31584
rect 4522 31520 4538 31584
rect 4602 31520 4618 31584
rect 4682 31520 4690 31584
rect 4370 30496 4690 31520
rect 4370 30432 4378 30496
rect 4442 30432 4458 30496
rect 4522 30432 4538 30496
rect 4602 30432 4618 30496
rect 4682 30432 4690 30496
rect 4370 29408 4690 30432
rect 4370 29344 4378 29408
rect 4442 29344 4458 29408
rect 4522 29344 4538 29408
rect 4602 29344 4618 29408
rect 4682 29344 4690 29408
rect 4370 28320 4690 29344
rect 4370 28256 4378 28320
rect 4442 28256 4458 28320
rect 4522 28256 4538 28320
rect 4602 28256 4618 28320
rect 4682 28256 4690 28320
rect 4370 27232 4690 28256
rect 4370 27168 4378 27232
rect 4442 27168 4458 27232
rect 4522 27168 4538 27232
rect 4602 27168 4618 27232
rect 4682 27168 4690 27232
rect 4370 26144 4690 27168
rect 5211 26484 5277 26485
rect 5211 26420 5212 26484
rect 5276 26420 5277 26484
rect 5211 26419 5277 26420
rect 4370 26080 4378 26144
rect 4442 26080 4458 26144
rect 4522 26080 4538 26144
rect 4602 26080 4618 26144
rect 4682 26080 4690 26144
rect 4370 25056 4690 26080
rect 4370 24992 4378 25056
rect 4442 24992 4458 25056
rect 4522 24992 4538 25056
rect 4602 24992 4618 25056
rect 4682 24992 4690 25056
rect 4370 23968 4690 24992
rect 4370 23904 4378 23968
rect 4442 23904 4458 23968
rect 4522 23904 4538 23968
rect 4602 23904 4618 23968
rect 4682 23904 4690 23968
rect 4370 22880 4690 23904
rect 4370 22816 4378 22880
rect 4442 22816 4458 22880
rect 4522 22816 4538 22880
rect 4602 22816 4618 22880
rect 4682 22816 4690 22880
rect 4370 21792 4690 22816
rect 4370 21728 4378 21792
rect 4442 21728 4458 21792
rect 4522 21728 4538 21792
rect 4602 21728 4618 21792
rect 4682 21728 4690 21792
rect 4370 20704 4690 21728
rect 4370 20640 4378 20704
rect 4442 20640 4458 20704
rect 4522 20640 4538 20704
rect 4602 20640 4618 20704
rect 4682 20640 4690 20704
rect 4370 19616 4690 20640
rect 4370 19552 4378 19616
rect 4442 19552 4458 19616
rect 4522 19552 4538 19616
rect 4602 19552 4618 19616
rect 4682 19552 4690 19616
rect 4370 18528 4690 19552
rect 4370 18464 4378 18528
rect 4442 18464 4458 18528
rect 4522 18464 4538 18528
rect 4602 18464 4618 18528
rect 4682 18464 4690 18528
rect 4370 17440 4690 18464
rect 4370 17376 4378 17440
rect 4442 17376 4458 17440
rect 4522 17376 4538 17440
rect 4602 17376 4618 17440
rect 4682 17376 4690 17440
rect 4370 16352 4690 17376
rect 4370 16288 4378 16352
rect 4442 16288 4458 16352
rect 4522 16288 4538 16352
rect 4602 16288 4618 16352
rect 4682 16288 4690 16352
rect 4370 15264 4690 16288
rect 4370 15200 4378 15264
rect 4442 15200 4458 15264
rect 4522 15200 4538 15264
rect 4602 15200 4618 15264
rect 4682 15200 4690 15264
rect 4370 14176 4690 15200
rect 4370 14112 4378 14176
rect 4442 14112 4458 14176
rect 4522 14112 4538 14176
rect 4602 14112 4618 14176
rect 4682 14112 4690 14176
rect 4370 13088 4690 14112
rect 4370 13024 4378 13088
rect 4442 13024 4458 13088
rect 4522 13024 4538 13088
rect 4602 13024 4618 13088
rect 4682 13024 4690 13088
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 2657 12480 2665 12544
rect 2729 12480 2745 12544
rect 2809 12480 2825 12544
rect 2889 12480 2905 12544
rect 2969 12480 2977 12544
rect 2657 11456 2977 12480
rect 2657 11392 2665 11456
rect 2729 11392 2745 11456
rect 2809 11392 2825 11456
rect 2889 11392 2905 11456
rect 2969 11392 2977 11456
rect 2657 10368 2977 11392
rect 2657 10304 2665 10368
rect 2729 10304 2745 10368
rect 2809 10304 2825 10368
rect 2889 10304 2905 10368
rect 2969 10304 2977 10368
rect 2657 9280 2977 10304
rect 2657 9216 2665 9280
rect 2729 9216 2745 9280
rect 2809 9216 2825 9280
rect 2889 9216 2905 9280
rect 2969 9216 2977 9280
rect 2657 8192 2977 9216
rect 2657 8128 2665 8192
rect 2729 8128 2745 8192
rect 2809 8128 2825 8192
rect 2889 8128 2905 8192
rect 2969 8128 2977 8192
rect 2657 7104 2977 8128
rect 2657 7040 2665 7104
rect 2729 7040 2745 7104
rect 2809 7040 2825 7104
rect 2889 7040 2905 7104
rect 2969 7040 2977 7104
rect 2657 6016 2977 7040
rect 2657 5952 2665 6016
rect 2729 5952 2745 6016
rect 2809 5952 2825 6016
rect 2889 5952 2905 6016
rect 2969 5952 2977 6016
rect 2657 4928 2977 5952
rect 2657 4864 2665 4928
rect 2729 4864 2745 4928
rect 2809 4864 2825 4928
rect 2889 4864 2905 4928
rect 2969 4864 2977 4928
rect 2657 3840 2977 4864
rect 2657 3776 2665 3840
rect 2729 3776 2745 3840
rect 2809 3776 2825 3840
rect 2889 3776 2905 3840
rect 2969 3776 2977 3840
rect 2657 2752 2977 3776
rect 2657 2688 2665 2752
rect 2729 2688 2745 2752
rect 2809 2688 2825 2752
rect 2889 2688 2905 2752
rect 2969 2688 2977 2752
rect 2657 1664 2977 2688
rect 2657 1600 2665 1664
rect 2729 1600 2745 1664
rect 2809 1600 2825 1664
rect 2889 1600 2905 1664
rect 2969 1600 2977 1664
rect 2657 1040 2977 1600
rect 4370 12000 4690 13024
rect 4370 11936 4378 12000
rect 4442 11936 4458 12000
rect 4522 11936 4538 12000
rect 4602 11936 4618 12000
rect 4682 11936 4690 12000
rect 4370 10912 4690 11936
rect 4370 10848 4378 10912
rect 4442 10848 4458 10912
rect 4522 10848 4538 10912
rect 4602 10848 4618 10912
rect 4682 10848 4690 10912
rect 4370 9824 4690 10848
rect 4370 9760 4378 9824
rect 4442 9760 4458 9824
rect 4522 9760 4538 9824
rect 4602 9760 4618 9824
rect 4682 9760 4690 9824
rect 4370 8736 4690 9760
rect 4370 8672 4378 8736
rect 4442 8672 4458 8736
rect 4522 8672 4538 8736
rect 4602 8672 4618 8736
rect 4682 8672 4690 8736
rect 4370 7648 4690 8672
rect 4370 7584 4378 7648
rect 4442 7584 4458 7648
rect 4522 7584 4538 7648
rect 4602 7584 4618 7648
rect 4682 7584 4690 7648
rect 4370 6560 4690 7584
rect 5214 6901 5274 26419
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 4370 6496 4378 6560
rect 4442 6496 4458 6560
rect 4522 6496 4538 6560
rect 4602 6496 4618 6560
rect 4682 6496 4690 6560
rect 4370 5472 4690 6496
rect 4370 5408 4378 5472
rect 4442 5408 4458 5472
rect 4522 5408 4538 5472
rect 4602 5408 4618 5472
rect 4682 5408 4690 5472
rect 4370 4384 4690 5408
rect 4370 4320 4378 4384
rect 4442 4320 4458 4384
rect 4522 4320 4538 4384
rect 4602 4320 4618 4384
rect 4682 4320 4690 4384
rect 4370 3296 4690 4320
rect 4370 3232 4378 3296
rect 4442 3232 4458 3296
rect 4522 3232 4538 3296
rect 4602 3232 4618 3296
rect 4682 3232 4690 3296
rect 4370 2208 4690 3232
rect 4370 2144 4378 2208
rect 4442 2144 4458 2208
rect 4522 2144 4538 2208
rect 4602 2144 4618 2208
rect 4682 2144 4690 2208
rect 4370 1120 4690 2144
rect 5398 1869 5458 42059
rect 6084 41920 6404 42944
rect 6084 41856 6092 41920
rect 6156 41856 6172 41920
rect 6236 41856 6252 41920
rect 6316 41856 6332 41920
rect 6396 41856 6404 41920
rect 5763 41852 5829 41853
rect 5763 41788 5764 41852
rect 5828 41788 5829 41852
rect 5763 41787 5829 41788
rect 5766 2685 5826 41787
rect 6084 40832 6404 41856
rect 7797 43552 8117 43568
rect 7797 43488 7805 43552
rect 7869 43488 7885 43552
rect 7949 43488 7965 43552
rect 8029 43488 8045 43552
rect 8109 43488 8117 43552
rect 7797 42464 8117 43488
rect 7797 42400 7805 42464
rect 7869 42400 7885 42464
rect 7949 42400 7965 42464
rect 8029 42400 8045 42464
rect 8109 42400 8117 42464
rect 6683 41852 6749 41853
rect 6683 41788 6684 41852
rect 6748 41788 6749 41852
rect 6683 41787 6749 41788
rect 7419 41852 7485 41853
rect 7419 41788 7420 41852
rect 7484 41788 7485 41852
rect 7419 41787 7485 41788
rect 6084 40768 6092 40832
rect 6156 40768 6172 40832
rect 6236 40768 6252 40832
rect 6316 40768 6332 40832
rect 6396 40768 6404 40832
rect 6084 39744 6404 40768
rect 6084 39680 6092 39744
rect 6156 39680 6172 39744
rect 6236 39680 6252 39744
rect 6316 39680 6332 39744
rect 6396 39680 6404 39744
rect 6084 38656 6404 39680
rect 6084 38592 6092 38656
rect 6156 38592 6172 38656
rect 6236 38592 6252 38656
rect 6316 38592 6332 38656
rect 6396 38592 6404 38656
rect 6084 37568 6404 38592
rect 6084 37504 6092 37568
rect 6156 37504 6172 37568
rect 6236 37504 6252 37568
rect 6316 37504 6332 37568
rect 6396 37504 6404 37568
rect 6084 36480 6404 37504
rect 6084 36416 6092 36480
rect 6156 36416 6172 36480
rect 6236 36416 6252 36480
rect 6316 36416 6332 36480
rect 6396 36416 6404 36480
rect 6084 35392 6404 36416
rect 6084 35328 6092 35392
rect 6156 35328 6172 35392
rect 6236 35328 6252 35392
rect 6316 35328 6332 35392
rect 6396 35328 6404 35392
rect 6084 34304 6404 35328
rect 6084 34240 6092 34304
rect 6156 34240 6172 34304
rect 6236 34240 6252 34304
rect 6316 34240 6332 34304
rect 6396 34240 6404 34304
rect 6084 33216 6404 34240
rect 6084 33152 6092 33216
rect 6156 33152 6172 33216
rect 6236 33152 6252 33216
rect 6316 33152 6332 33216
rect 6396 33152 6404 33216
rect 6084 32128 6404 33152
rect 6084 32064 6092 32128
rect 6156 32064 6172 32128
rect 6236 32064 6252 32128
rect 6316 32064 6332 32128
rect 6396 32064 6404 32128
rect 6084 31040 6404 32064
rect 6084 30976 6092 31040
rect 6156 30976 6172 31040
rect 6236 30976 6252 31040
rect 6316 30976 6332 31040
rect 6396 30976 6404 31040
rect 6084 29952 6404 30976
rect 6084 29888 6092 29952
rect 6156 29888 6172 29952
rect 6236 29888 6252 29952
rect 6316 29888 6332 29952
rect 6396 29888 6404 29952
rect 6084 28864 6404 29888
rect 6084 28800 6092 28864
rect 6156 28800 6172 28864
rect 6236 28800 6252 28864
rect 6316 28800 6332 28864
rect 6396 28800 6404 28864
rect 6084 27776 6404 28800
rect 6084 27712 6092 27776
rect 6156 27712 6172 27776
rect 6236 27712 6252 27776
rect 6316 27712 6332 27776
rect 6396 27712 6404 27776
rect 6084 26688 6404 27712
rect 6084 26624 6092 26688
rect 6156 26624 6172 26688
rect 6236 26624 6252 26688
rect 6316 26624 6332 26688
rect 6396 26624 6404 26688
rect 6084 25600 6404 26624
rect 6084 25536 6092 25600
rect 6156 25536 6172 25600
rect 6236 25536 6252 25600
rect 6316 25536 6332 25600
rect 6396 25536 6404 25600
rect 6084 24512 6404 25536
rect 6084 24448 6092 24512
rect 6156 24448 6172 24512
rect 6236 24448 6252 24512
rect 6316 24448 6332 24512
rect 6396 24448 6404 24512
rect 6084 23424 6404 24448
rect 6084 23360 6092 23424
rect 6156 23360 6172 23424
rect 6236 23360 6252 23424
rect 6316 23360 6332 23424
rect 6396 23360 6404 23424
rect 6084 22336 6404 23360
rect 6084 22272 6092 22336
rect 6156 22272 6172 22336
rect 6236 22272 6252 22336
rect 6316 22272 6332 22336
rect 6396 22272 6404 22336
rect 6084 21248 6404 22272
rect 6084 21184 6092 21248
rect 6156 21184 6172 21248
rect 6236 21184 6252 21248
rect 6316 21184 6332 21248
rect 6396 21184 6404 21248
rect 6084 20160 6404 21184
rect 6084 20096 6092 20160
rect 6156 20096 6172 20160
rect 6236 20096 6252 20160
rect 6316 20096 6332 20160
rect 6396 20096 6404 20160
rect 6084 19072 6404 20096
rect 6084 19008 6092 19072
rect 6156 19008 6172 19072
rect 6236 19008 6252 19072
rect 6316 19008 6332 19072
rect 6396 19008 6404 19072
rect 6084 17984 6404 19008
rect 6084 17920 6092 17984
rect 6156 17920 6172 17984
rect 6236 17920 6252 17984
rect 6316 17920 6332 17984
rect 6396 17920 6404 17984
rect 6084 16896 6404 17920
rect 6084 16832 6092 16896
rect 6156 16832 6172 16896
rect 6236 16832 6252 16896
rect 6316 16832 6332 16896
rect 6396 16832 6404 16896
rect 6084 15808 6404 16832
rect 6084 15744 6092 15808
rect 6156 15744 6172 15808
rect 6236 15744 6252 15808
rect 6316 15744 6332 15808
rect 6396 15744 6404 15808
rect 6084 14720 6404 15744
rect 6084 14656 6092 14720
rect 6156 14656 6172 14720
rect 6236 14656 6252 14720
rect 6316 14656 6332 14720
rect 6396 14656 6404 14720
rect 6084 13632 6404 14656
rect 6084 13568 6092 13632
rect 6156 13568 6172 13632
rect 6236 13568 6252 13632
rect 6316 13568 6332 13632
rect 6396 13568 6404 13632
rect 6084 12544 6404 13568
rect 6084 12480 6092 12544
rect 6156 12480 6172 12544
rect 6236 12480 6252 12544
rect 6316 12480 6332 12544
rect 6396 12480 6404 12544
rect 6084 11456 6404 12480
rect 6084 11392 6092 11456
rect 6156 11392 6172 11456
rect 6236 11392 6252 11456
rect 6316 11392 6332 11456
rect 6396 11392 6404 11456
rect 6084 10368 6404 11392
rect 6084 10304 6092 10368
rect 6156 10304 6172 10368
rect 6236 10304 6252 10368
rect 6316 10304 6332 10368
rect 6396 10304 6404 10368
rect 6084 9280 6404 10304
rect 6084 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6332 9280
rect 6396 9216 6404 9280
rect 6084 8192 6404 9216
rect 6084 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6332 8192
rect 6396 8128 6404 8192
rect 6084 7104 6404 8128
rect 6084 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6332 7104
rect 6396 7040 6404 7104
rect 6084 6016 6404 7040
rect 6084 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6332 6016
rect 6396 5952 6404 6016
rect 6084 4928 6404 5952
rect 6084 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6332 4928
rect 6396 4864 6404 4928
rect 6084 3840 6404 4864
rect 6084 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6332 3840
rect 6396 3776 6404 3840
rect 6084 2752 6404 3776
rect 6084 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6332 2752
rect 6396 2688 6404 2752
rect 5763 2684 5829 2685
rect 5763 2620 5764 2684
rect 5828 2620 5829 2684
rect 5763 2619 5829 2620
rect 5395 1868 5461 1869
rect 5395 1804 5396 1868
rect 5460 1804 5461 1868
rect 5395 1803 5461 1804
rect 4370 1056 4378 1120
rect 4442 1056 4458 1120
rect 4522 1056 4538 1120
rect 4602 1056 4618 1120
rect 4682 1056 4690 1120
rect 4370 1040 4690 1056
rect 6084 1664 6404 2688
rect 6686 2685 6746 41787
rect 7235 20364 7301 20365
rect 7235 20300 7236 20364
rect 7300 20300 7301 20364
rect 7235 20299 7301 20300
rect 7238 11797 7298 20299
rect 7235 11796 7301 11797
rect 7235 11732 7236 11796
rect 7300 11732 7301 11796
rect 7235 11731 7301 11732
rect 7422 2685 7482 41787
rect 7797 41376 8117 42400
rect 7797 41312 7805 41376
rect 7869 41312 7885 41376
rect 7949 41312 7965 41376
rect 8029 41312 8045 41376
rect 8109 41312 8117 41376
rect 7797 40288 8117 41312
rect 7797 40224 7805 40288
rect 7869 40224 7885 40288
rect 7949 40224 7965 40288
rect 8029 40224 8045 40288
rect 8109 40224 8117 40288
rect 7797 39200 8117 40224
rect 7797 39136 7805 39200
rect 7869 39136 7885 39200
rect 7949 39136 7965 39200
rect 8029 39136 8045 39200
rect 8109 39136 8117 39200
rect 7797 38112 8117 39136
rect 7797 38048 7805 38112
rect 7869 38048 7885 38112
rect 7949 38048 7965 38112
rect 8029 38048 8045 38112
rect 8109 38048 8117 38112
rect 7797 37024 8117 38048
rect 7797 36960 7805 37024
rect 7869 36960 7885 37024
rect 7949 36960 7965 37024
rect 8029 36960 8045 37024
rect 8109 36960 8117 37024
rect 7797 35936 8117 36960
rect 7797 35872 7805 35936
rect 7869 35872 7885 35936
rect 7949 35872 7965 35936
rect 8029 35872 8045 35936
rect 8109 35872 8117 35936
rect 7797 34848 8117 35872
rect 7797 34784 7805 34848
rect 7869 34784 7885 34848
rect 7949 34784 7965 34848
rect 8029 34784 8045 34848
rect 8109 34784 8117 34848
rect 7797 33760 8117 34784
rect 7797 33696 7805 33760
rect 7869 33696 7885 33760
rect 7949 33696 7965 33760
rect 8029 33696 8045 33760
rect 8109 33696 8117 33760
rect 7797 32672 8117 33696
rect 7797 32608 7805 32672
rect 7869 32608 7885 32672
rect 7949 32608 7965 32672
rect 8029 32608 8045 32672
rect 8109 32608 8117 32672
rect 7797 31584 8117 32608
rect 7797 31520 7805 31584
rect 7869 31520 7885 31584
rect 7949 31520 7965 31584
rect 8029 31520 8045 31584
rect 8109 31520 8117 31584
rect 7797 30496 8117 31520
rect 7797 30432 7805 30496
rect 7869 30432 7885 30496
rect 7949 30432 7965 30496
rect 8029 30432 8045 30496
rect 8109 30432 8117 30496
rect 7797 29408 8117 30432
rect 7797 29344 7805 29408
rect 7869 29344 7885 29408
rect 7949 29344 7965 29408
rect 8029 29344 8045 29408
rect 8109 29344 8117 29408
rect 7797 28320 8117 29344
rect 9511 43008 9831 43568
rect 9511 42944 9519 43008
rect 9583 42944 9599 43008
rect 9663 42944 9679 43008
rect 9743 42944 9759 43008
rect 9823 42944 9831 43008
rect 9511 41920 9831 42944
rect 9511 41856 9519 41920
rect 9583 41856 9599 41920
rect 9663 41856 9679 41920
rect 9743 41856 9759 41920
rect 9823 41856 9831 41920
rect 9511 40832 9831 41856
rect 11224 43552 11544 43568
rect 11224 43488 11232 43552
rect 11296 43488 11312 43552
rect 11376 43488 11392 43552
rect 11456 43488 11472 43552
rect 11536 43488 11544 43552
rect 11224 42464 11544 43488
rect 11224 42400 11232 42464
rect 11296 42400 11312 42464
rect 11376 42400 11392 42464
rect 11456 42400 11472 42464
rect 11536 42400 11544 42464
rect 10915 41852 10981 41853
rect 10915 41788 10916 41852
rect 10980 41788 10981 41852
rect 10915 41787 10981 41788
rect 10731 41580 10797 41581
rect 10731 41516 10732 41580
rect 10796 41516 10797 41580
rect 10731 41515 10797 41516
rect 9511 40768 9519 40832
rect 9583 40768 9599 40832
rect 9663 40768 9679 40832
rect 9743 40768 9759 40832
rect 9823 40768 9831 40832
rect 9511 39744 9831 40768
rect 9511 39680 9519 39744
rect 9583 39680 9599 39744
rect 9663 39680 9679 39744
rect 9743 39680 9759 39744
rect 9823 39680 9831 39744
rect 9511 38656 9831 39680
rect 9511 38592 9519 38656
rect 9583 38592 9599 38656
rect 9663 38592 9679 38656
rect 9743 38592 9759 38656
rect 9823 38592 9831 38656
rect 9511 37568 9831 38592
rect 9511 37504 9519 37568
rect 9583 37504 9599 37568
rect 9663 37504 9679 37568
rect 9743 37504 9759 37568
rect 9823 37504 9831 37568
rect 9511 36480 9831 37504
rect 9511 36416 9519 36480
rect 9583 36416 9599 36480
rect 9663 36416 9679 36480
rect 9743 36416 9759 36480
rect 9823 36416 9831 36480
rect 9511 35392 9831 36416
rect 9511 35328 9519 35392
rect 9583 35328 9599 35392
rect 9663 35328 9679 35392
rect 9743 35328 9759 35392
rect 9823 35328 9831 35392
rect 9511 34304 9831 35328
rect 9511 34240 9519 34304
rect 9583 34240 9599 34304
rect 9663 34240 9679 34304
rect 9743 34240 9759 34304
rect 9823 34240 9831 34304
rect 9511 33216 9831 34240
rect 9511 33152 9519 33216
rect 9583 33152 9599 33216
rect 9663 33152 9679 33216
rect 9743 33152 9759 33216
rect 9823 33152 9831 33216
rect 9511 32128 9831 33152
rect 9511 32064 9519 32128
rect 9583 32064 9599 32128
rect 9663 32064 9679 32128
rect 9743 32064 9759 32128
rect 9823 32064 9831 32128
rect 9511 31040 9831 32064
rect 9511 30976 9519 31040
rect 9583 30976 9599 31040
rect 9663 30976 9679 31040
rect 9743 30976 9759 31040
rect 9823 30976 9831 31040
rect 9511 29952 9831 30976
rect 9511 29888 9519 29952
rect 9583 29888 9599 29952
rect 9663 29888 9679 29952
rect 9743 29888 9759 29952
rect 9823 29888 9831 29952
rect 9075 29068 9141 29069
rect 9075 29004 9076 29068
rect 9140 29004 9141 29068
rect 9075 29003 9141 29004
rect 9259 29068 9325 29069
rect 9259 29004 9260 29068
rect 9324 29004 9325 29068
rect 9259 29003 9325 29004
rect 7797 28256 7805 28320
rect 7869 28256 7885 28320
rect 7949 28256 7965 28320
rect 8029 28256 8045 28320
rect 8109 28256 8117 28320
rect 7797 27232 8117 28256
rect 7797 27168 7805 27232
rect 7869 27168 7885 27232
rect 7949 27168 7965 27232
rect 8029 27168 8045 27232
rect 8109 27168 8117 27232
rect 7797 26144 8117 27168
rect 8891 26348 8957 26349
rect 8891 26284 8892 26348
rect 8956 26284 8957 26348
rect 8891 26283 8957 26284
rect 7797 26080 7805 26144
rect 7869 26080 7885 26144
rect 7949 26080 7965 26144
rect 8029 26080 8045 26144
rect 8109 26080 8117 26144
rect 7797 25056 8117 26080
rect 7797 24992 7805 25056
rect 7869 24992 7885 25056
rect 7949 24992 7965 25056
rect 8029 24992 8045 25056
rect 8109 24992 8117 25056
rect 7797 23968 8117 24992
rect 7797 23904 7805 23968
rect 7869 23904 7885 23968
rect 7949 23904 7965 23968
rect 8029 23904 8045 23968
rect 8109 23904 8117 23968
rect 7797 22880 8117 23904
rect 7797 22816 7805 22880
rect 7869 22816 7885 22880
rect 7949 22816 7965 22880
rect 8029 22816 8045 22880
rect 8109 22816 8117 22880
rect 7797 21792 8117 22816
rect 7797 21728 7805 21792
rect 7869 21728 7885 21792
rect 7949 21728 7965 21792
rect 8029 21728 8045 21792
rect 8109 21728 8117 21792
rect 7797 20704 8117 21728
rect 7797 20640 7805 20704
rect 7869 20640 7885 20704
rect 7949 20640 7965 20704
rect 8029 20640 8045 20704
rect 8109 20640 8117 20704
rect 7797 19616 8117 20640
rect 8707 20500 8773 20501
rect 8707 20436 8708 20500
rect 8772 20436 8773 20500
rect 8707 20435 8773 20436
rect 8710 19821 8770 20435
rect 8707 19820 8773 19821
rect 8707 19756 8708 19820
rect 8772 19756 8773 19820
rect 8707 19755 8773 19756
rect 7797 19552 7805 19616
rect 7869 19552 7885 19616
rect 7949 19552 7965 19616
rect 8029 19552 8045 19616
rect 8109 19552 8117 19616
rect 7797 18528 8117 19552
rect 7797 18464 7805 18528
rect 7869 18464 7885 18528
rect 7949 18464 7965 18528
rect 8029 18464 8045 18528
rect 8109 18464 8117 18528
rect 7797 17440 8117 18464
rect 7797 17376 7805 17440
rect 7869 17376 7885 17440
rect 7949 17376 7965 17440
rect 8029 17376 8045 17440
rect 8109 17376 8117 17440
rect 7797 16352 8117 17376
rect 7797 16288 7805 16352
rect 7869 16288 7885 16352
rect 7949 16288 7965 16352
rect 8029 16288 8045 16352
rect 8109 16288 8117 16352
rect 7797 15264 8117 16288
rect 7797 15200 7805 15264
rect 7869 15200 7885 15264
rect 7949 15200 7965 15264
rect 8029 15200 8045 15264
rect 8109 15200 8117 15264
rect 7797 14176 8117 15200
rect 7797 14112 7805 14176
rect 7869 14112 7885 14176
rect 7949 14112 7965 14176
rect 8029 14112 8045 14176
rect 8109 14112 8117 14176
rect 7797 13088 8117 14112
rect 7797 13024 7805 13088
rect 7869 13024 7885 13088
rect 7949 13024 7965 13088
rect 8029 13024 8045 13088
rect 8109 13024 8117 13088
rect 7797 12000 8117 13024
rect 7797 11936 7805 12000
rect 7869 11936 7885 12000
rect 7949 11936 7965 12000
rect 8029 11936 8045 12000
rect 8109 11936 8117 12000
rect 7797 10912 8117 11936
rect 7797 10848 7805 10912
rect 7869 10848 7885 10912
rect 7949 10848 7965 10912
rect 8029 10848 8045 10912
rect 8109 10848 8117 10912
rect 7797 9824 8117 10848
rect 7797 9760 7805 9824
rect 7869 9760 7885 9824
rect 7949 9760 7965 9824
rect 8029 9760 8045 9824
rect 8109 9760 8117 9824
rect 7797 8736 8117 9760
rect 7797 8672 7805 8736
rect 7869 8672 7885 8736
rect 7949 8672 7965 8736
rect 8029 8672 8045 8736
rect 8109 8672 8117 8736
rect 7797 7648 8117 8672
rect 7797 7584 7805 7648
rect 7869 7584 7885 7648
rect 7949 7584 7965 7648
rect 8029 7584 8045 7648
rect 8109 7584 8117 7648
rect 7797 6560 8117 7584
rect 7797 6496 7805 6560
rect 7869 6496 7885 6560
rect 7949 6496 7965 6560
rect 8029 6496 8045 6560
rect 8109 6496 8117 6560
rect 7797 5472 8117 6496
rect 7797 5408 7805 5472
rect 7869 5408 7885 5472
rect 7949 5408 7965 5472
rect 8029 5408 8045 5472
rect 8109 5408 8117 5472
rect 7797 4384 8117 5408
rect 7797 4320 7805 4384
rect 7869 4320 7885 4384
rect 7949 4320 7965 4384
rect 8029 4320 8045 4384
rect 8109 4320 8117 4384
rect 7797 3296 8117 4320
rect 8710 4045 8770 19755
rect 8894 16149 8954 26283
rect 9078 20093 9138 29003
rect 9075 20092 9141 20093
rect 9075 20028 9076 20092
rect 9140 20028 9141 20092
rect 9075 20027 9141 20028
rect 9078 19685 9138 20027
rect 9262 19957 9322 29003
rect 9511 28864 9831 29888
rect 9511 28800 9519 28864
rect 9583 28800 9599 28864
rect 9663 28800 9679 28864
rect 9743 28800 9759 28864
rect 9823 28800 9831 28864
rect 9511 27776 9831 28800
rect 9511 27712 9519 27776
rect 9583 27712 9599 27776
rect 9663 27712 9679 27776
rect 9743 27712 9759 27776
rect 9823 27712 9831 27776
rect 9511 26688 9831 27712
rect 9511 26624 9519 26688
rect 9583 26624 9599 26688
rect 9663 26624 9679 26688
rect 9743 26624 9759 26688
rect 9823 26624 9831 26688
rect 9511 25600 9831 26624
rect 9511 25536 9519 25600
rect 9583 25536 9599 25600
rect 9663 25536 9679 25600
rect 9743 25536 9759 25600
rect 9823 25536 9831 25600
rect 9511 24512 9831 25536
rect 9511 24448 9519 24512
rect 9583 24448 9599 24512
rect 9663 24448 9679 24512
rect 9743 24448 9759 24512
rect 9823 24448 9831 24512
rect 9511 23424 9831 24448
rect 9511 23360 9519 23424
rect 9583 23360 9599 23424
rect 9663 23360 9679 23424
rect 9743 23360 9759 23424
rect 9823 23360 9831 23424
rect 9511 22336 9831 23360
rect 9511 22272 9519 22336
rect 9583 22272 9599 22336
rect 9663 22272 9679 22336
rect 9743 22272 9759 22336
rect 9823 22272 9831 22336
rect 9511 21248 9831 22272
rect 9511 21184 9519 21248
rect 9583 21184 9599 21248
rect 9663 21184 9679 21248
rect 9743 21184 9759 21248
rect 9823 21184 9831 21248
rect 9511 20160 9831 21184
rect 9511 20096 9519 20160
rect 9583 20096 9599 20160
rect 9663 20096 9679 20160
rect 9743 20096 9759 20160
rect 9823 20096 9831 20160
rect 9259 19956 9325 19957
rect 9259 19892 9260 19956
rect 9324 19892 9325 19956
rect 9259 19891 9325 19892
rect 9075 19684 9141 19685
rect 9075 19620 9076 19684
rect 9140 19620 9141 19684
rect 9075 19619 9141 19620
rect 9511 19072 9831 20096
rect 10547 19276 10613 19277
rect 10547 19212 10548 19276
rect 10612 19212 10613 19276
rect 10547 19211 10613 19212
rect 9511 19008 9519 19072
rect 9583 19008 9599 19072
rect 9663 19008 9679 19072
rect 9743 19008 9759 19072
rect 9823 19008 9831 19072
rect 9511 17984 9831 19008
rect 10363 18188 10429 18189
rect 10363 18124 10364 18188
rect 10428 18124 10429 18188
rect 10363 18123 10429 18124
rect 9511 17920 9519 17984
rect 9583 17920 9599 17984
rect 9663 17920 9679 17984
rect 9743 17920 9759 17984
rect 9823 17920 9831 17984
rect 9511 16896 9831 17920
rect 9511 16832 9519 16896
rect 9583 16832 9599 16896
rect 9663 16832 9679 16896
rect 9743 16832 9759 16896
rect 9823 16832 9831 16896
rect 8891 16148 8957 16149
rect 8891 16084 8892 16148
rect 8956 16084 8957 16148
rect 8891 16083 8957 16084
rect 9511 15808 9831 16832
rect 9511 15744 9519 15808
rect 9583 15744 9599 15808
rect 9663 15744 9679 15808
rect 9743 15744 9759 15808
rect 9823 15744 9831 15808
rect 9511 14720 9831 15744
rect 9511 14656 9519 14720
rect 9583 14656 9599 14720
rect 9663 14656 9679 14720
rect 9743 14656 9759 14720
rect 9823 14656 9831 14720
rect 9511 13632 9831 14656
rect 10366 14517 10426 18123
rect 10550 16557 10610 19211
rect 10547 16556 10613 16557
rect 10547 16492 10548 16556
rect 10612 16492 10613 16556
rect 10547 16491 10613 16492
rect 10363 14516 10429 14517
rect 10363 14452 10364 14516
rect 10428 14452 10429 14516
rect 10363 14451 10429 14452
rect 9511 13568 9519 13632
rect 9583 13568 9599 13632
rect 9663 13568 9679 13632
rect 9743 13568 9759 13632
rect 9823 13568 9831 13632
rect 9511 12544 9831 13568
rect 10734 13565 10794 41515
rect 10731 13564 10797 13565
rect 10731 13500 10732 13564
rect 10796 13500 10797 13564
rect 10731 13499 10797 13500
rect 9511 12480 9519 12544
rect 9583 12480 9599 12544
rect 9663 12480 9679 12544
rect 9743 12480 9759 12544
rect 9823 12480 9831 12544
rect 9511 11456 9831 12480
rect 9511 11392 9519 11456
rect 9583 11392 9599 11456
rect 9663 11392 9679 11456
rect 9743 11392 9759 11456
rect 9823 11392 9831 11456
rect 9511 10368 9831 11392
rect 9511 10304 9519 10368
rect 9583 10304 9599 10368
rect 9663 10304 9679 10368
rect 9743 10304 9759 10368
rect 9823 10304 9831 10368
rect 9511 9280 9831 10304
rect 10731 9892 10797 9893
rect 10731 9828 10732 9892
rect 10796 9828 10797 9892
rect 10731 9827 10797 9828
rect 9511 9216 9519 9280
rect 9583 9216 9599 9280
rect 9663 9216 9679 9280
rect 9743 9216 9759 9280
rect 9823 9216 9831 9280
rect 9511 8192 9831 9216
rect 10547 9212 10613 9213
rect 10547 9148 10548 9212
rect 10612 9148 10613 9212
rect 10547 9147 10613 9148
rect 9511 8128 9519 8192
rect 9583 8128 9599 8192
rect 9663 8128 9679 8192
rect 9743 8128 9759 8192
rect 9823 8128 9831 8192
rect 9511 7104 9831 8128
rect 10550 7853 10610 9147
rect 10547 7852 10613 7853
rect 10547 7788 10548 7852
rect 10612 7788 10613 7852
rect 10547 7787 10613 7788
rect 9511 7040 9519 7104
rect 9583 7040 9599 7104
rect 9663 7040 9679 7104
rect 9743 7040 9759 7104
rect 9823 7040 9831 7104
rect 9511 6016 9831 7040
rect 9511 5952 9519 6016
rect 9583 5952 9599 6016
rect 9663 5952 9679 6016
rect 9743 5952 9759 6016
rect 9823 5952 9831 6016
rect 9511 4928 9831 5952
rect 10734 5269 10794 9827
rect 10731 5268 10797 5269
rect 10731 5204 10732 5268
rect 10796 5204 10797 5268
rect 10731 5203 10797 5204
rect 9511 4864 9519 4928
rect 9583 4864 9599 4928
rect 9663 4864 9679 4928
rect 9743 4864 9759 4928
rect 9823 4864 9831 4928
rect 8707 4044 8773 4045
rect 8707 3980 8708 4044
rect 8772 3980 8773 4044
rect 8707 3979 8773 3980
rect 7797 3232 7805 3296
rect 7869 3232 7885 3296
rect 7949 3232 7965 3296
rect 8029 3232 8045 3296
rect 8109 3232 8117 3296
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 6084 1600 6092 1664
rect 6156 1600 6172 1664
rect 6236 1600 6252 1664
rect 6316 1600 6332 1664
rect 6396 1600 6404 1664
rect 6084 1040 6404 1600
rect 7797 2208 8117 3232
rect 7797 2144 7805 2208
rect 7869 2144 7885 2208
rect 7949 2144 7965 2208
rect 8029 2144 8045 2208
rect 8109 2144 8117 2208
rect 7797 1120 8117 2144
rect 7797 1056 7805 1120
rect 7869 1056 7885 1120
rect 7949 1056 7965 1120
rect 8029 1056 8045 1120
rect 8109 1056 8117 1120
rect 7797 1040 8117 1056
rect 9511 3840 9831 4864
rect 9511 3776 9519 3840
rect 9583 3776 9599 3840
rect 9663 3776 9679 3840
rect 9743 3776 9759 3840
rect 9823 3776 9831 3840
rect 9511 2752 9831 3776
rect 9511 2688 9519 2752
rect 9583 2688 9599 2752
rect 9663 2688 9679 2752
rect 9743 2688 9759 2752
rect 9823 2688 9831 2752
rect 9511 1664 9831 2688
rect 10918 2685 10978 41787
rect 11224 41376 11544 42400
rect 11224 41312 11232 41376
rect 11296 41312 11312 41376
rect 11376 41312 11392 41376
rect 11456 41312 11472 41376
rect 11536 41312 11544 41376
rect 11224 40288 11544 41312
rect 11224 40224 11232 40288
rect 11296 40224 11312 40288
rect 11376 40224 11392 40288
rect 11456 40224 11472 40288
rect 11536 40224 11544 40288
rect 11224 39200 11544 40224
rect 11224 39136 11232 39200
rect 11296 39136 11312 39200
rect 11376 39136 11392 39200
rect 11456 39136 11472 39200
rect 11536 39136 11544 39200
rect 11224 38112 11544 39136
rect 11224 38048 11232 38112
rect 11296 38048 11312 38112
rect 11376 38048 11392 38112
rect 11456 38048 11472 38112
rect 11536 38048 11544 38112
rect 11224 37024 11544 38048
rect 11224 36960 11232 37024
rect 11296 36960 11312 37024
rect 11376 36960 11392 37024
rect 11456 36960 11472 37024
rect 11536 36960 11544 37024
rect 11224 35936 11544 36960
rect 11224 35872 11232 35936
rect 11296 35872 11312 35936
rect 11376 35872 11392 35936
rect 11456 35872 11472 35936
rect 11536 35872 11544 35936
rect 11224 34848 11544 35872
rect 11224 34784 11232 34848
rect 11296 34784 11312 34848
rect 11376 34784 11392 34848
rect 11456 34784 11472 34848
rect 11536 34784 11544 34848
rect 11224 33760 11544 34784
rect 11224 33696 11232 33760
rect 11296 33696 11312 33760
rect 11376 33696 11392 33760
rect 11456 33696 11472 33760
rect 11536 33696 11544 33760
rect 11224 32672 11544 33696
rect 11224 32608 11232 32672
rect 11296 32608 11312 32672
rect 11376 32608 11392 32672
rect 11456 32608 11472 32672
rect 11536 32608 11544 32672
rect 11224 31584 11544 32608
rect 12938 43008 13258 43568
rect 12938 42944 12946 43008
rect 13010 42944 13026 43008
rect 13090 42944 13106 43008
rect 13170 42944 13186 43008
rect 13250 42944 13258 43008
rect 12938 41920 13258 42944
rect 12938 41856 12946 41920
rect 13010 41856 13026 41920
rect 13090 41856 13106 41920
rect 13170 41856 13186 41920
rect 13250 41856 13258 41920
rect 12938 40832 13258 41856
rect 12938 40768 12946 40832
rect 13010 40768 13026 40832
rect 13090 40768 13106 40832
rect 13170 40768 13186 40832
rect 13250 40768 13258 40832
rect 12938 39744 13258 40768
rect 12938 39680 12946 39744
rect 13010 39680 13026 39744
rect 13090 39680 13106 39744
rect 13170 39680 13186 39744
rect 13250 39680 13258 39744
rect 12938 38656 13258 39680
rect 12938 38592 12946 38656
rect 13010 38592 13026 38656
rect 13090 38592 13106 38656
rect 13170 38592 13186 38656
rect 13250 38592 13258 38656
rect 12938 37568 13258 38592
rect 12938 37504 12946 37568
rect 13010 37504 13026 37568
rect 13090 37504 13106 37568
rect 13170 37504 13186 37568
rect 13250 37504 13258 37568
rect 12938 36480 13258 37504
rect 12938 36416 12946 36480
rect 13010 36416 13026 36480
rect 13090 36416 13106 36480
rect 13170 36416 13186 36480
rect 13250 36416 13258 36480
rect 12938 35392 13258 36416
rect 12938 35328 12946 35392
rect 13010 35328 13026 35392
rect 13090 35328 13106 35392
rect 13170 35328 13186 35392
rect 13250 35328 13258 35392
rect 12938 34304 13258 35328
rect 12938 34240 12946 34304
rect 13010 34240 13026 34304
rect 13090 34240 13106 34304
rect 13170 34240 13186 34304
rect 13250 34240 13258 34304
rect 12938 33216 13258 34240
rect 12938 33152 12946 33216
rect 13010 33152 13026 33216
rect 13090 33152 13106 33216
rect 13170 33152 13186 33216
rect 13250 33152 13258 33216
rect 12019 32468 12085 32469
rect 12019 32404 12020 32468
rect 12084 32404 12085 32468
rect 12019 32403 12085 32404
rect 11835 32332 11901 32333
rect 11835 32268 11836 32332
rect 11900 32268 11901 32332
rect 11835 32267 11901 32268
rect 11224 31520 11232 31584
rect 11296 31520 11312 31584
rect 11376 31520 11392 31584
rect 11456 31520 11472 31584
rect 11536 31520 11544 31584
rect 11224 30496 11544 31520
rect 11224 30432 11232 30496
rect 11296 30432 11312 30496
rect 11376 30432 11392 30496
rect 11456 30432 11472 30496
rect 11536 30432 11544 30496
rect 11224 29408 11544 30432
rect 11224 29344 11232 29408
rect 11296 29344 11312 29408
rect 11376 29344 11392 29408
rect 11456 29344 11472 29408
rect 11536 29344 11544 29408
rect 11224 28320 11544 29344
rect 11224 28256 11232 28320
rect 11296 28256 11312 28320
rect 11376 28256 11392 28320
rect 11456 28256 11472 28320
rect 11536 28256 11544 28320
rect 11224 27232 11544 28256
rect 11224 27168 11232 27232
rect 11296 27168 11312 27232
rect 11376 27168 11392 27232
rect 11456 27168 11472 27232
rect 11536 27168 11544 27232
rect 11224 26144 11544 27168
rect 11224 26080 11232 26144
rect 11296 26080 11312 26144
rect 11376 26080 11392 26144
rect 11456 26080 11472 26144
rect 11536 26080 11544 26144
rect 11224 25056 11544 26080
rect 11224 24992 11232 25056
rect 11296 24992 11312 25056
rect 11376 24992 11392 25056
rect 11456 24992 11472 25056
rect 11536 24992 11544 25056
rect 11224 23968 11544 24992
rect 11224 23904 11232 23968
rect 11296 23904 11312 23968
rect 11376 23904 11392 23968
rect 11456 23904 11472 23968
rect 11536 23904 11544 23968
rect 11224 22880 11544 23904
rect 11224 22816 11232 22880
rect 11296 22816 11312 22880
rect 11376 22816 11392 22880
rect 11456 22816 11472 22880
rect 11536 22816 11544 22880
rect 11224 21792 11544 22816
rect 11838 21997 11898 32267
rect 12022 28933 12082 32403
rect 12938 32128 13258 33152
rect 12938 32064 12946 32128
rect 13010 32064 13026 32128
rect 13090 32064 13106 32128
rect 13170 32064 13186 32128
rect 13250 32064 13258 32128
rect 12571 31788 12637 31789
rect 12571 31724 12572 31788
rect 12636 31724 12637 31788
rect 12571 31723 12637 31724
rect 12019 28932 12085 28933
rect 12019 28868 12020 28932
rect 12084 28868 12085 28932
rect 12019 28867 12085 28868
rect 12574 21997 12634 31723
rect 12938 31040 13258 32064
rect 12938 30976 12946 31040
rect 13010 30976 13026 31040
rect 13090 30976 13106 31040
rect 13170 30976 13186 31040
rect 13250 30976 13258 31040
rect 12938 29952 13258 30976
rect 12938 29888 12946 29952
rect 13010 29888 13026 29952
rect 13090 29888 13106 29952
rect 13170 29888 13186 29952
rect 13250 29888 13258 29952
rect 12938 28864 13258 29888
rect 12938 28800 12946 28864
rect 13010 28800 13026 28864
rect 13090 28800 13106 28864
rect 13170 28800 13186 28864
rect 13250 28800 13258 28864
rect 12938 27776 13258 28800
rect 12938 27712 12946 27776
rect 13010 27712 13026 27776
rect 13090 27712 13106 27776
rect 13170 27712 13186 27776
rect 13250 27712 13258 27776
rect 12938 26688 13258 27712
rect 12938 26624 12946 26688
rect 13010 26624 13026 26688
rect 13090 26624 13106 26688
rect 13170 26624 13186 26688
rect 13250 26624 13258 26688
rect 12938 25600 13258 26624
rect 12938 25536 12946 25600
rect 13010 25536 13026 25600
rect 13090 25536 13106 25600
rect 13170 25536 13186 25600
rect 13250 25536 13258 25600
rect 12938 24512 13258 25536
rect 12938 24448 12946 24512
rect 13010 24448 13026 24512
rect 13090 24448 13106 24512
rect 13170 24448 13186 24512
rect 13250 24448 13258 24512
rect 12938 23424 13258 24448
rect 14651 43552 14971 43568
rect 14651 43488 14659 43552
rect 14723 43488 14739 43552
rect 14803 43488 14819 43552
rect 14883 43488 14899 43552
rect 14963 43488 14971 43552
rect 14651 42464 14971 43488
rect 14651 42400 14659 42464
rect 14723 42400 14739 42464
rect 14803 42400 14819 42464
rect 14883 42400 14899 42464
rect 14963 42400 14971 42464
rect 14651 41376 14971 42400
rect 14651 41312 14659 41376
rect 14723 41312 14739 41376
rect 14803 41312 14819 41376
rect 14883 41312 14899 41376
rect 14963 41312 14971 41376
rect 14651 40288 14971 41312
rect 14651 40224 14659 40288
rect 14723 40224 14739 40288
rect 14803 40224 14819 40288
rect 14883 40224 14899 40288
rect 14963 40224 14971 40288
rect 14651 39200 14971 40224
rect 14651 39136 14659 39200
rect 14723 39136 14739 39200
rect 14803 39136 14819 39200
rect 14883 39136 14899 39200
rect 14963 39136 14971 39200
rect 14651 38112 14971 39136
rect 14651 38048 14659 38112
rect 14723 38048 14739 38112
rect 14803 38048 14819 38112
rect 14883 38048 14899 38112
rect 14963 38048 14971 38112
rect 14651 37024 14971 38048
rect 14651 36960 14659 37024
rect 14723 36960 14739 37024
rect 14803 36960 14819 37024
rect 14883 36960 14899 37024
rect 14963 36960 14971 37024
rect 14651 35936 14971 36960
rect 14651 35872 14659 35936
rect 14723 35872 14739 35936
rect 14803 35872 14819 35936
rect 14883 35872 14899 35936
rect 14963 35872 14971 35936
rect 14651 34848 14971 35872
rect 14651 34784 14659 34848
rect 14723 34784 14739 34848
rect 14803 34784 14819 34848
rect 14883 34784 14899 34848
rect 14963 34784 14971 34848
rect 14651 33760 14971 34784
rect 14651 33696 14659 33760
rect 14723 33696 14739 33760
rect 14803 33696 14819 33760
rect 14883 33696 14899 33760
rect 14963 33696 14971 33760
rect 14651 32672 14971 33696
rect 14651 32608 14659 32672
rect 14723 32608 14739 32672
rect 14803 32608 14819 32672
rect 14883 32608 14899 32672
rect 14963 32608 14971 32672
rect 14651 31584 14971 32608
rect 14651 31520 14659 31584
rect 14723 31520 14739 31584
rect 14803 31520 14819 31584
rect 14883 31520 14899 31584
rect 14963 31520 14971 31584
rect 14651 30496 14971 31520
rect 14651 30432 14659 30496
rect 14723 30432 14739 30496
rect 14803 30432 14819 30496
rect 14883 30432 14899 30496
rect 14963 30432 14971 30496
rect 14651 29408 14971 30432
rect 14651 29344 14659 29408
rect 14723 29344 14739 29408
rect 14803 29344 14819 29408
rect 14883 29344 14899 29408
rect 14963 29344 14971 29408
rect 14651 28320 14971 29344
rect 14651 28256 14659 28320
rect 14723 28256 14739 28320
rect 14803 28256 14819 28320
rect 14883 28256 14899 28320
rect 14963 28256 14971 28320
rect 14651 27232 14971 28256
rect 14651 27168 14659 27232
rect 14723 27168 14739 27232
rect 14803 27168 14819 27232
rect 14883 27168 14899 27232
rect 14963 27168 14971 27232
rect 14651 26144 14971 27168
rect 14651 26080 14659 26144
rect 14723 26080 14739 26144
rect 14803 26080 14819 26144
rect 14883 26080 14899 26144
rect 14963 26080 14971 26144
rect 14651 25056 14971 26080
rect 14651 24992 14659 25056
rect 14723 24992 14739 25056
rect 14803 24992 14819 25056
rect 14883 24992 14899 25056
rect 14963 24992 14971 25056
rect 14651 23968 14971 24992
rect 14651 23904 14659 23968
rect 14723 23904 14739 23968
rect 14803 23904 14819 23968
rect 14883 23904 14899 23968
rect 14963 23904 14971 23968
rect 13491 23900 13557 23901
rect 13491 23836 13492 23900
rect 13556 23836 13557 23900
rect 13491 23835 13557 23836
rect 12938 23360 12946 23424
rect 13010 23360 13026 23424
rect 13090 23360 13106 23424
rect 13170 23360 13186 23424
rect 13250 23360 13258 23424
rect 12938 22336 13258 23360
rect 12938 22272 12946 22336
rect 13010 22272 13026 22336
rect 13090 22272 13106 22336
rect 13170 22272 13186 22336
rect 13250 22272 13258 22336
rect 11835 21996 11901 21997
rect 11835 21932 11836 21996
rect 11900 21932 11901 21996
rect 11835 21931 11901 21932
rect 12571 21996 12637 21997
rect 12571 21932 12572 21996
rect 12636 21932 12637 21996
rect 12571 21931 12637 21932
rect 11224 21728 11232 21792
rect 11296 21728 11312 21792
rect 11376 21728 11392 21792
rect 11456 21728 11472 21792
rect 11536 21728 11544 21792
rect 11224 20704 11544 21728
rect 11224 20640 11232 20704
rect 11296 20640 11312 20704
rect 11376 20640 11392 20704
rect 11456 20640 11472 20704
rect 11536 20640 11544 20704
rect 11224 19616 11544 20640
rect 11224 19552 11232 19616
rect 11296 19552 11312 19616
rect 11376 19552 11392 19616
rect 11456 19552 11472 19616
rect 11536 19552 11544 19616
rect 11224 18528 11544 19552
rect 11224 18464 11232 18528
rect 11296 18464 11312 18528
rect 11376 18464 11392 18528
rect 11456 18464 11472 18528
rect 11536 18464 11544 18528
rect 11224 17440 11544 18464
rect 11838 17917 11898 21931
rect 11835 17916 11901 17917
rect 11835 17852 11836 17916
rect 11900 17852 11901 17916
rect 11835 17851 11901 17852
rect 11224 17376 11232 17440
rect 11296 17376 11312 17440
rect 11376 17376 11392 17440
rect 11456 17376 11472 17440
rect 11536 17376 11544 17440
rect 11224 16352 11544 17376
rect 11224 16288 11232 16352
rect 11296 16288 11312 16352
rect 11376 16288 11392 16352
rect 11456 16288 11472 16352
rect 11536 16288 11544 16352
rect 11224 15264 11544 16288
rect 12574 15877 12634 21931
rect 12938 21248 13258 22272
rect 12938 21184 12946 21248
rect 13010 21184 13026 21248
rect 13090 21184 13106 21248
rect 13170 21184 13186 21248
rect 13250 21184 13258 21248
rect 12755 20772 12821 20773
rect 12755 20708 12756 20772
rect 12820 20708 12821 20772
rect 12755 20707 12821 20708
rect 12758 16149 12818 20707
rect 12938 20160 13258 21184
rect 13494 21181 13554 23835
rect 14651 22880 14971 23904
rect 14651 22816 14659 22880
rect 14723 22816 14739 22880
rect 14803 22816 14819 22880
rect 14883 22816 14899 22880
rect 14963 22816 14971 22880
rect 13859 22404 13925 22405
rect 13859 22340 13860 22404
rect 13924 22340 13925 22404
rect 13859 22339 13925 22340
rect 13491 21180 13557 21181
rect 13491 21116 13492 21180
rect 13556 21116 13557 21180
rect 13491 21115 13557 21116
rect 12938 20096 12946 20160
rect 13010 20096 13026 20160
rect 13090 20096 13106 20160
rect 13170 20096 13186 20160
rect 13250 20096 13258 20160
rect 12938 19072 13258 20096
rect 12938 19008 12946 19072
rect 13010 19008 13026 19072
rect 13090 19008 13106 19072
rect 13170 19008 13186 19072
rect 13250 19008 13258 19072
rect 12938 17984 13258 19008
rect 13491 18188 13557 18189
rect 13491 18124 13492 18188
rect 13556 18124 13557 18188
rect 13491 18123 13557 18124
rect 12938 17920 12946 17984
rect 13010 17920 13026 17984
rect 13090 17920 13106 17984
rect 13170 17920 13186 17984
rect 13250 17920 13258 17984
rect 12938 16896 13258 17920
rect 12938 16832 12946 16896
rect 13010 16832 13026 16896
rect 13090 16832 13106 16896
rect 13170 16832 13186 16896
rect 13250 16832 13258 16896
rect 12755 16148 12821 16149
rect 12755 16084 12756 16148
rect 12820 16084 12821 16148
rect 12755 16083 12821 16084
rect 12571 15876 12637 15877
rect 12571 15812 12572 15876
rect 12636 15812 12637 15876
rect 12571 15811 12637 15812
rect 12938 15808 13258 16832
rect 13494 16285 13554 18123
rect 13862 17237 13922 22339
rect 14651 21792 14971 22816
rect 15331 21996 15397 21997
rect 15331 21932 15332 21996
rect 15396 21932 15397 21996
rect 15331 21931 15397 21932
rect 14651 21728 14659 21792
rect 14723 21728 14739 21792
rect 14803 21728 14819 21792
rect 14883 21728 14899 21792
rect 14963 21728 14971 21792
rect 14651 20704 14971 21728
rect 14651 20640 14659 20704
rect 14723 20640 14739 20704
rect 14803 20640 14819 20704
rect 14883 20640 14899 20704
rect 14963 20640 14971 20704
rect 14651 19616 14971 20640
rect 14651 19552 14659 19616
rect 14723 19552 14739 19616
rect 14803 19552 14819 19616
rect 14883 19552 14899 19616
rect 14963 19552 14971 19616
rect 14651 18528 14971 19552
rect 14651 18464 14659 18528
rect 14723 18464 14739 18528
rect 14803 18464 14819 18528
rect 14883 18464 14899 18528
rect 14963 18464 14971 18528
rect 14651 17440 14971 18464
rect 14651 17376 14659 17440
rect 14723 17376 14739 17440
rect 14803 17376 14819 17440
rect 14883 17376 14899 17440
rect 14963 17376 14971 17440
rect 13859 17236 13925 17237
rect 13859 17172 13860 17236
rect 13924 17172 13925 17236
rect 13859 17171 13925 17172
rect 14651 16352 14971 17376
rect 14651 16288 14659 16352
rect 14723 16288 14739 16352
rect 14803 16288 14819 16352
rect 14883 16288 14899 16352
rect 14963 16288 14971 16352
rect 13491 16284 13557 16285
rect 13491 16220 13492 16284
rect 13556 16220 13557 16284
rect 13491 16219 13557 16220
rect 13859 16284 13925 16285
rect 13859 16220 13860 16284
rect 13924 16220 13925 16284
rect 13859 16219 13925 16220
rect 12938 15744 12946 15808
rect 13010 15744 13026 15808
rect 13090 15744 13106 15808
rect 13170 15744 13186 15808
rect 13250 15744 13258 15808
rect 11651 15604 11717 15605
rect 11651 15540 11652 15604
rect 11716 15540 11717 15604
rect 11651 15539 11717 15540
rect 11224 15200 11232 15264
rect 11296 15200 11312 15264
rect 11376 15200 11392 15264
rect 11456 15200 11472 15264
rect 11536 15200 11544 15264
rect 11224 14176 11544 15200
rect 11224 14112 11232 14176
rect 11296 14112 11312 14176
rect 11376 14112 11392 14176
rect 11456 14112 11472 14176
rect 11536 14112 11544 14176
rect 11224 13088 11544 14112
rect 11224 13024 11232 13088
rect 11296 13024 11312 13088
rect 11376 13024 11392 13088
rect 11456 13024 11472 13088
rect 11536 13024 11544 13088
rect 11224 12000 11544 13024
rect 11654 12341 11714 15539
rect 12938 14720 13258 15744
rect 12938 14656 12946 14720
rect 13010 14656 13026 14720
rect 13090 14656 13106 14720
rect 13170 14656 13186 14720
rect 13250 14656 13258 14720
rect 12938 13632 13258 14656
rect 13675 13836 13741 13837
rect 13675 13772 13676 13836
rect 13740 13772 13741 13836
rect 13675 13771 13741 13772
rect 12938 13568 12946 13632
rect 13010 13568 13026 13632
rect 13090 13568 13106 13632
rect 13170 13568 13186 13632
rect 13250 13568 13258 13632
rect 11835 13564 11901 13565
rect 11835 13500 11836 13564
rect 11900 13500 11901 13564
rect 11835 13499 11901 13500
rect 11651 12340 11717 12341
rect 11651 12276 11652 12340
rect 11716 12276 11717 12340
rect 11651 12275 11717 12276
rect 11224 11936 11232 12000
rect 11296 11936 11312 12000
rect 11376 11936 11392 12000
rect 11456 11936 11472 12000
rect 11536 11936 11544 12000
rect 11224 10912 11544 11936
rect 11224 10848 11232 10912
rect 11296 10848 11312 10912
rect 11376 10848 11392 10912
rect 11456 10848 11472 10912
rect 11536 10848 11544 10912
rect 11224 9824 11544 10848
rect 11224 9760 11232 9824
rect 11296 9760 11312 9824
rect 11376 9760 11392 9824
rect 11456 9760 11472 9824
rect 11536 9760 11544 9824
rect 11224 8736 11544 9760
rect 11651 9348 11717 9349
rect 11651 9284 11652 9348
rect 11716 9284 11717 9348
rect 11651 9283 11717 9284
rect 11224 8672 11232 8736
rect 11296 8672 11312 8736
rect 11376 8672 11392 8736
rect 11456 8672 11472 8736
rect 11536 8672 11544 8736
rect 11224 7648 11544 8672
rect 11224 7584 11232 7648
rect 11296 7584 11312 7648
rect 11376 7584 11392 7648
rect 11456 7584 11472 7648
rect 11536 7584 11544 7648
rect 11224 6560 11544 7584
rect 11224 6496 11232 6560
rect 11296 6496 11312 6560
rect 11376 6496 11392 6560
rect 11456 6496 11472 6560
rect 11536 6496 11544 6560
rect 11224 5472 11544 6496
rect 11654 5949 11714 9283
rect 11838 8805 11898 13499
rect 12571 12612 12637 12613
rect 12571 12548 12572 12612
rect 12636 12548 12637 12612
rect 12571 12547 12637 12548
rect 12203 10436 12269 10437
rect 12203 10372 12204 10436
rect 12268 10372 12269 10436
rect 12203 10371 12269 10372
rect 12206 9485 12266 10371
rect 12203 9484 12269 9485
rect 12203 9420 12204 9484
rect 12268 9420 12269 9484
rect 12203 9419 12269 9420
rect 12203 9348 12269 9349
rect 12203 9284 12204 9348
rect 12268 9284 12269 9348
rect 12203 9283 12269 9284
rect 11835 8804 11901 8805
rect 11835 8740 11836 8804
rect 11900 8740 11901 8804
rect 11835 8739 11901 8740
rect 12206 8669 12266 9283
rect 12203 8668 12269 8669
rect 12203 8604 12204 8668
rect 12268 8604 12269 8668
rect 12203 8603 12269 8604
rect 12574 7853 12634 12547
rect 12938 12544 13258 13568
rect 12938 12480 12946 12544
rect 13010 12480 13026 12544
rect 13090 12480 13106 12544
rect 13170 12480 13186 12544
rect 13250 12480 13258 12544
rect 12755 12476 12821 12477
rect 12755 12412 12756 12476
rect 12820 12412 12821 12476
rect 12755 12411 12821 12412
rect 12758 9213 12818 12411
rect 12938 11456 13258 12480
rect 12938 11392 12946 11456
rect 13010 11392 13026 11456
rect 13090 11392 13106 11456
rect 13170 11392 13186 11456
rect 13250 11392 13258 11456
rect 12938 10368 13258 11392
rect 12938 10304 12946 10368
rect 13010 10304 13026 10368
rect 13090 10304 13106 10368
rect 13170 10304 13186 10368
rect 13250 10304 13258 10368
rect 12938 9280 13258 10304
rect 12938 9216 12946 9280
rect 13010 9216 13026 9280
rect 13090 9216 13106 9280
rect 13170 9216 13186 9280
rect 13250 9216 13258 9280
rect 12755 9212 12821 9213
rect 12755 9148 12756 9212
rect 12820 9148 12821 9212
rect 12755 9147 12821 9148
rect 12938 8192 13258 9216
rect 13678 8261 13738 13771
rect 13862 12477 13922 16219
rect 14651 15264 14971 16288
rect 14651 15200 14659 15264
rect 14723 15200 14739 15264
rect 14803 15200 14819 15264
rect 14883 15200 14899 15264
rect 14963 15200 14971 15264
rect 14651 14176 14971 15200
rect 14651 14112 14659 14176
rect 14723 14112 14739 14176
rect 14803 14112 14819 14176
rect 14883 14112 14899 14176
rect 14963 14112 14971 14176
rect 14651 13088 14971 14112
rect 15334 13565 15394 21931
rect 15331 13564 15397 13565
rect 15331 13500 15332 13564
rect 15396 13500 15397 13564
rect 15331 13499 15397 13500
rect 14651 13024 14659 13088
rect 14723 13024 14739 13088
rect 14803 13024 14819 13088
rect 14883 13024 14899 13088
rect 14963 13024 14971 13088
rect 13859 12476 13925 12477
rect 13859 12412 13860 12476
rect 13924 12412 13925 12476
rect 13859 12411 13925 12412
rect 14651 12000 14971 13024
rect 14651 11936 14659 12000
rect 14723 11936 14739 12000
rect 14803 11936 14819 12000
rect 14883 11936 14899 12000
rect 14963 11936 14971 12000
rect 14651 10912 14971 11936
rect 14651 10848 14659 10912
rect 14723 10848 14739 10912
rect 14803 10848 14819 10912
rect 14883 10848 14899 10912
rect 14963 10848 14971 10912
rect 14651 9824 14971 10848
rect 14651 9760 14659 9824
rect 14723 9760 14739 9824
rect 14803 9760 14819 9824
rect 14883 9760 14899 9824
rect 14963 9760 14971 9824
rect 14651 8736 14971 9760
rect 14651 8672 14659 8736
rect 14723 8672 14739 8736
rect 14803 8672 14819 8736
rect 14883 8672 14899 8736
rect 14963 8672 14971 8736
rect 13675 8260 13741 8261
rect 13675 8196 13676 8260
rect 13740 8196 13741 8260
rect 13675 8195 13741 8196
rect 12938 8128 12946 8192
rect 13010 8128 13026 8192
rect 13090 8128 13106 8192
rect 13170 8128 13186 8192
rect 13250 8128 13258 8192
rect 12571 7852 12637 7853
rect 12571 7788 12572 7852
rect 12636 7788 12637 7852
rect 12571 7787 12637 7788
rect 12574 6085 12634 7787
rect 12938 7104 13258 8128
rect 12938 7040 12946 7104
rect 13010 7040 13026 7104
rect 13090 7040 13106 7104
rect 13170 7040 13186 7104
rect 13250 7040 13258 7104
rect 12571 6084 12637 6085
rect 12571 6020 12572 6084
rect 12636 6020 12637 6084
rect 12571 6019 12637 6020
rect 12938 6016 13258 7040
rect 12938 5952 12946 6016
rect 13010 5952 13026 6016
rect 13090 5952 13106 6016
rect 13170 5952 13186 6016
rect 13250 5952 13258 6016
rect 11651 5948 11717 5949
rect 11651 5884 11652 5948
rect 11716 5884 11717 5948
rect 11651 5883 11717 5884
rect 11224 5408 11232 5472
rect 11296 5408 11312 5472
rect 11376 5408 11392 5472
rect 11456 5408 11472 5472
rect 11536 5408 11544 5472
rect 11224 4384 11544 5408
rect 11224 4320 11232 4384
rect 11296 4320 11312 4384
rect 11376 4320 11392 4384
rect 11456 4320 11472 4384
rect 11536 4320 11544 4384
rect 11224 3296 11544 4320
rect 11224 3232 11232 3296
rect 11296 3232 11312 3296
rect 11376 3232 11392 3296
rect 11456 3232 11472 3296
rect 11536 3232 11544 3296
rect 10915 2684 10981 2685
rect 10915 2620 10916 2684
rect 10980 2620 10981 2684
rect 10915 2619 10981 2620
rect 9511 1600 9519 1664
rect 9583 1600 9599 1664
rect 9663 1600 9679 1664
rect 9743 1600 9759 1664
rect 9823 1600 9831 1664
rect 9511 1040 9831 1600
rect 11224 2208 11544 3232
rect 11224 2144 11232 2208
rect 11296 2144 11312 2208
rect 11376 2144 11392 2208
rect 11456 2144 11472 2208
rect 11536 2144 11544 2208
rect 11224 1120 11544 2144
rect 11224 1056 11232 1120
rect 11296 1056 11312 1120
rect 11376 1056 11392 1120
rect 11456 1056 11472 1120
rect 11536 1056 11544 1120
rect 11224 1040 11544 1056
rect 12938 4928 13258 5952
rect 12938 4864 12946 4928
rect 13010 4864 13026 4928
rect 13090 4864 13106 4928
rect 13170 4864 13186 4928
rect 13250 4864 13258 4928
rect 12938 3840 13258 4864
rect 12938 3776 12946 3840
rect 13010 3776 13026 3840
rect 13090 3776 13106 3840
rect 13170 3776 13186 3840
rect 13250 3776 13258 3840
rect 12938 2752 13258 3776
rect 12938 2688 12946 2752
rect 13010 2688 13026 2752
rect 13090 2688 13106 2752
rect 13170 2688 13186 2752
rect 13250 2688 13258 2752
rect 12938 1664 13258 2688
rect 12938 1600 12946 1664
rect 13010 1600 13026 1664
rect 13090 1600 13106 1664
rect 13170 1600 13186 1664
rect 13250 1600 13258 1664
rect 12938 1040 13258 1600
rect 14651 7648 14971 8672
rect 14651 7584 14659 7648
rect 14723 7584 14739 7648
rect 14803 7584 14819 7648
rect 14883 7584 14899 7648
rect 14963 7584 14971 7648
rect 14651 6560 14971 7584
rect 14651 6496 14659 6560
rect 14723 6496 14739 6560
rect 14803 6496 14819 6560
rect 14883 6496 14899 6560
rect 14963 6496 14971 6560
rect 14651 5472 14971 6496
rect 14651 5408 14659 5472
rect 14723 5408 14739 5472
rect 14803 5408 14819 5472
rect 14883 5408 14899 5472
rect 14963 5408 14971 5472
rect 14651 4384 14971 5408
rect 14651 4320 14659 4384
rect 14723 4320 14739 4384
rect 14803 4320 14819 4384
rect 14883 4320 14899 4384
rect 14963 4320 14971 4384
rect 14651 3296 14971 4320
rect 14651 3232 14659 3296
rect 14723 3232 14739 3296
rect 14803 3232 14819 3296
rect 14883 3232 14899 3296
rect 14963 3232 14971 3296
rect 14651 2208 14971 3232
rect 14651 2144 14659 2208
rect 14723 2144 14739 2208
rect 14803 2144 14819 2208
rect 14883 2144 14899 2208
rect 14963 2144 14971 2208
rect 14651 1120 14971 2144
rect 14651 1056 14659 1120
rect 14723 1056 14739 1120
rect 14803 1056 14819 1120
rect 14883 1056 14899 1120
rect 14963 1056 14971 1120
rect 14651 1040 14971 1056
use sky130_fd_sc_hd__clkbuf_1  _00_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _01_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _02_
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1688980957
transform 1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1688980957
transform 1 0 13156 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1688980957
transform 1 0 11776 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1688980957
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1688980957
transform 1 0 12328 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1688980957
transform 1 0 11960 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1688980957
transform 1 0 12144 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1688980957
transform 1 0 9844 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _16_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1688980957
transform 1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1688980957
transform 1 0 13248 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1688980957
transform 1 0 13524 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1688980957
transform 1 0 11868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1688980957
transform 1 0 12972 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1688980957
transform 1 0 14168 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1688980957
transform 1 0 12696 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1688980957
transform 1 0 12420 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1688980957
transform 1 0 11316 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1688980957
transform 1 0 12972 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1688980957
transform 1 0 12052 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1688980957
transform 1 0 10672 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1688980957
transform 1 0 11500 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1688980957
transform 1 0 13064 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1688980957
transform 1 0 13156 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1688980957
transform 1 0 12144 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1688980957
transform 1 0 13064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1688980957
transform 1 0 13156 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1688980957
transform 1 0 11776 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1688980957
transform 1 0 12604 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1688980957
transform 1 0 11776 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1688980957
transform 1 0 13524 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1688980957
transform 1 0 10948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1688980957
transform 1 0 12788 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1688980957
transform 1 0 12144 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1688980957
transform 1 0 11868 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1688980957
transform 1 0 11684 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1688980957
transform 1 0 13156 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1688980957
transform 1 0 10948 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1688980957
transform 1 0 13156 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1688980957
transform 1 0 10948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1688980957
transform 1 0 9292 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1688980957
transform 1 0 10488 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1688980957
transform 1 0 11960 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1688980957
transform 1 0 12880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1688980957
transform 1 0 10212 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1688980957
transform 1 0 10488 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1688980957
transform 1 0 12144 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1688980957
transform 1 0 12328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1688980957
transform 1 0 12972 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1688980957
transform 1 0 12512 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1688980957
transform 1 0 12788 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1688980957
transform 1 0 12788 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1688980957
transform 1 0 12512 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1688980957
transform 1 0 1748 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1688980957
transform 1 0 2760 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1688980957
transform 1 0 3312 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1688980957
transform 1 0 4140 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1688980957
transform 1 0 4968 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1688980957
transform 1 0 5704 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1688980957
transform 1 0 6440 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _88_
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _89_
timestamp 1688980957
transform 1 0 7820 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _90_
timestamp 1688980957
transform 1 0 8556 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _91_
timestamp 1688980957
transform 1 0 9292 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _92_
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _93_
timestamp 1688980957
transform 1 0 10764 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _94_
timestamp 1688980957
transform 1 0 11500 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _95_
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _96_
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _97_
timestamp 1688980957
transform 1 0 14260 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _98_
timestamp 1688980957
transform 1 0 12696 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _99_
timestamp 1688980957
transform 1 0 13984 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 13340 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 11776 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 12604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 11684 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 12880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 11408 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 9568 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 9844 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 8096 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 11592 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 12052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 9016 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 12420 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 13156 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 12788 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 13156 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 12144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 9936 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 12512 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 12236 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 7360 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 8372 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 9476 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 10948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 12052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 12512 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 11132 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 12972 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 12972 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 11960 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 10856 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 12328 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 10396 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 12604 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 10212 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 10488 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 9200 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 9752 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 12512 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 9752 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 12880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 11592 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 11868 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 12328 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 10764 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 11868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 13064 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 11960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 8096 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 9200 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_38 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_42
timestamp 1688980957
transform 1 0 4968 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_46
timestamp 1688980957
transform 1 0 5336 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_50
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_62
timestamp 1688980957
transform 1 0 6808 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_66
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_70
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_74
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_78 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_94
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_98
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_102
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_106
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_118
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_122
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_126
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_23
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_31
timestamp 1688980957
transform 1 0 3956 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_45
timestamp 1688980957
transform 1 0 5244 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_53
timestamp 1688980957
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_68
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_76
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_100
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_108
timestamp 1688980957
transform 1 0 11040 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_124
timestamp 1688980957
transform 1 0 12512 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_33
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_38
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_50
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_62
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_74
timestamp 1688980957
transform 1 0 7912 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_82
timestamp 1688980957
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_145
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_117
timestamp 1688980957
transform 1 0 11868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_134
timestamp 1688980957
transform 1 0 13432 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_42
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_77
timestamp 1688980957
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_95
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_144
timestamp 1688980957
transform 1 0 14352 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_93
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_14
timestamp 1688980957
transform 1 0 2392 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_26
timestamp 1688980957
transform 1 0 3496 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_38
timestamp 1688980957
transform 1 0 4600 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_50
timestamp 1688980957
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_90
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_102
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1688980957
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_136
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_16
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_28
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_40
timestamp 1688980957
transform 1 0 4784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1688980957
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_104
timestamp 1688980957
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_119
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_138
timestamp 1688980957
transform 1 0 13800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_142
timestamp 1688980957
transform 1 0 14168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_115
timestamp 1688980957
transform 1 0 11684 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_48
timestamp 1688980957
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_95
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_89
timestamp 1688980957
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_130
timestamp 1688980957
transform 1 0 13064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_14
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_84
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_134
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_138
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_14
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_26
timestamp 1688980957
transform 1 0 3496 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_38
timestamp 1688980957
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_47
timestamp 1688980957
transform 1 0 5428 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_86
timestamp 1688980957
transform 1 0 9016 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_90
timestamp 1688980957
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_88
timestamp 1688980957
transform 1 0 9200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_12
timestamp 1688980957
transform 1 0 2208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_24
timestamp 1688980957
transform 1 0 3312 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_32
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_49
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_74
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_80
timestamp 1688980957
transform 1 0 8464 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_92
timestamp 1688980957
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_96
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_142
timestamp 1688980957
transform 1 0 14168 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_64
timestamp 1688980957
transform 1 0 6992 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_76
timestamp 1688980957
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_76
timestamp 1688980957
transform 1 0 8096 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_99
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_145
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_16
timestamp 1688980957
transform 1 0 2576 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_61
timestamp 1688980957
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1688980957
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_110
timestamp 1688980957
transform 1 0 11224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_106
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_18
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_108
timestamp 1688980957
transform 1 0 11040 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_116
timestamp 1688980957
transform 1 0 11776 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_144
timestamp 1688980957
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_19
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_72
timestamp 1688980957
transform 1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_16
timestamp 1688980957
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_73
timestamp 1688980957
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_100
timestamp 1688980957
transform 1 0 10304 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_18
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_30
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_84
timestamp 1688980957
transform 1 0 8832 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_90
timestamp 1688980957
transform 1 0 9384 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_121
timestamp 1688980957
transform 1 0 12236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_18
timestamp 1688980957
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_47
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_63
timestamp 1688980957
transform 1 0 6900 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 1688980957
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_114
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_7
timestamp 1688980957
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_19
timestamp 1688980957
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_31
timestamp 1688980957
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_7
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_63
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_80
timestamp 1688980957
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_89
timestamp 1688980957
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_113
timestamp 1688980957
transform 1 0 11500 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_7
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_31
timestamp 1688980957
transform 1 0 3956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_73
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_85
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_144
timestamp 1688980957
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_46
timestamp 1688980957
transform 1 0 5336 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_68
timestamp 1688980957
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_80
timestamp 1688980957
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_120
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_49
timestamp 1688980957
transform 1 0 5612 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_60
timestamp 1688980957
transform 1 0 6624 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_72
timestamp 1688980957
transform 1 0 7728 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_94
timestamp 1688980957
transform 1 0 9752 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_98
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_102
timestamp 1688980957
transform 1 0 10488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_128
timestamp 1688980957
transform 1 0 12880 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_138
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_92
timestamp 1688980957
transform 1 0 9568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_114
timestamp 1688980957
transform 1 0 11592 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_144
timestamp 1688980957
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_47
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_63
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_79
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_85
timestamp 1688980957
transform 1 0 8924 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_135
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_63
timestamp 1688980957
transform 1 0 6900 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_68
timestamp 1688980957
transform 1 0 7360 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_80
timestamp 1688980957
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_101
timestamp 1688980957
transform 1 0 10396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_113
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_130
timestamp 1688980957
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_7
timestamp 1688980957
transform 1 0 1748 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_19
timestamp 1688980957
transform 1 0 2852 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_31
timestamp 1688980957
transform 1 0 3956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_43
timestamp 1688980957
transform 1 0 5060 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_50
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_63
timestamp 1688980957
transform 1 0 6900 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_80
timestamp 1688980957
transform 1 0 8464 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_92
timestamp 1688980957
transform 1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_100
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_7
timestamp 1688980957
transform 1 0 1748 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_19
timestamp 1688980957
transform 1 0 2852 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_35
timestamp 1688980957
transform 1 0 4324 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_67
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_119
timestamp 1688980957
transform 1 0 12052 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_26
timestamp 1688980957
transform 1 0 3496 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_38
timestamp 1688980957
transform 1 0 4600 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_50
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_90
timestamp 1688980957
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_94
timestamp 1688980957
transform 1 0 9752 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_101
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_7
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_19
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_25
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_104
timestamp 1688980957
transform 1 0 10672 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_144
timestamp 1688980957
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_7
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_33
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_70
timestamp 1688980957
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_129
timestamp 1688980957
transform 1 0 12972 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_13
timestamp 1688980957
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_25
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_37
timestamp 1688980957
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_49
timestamp 1688980957
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_86
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_102
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_117
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_139
timestamp 1688980957
transform 1 0 13892 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_129
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_144
timestamp 1688980957
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_13
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_25
timestamp 1688980957
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_33
timestamp 1688980957
transform 1 0 4140 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_70
timestamp 1688980957
transform 1 0 7544 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_82
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_138
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_72
timestamp 1688980957
transform 1 0 7728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_90
timestamp 1688980957
transform 1 0 9384 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_96
timestamp 1688980957
transform 1 0 9936 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_7
timestamp 1688980957
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_19
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_57
timestamp 1688980957
transform 1 0 6348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_73
timestamp 1688980957
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_7
timestamp 1688980957
transform 1 0 1748 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_19
timestamp 1688980957
transform 1 0 2852 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_31
timestamp 1688980957
transform 1 0 3956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_43
timestamp 1688980957
transform 1 0 5060 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_102
timestamp 1688980957
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_69
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_100
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_108
timestamp 1688980957
transform 1 0 11040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_19
timestamp 1688980957
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_43
timestamp 1688980957
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_90
timestamp 1688980957
transform 1 0 9384 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_108
timestamp 1688980957
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_130
timestamp 1688980957
transform 1 0 13064 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_144
timestamp 1688980957
transform 1 0 14352 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_7
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_19
timestamp 1688980957
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_59
timestamp 1688980957
transform 1 0 6532 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_75
timestamp 1688980957
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_61
timestamp 1688980957
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_98
timestamp 1688980957
transform 1 0 10120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_122
timestamp 1688980957
transform 1 0 12328 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_144
timestamp 1688980957
transform 1 0 14352 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_19
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_47
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_144
timestamp 1688980957
transform 1 0 14352 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_7
timestamp 1688980957
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_19
timestamp 1688980957
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_31
timestamp 1688980957
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_43
timestamp 1688980957
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_72
timestamp 1688980957
transform 1 0 7728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_84
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_109
timestamp 1688980957
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_135
timestamp 1688980957
transform 1 0 13524 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_145
timestamp 1688980957
transform 1 0 14444 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_94
timestamp 1688980957
transform 1 0 9752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_103
timestamp 1688980957
transform 1 0 10580 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_110
timestamp 1688980957
transform 1 0 11224 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_7
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_19
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_31
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_43
timestamp 1688980957
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_65
timestamp 1688980957
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_97
timestamp 1688980957
transform 1 0 10028 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_110
timestamp 1688980957
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_131
timestamp 1688980957
transform 1 0 13156 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_144
timestamp 1688980957
transform 1 0 14352 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_7
timestamp 1688980957
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_19
timestamp 1688980957
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_61
timestamp 1688980957
transform 1 0 6716 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_78
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_145
timestamp 1688980957
transform 1 0 14444 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_128
timestamp 1688980957
transform 1 0 12880 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_7
timestamp 1688980957
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_19
timestamp 1688980957
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_100
timestamp 1688980957
transform 1 0 10304 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_130
timestamp 1688980957
transform 1 0 13064 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_145
timestamp 1688980957
transform 1 0 14444 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_7
timestamp 1688980957
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_19
timestamp 1688980957
transform 1 0 2852 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_31
timestamp 1688980957
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_43
timestamp 1688980957
transform 1 0 5060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_75
timestamp 1688980957
transform 1 0 8004 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_79
timestamp 1688980957
transform 1 0 8372 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_91
timestamp 1688980957
transform 1 0 9476 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_98
timestamp 1688980957
transform 1 0 10120 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_104
timestamp 1688980957
transform 1 0 10672 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_110
timestamp 1688980957
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_144
timestamp 1688980957
transform 1 0 14352 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_8
timestamp 1688980957
transform 1 0 1840 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_20
timestamp 1688980957
transform 1 0 2944 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_91
timestamp 1688980957
transform 1 0 9476 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_108
timestamp 1688980957
transform 1 0 11040 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_132
timestamp 1688980957
transform 1 0 13248 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_10
timestamp 1688980957
transform 1 0 2024 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_22
timestamp 1688980957
transform 1 0 3128 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_34
timestamp 1688980957
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_46
timestamp 1688980957
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_54
timestamp 1688980957
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_92
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_97
timestamp 1688980957
transform 1 0 10028 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_101
timestamp 1688980957
transform 1 0 10396 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_110
timestamp 1688980957
transform 1 0 11224 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_117
timestamp 1688980957
transform 1 0 11868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_128
timestamp 1688980957
transform 1 0 12880 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_144
timestamp 1688980957
transform 1 0 14352 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_10
timestamp 1688980957
transform 1 0 2024 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_22
timestamp 1688980957
transform 1 0 3128 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_124
timestamp 1688980957
transform 1 0 12512 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_144
timestamp 1688980957
transform 1 0 14352 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_7
timestamp 1688980957
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_19
timestamp 1688980957
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_117
timestamp 1688980957
transform 1 0 11868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_126
timestamp 1688980957
transform 1 0 12696 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_7
timestamp 1688980957
transform 1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_14
timestamp 1688980957
transform 1 0 2392 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_26
timestamp 1688980957
transform 1 0 3496 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_38
timestamp 1688980957
transform 1 0 4600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_50
timestamp 1688980957
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_99
timestamp 1688980957
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_123
timestamp 1688980957
transform 1 0 12420 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_130
timestamp 1688980957
transform 1 0 13064 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_108
timestamp 1688980957
transform 1 0 11040 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_112
timestamp 1688980957
transform 1 0 11408 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_120
timestamp 1688980957
transform 1 0 12144 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_7
timestamp 1688980957
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_19
timestamp 1688980957
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_31
timestamp 1688980957
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_43
timestamp 1688980957
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_116
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_120
timestamp 1688980957
transform 1 0 12144 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_131
timestamp 1688980957
transform 1 0 13156 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_144
timestamp 1688980957
transform 1 0 14352 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_7
timestamp 1688980957
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_19
timestamp 1688980957
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_37
timestamp 1688980957
transform 1 0 4508 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_43
timestamp 1688980957
transform 1 0 5060 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_55
timestamp 1688980957
transform 1 0 6164 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_67
timestamp 1688980957
transform 1 0 7268 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_79
timestamp 1688980957
transform 1 0 8372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_127
timestamp 1688980957
transform 1 0 12788 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_132
timestamp 1688980957
transform 1 0 13248 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_45
timestamp 1688980957
transform 1 0 5244 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_53
timestamp 1688980957
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_117
timestamp 1688980957
transform 1 0 11868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_130
timestamp 1688980957
transform 1 0 13064 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_144
timestamp 1688980957
transform 1 0 14352 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_7
timestamp 1688980957
transform 1 0 1748 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_19
timestamp 1688980957
transform 1 0 2852 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_71
timestamp 1688980957
transform 1 0 7636 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_75
timestamp 1688980957
transform 1 0 8004 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_82
timestamp 1688980957
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_94
timestamp 1688980957
transform 1 0 9752 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_118
timestamp 1688980957
transform 1 0 11960 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_7
timestamp 1688980957
transform 1 0 1748 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_19
timestamp 1688980957
transform 1 0 2852 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_31
timestamp 1688980957
transform 1 0 3956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_43
timestamp 1688980957
transform 1 0 5060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_131
timestamp 1688980957
transform 1 0 13156 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_144
timestamp 1688980957
transform 1 0 14352 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_145
timestamp 1688980957
transform 1 0 14444 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_7
timestamp 1688980957
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_19
timestamp 1688980957
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_31
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_43
timestamp 1688980957
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_145
timestamp 1688980957
transform 1 0 14444 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_22
timestamp 1688980957
transform 1 0 3128 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_9
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_13
timestamp 1688980957
transform 1 0 2300 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_22
timestamp 1688980957
transform 1 0 3128 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_34
timestamp 1688980957
transform 1 0 4232 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_46
timestamp 1688980957
transform 1 0 5336 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_60
timestamp 1688980957
transform 1 0 6624 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_64
timestamp 1688980957
transform 1 0 6992 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_68
timestamp 1688980957
transform 1 0 7360 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_77
timestamp 1688980957
transform 1 0 8188 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_85
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_92
timestamp 1688980957
transform 1 0 9568 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_101
timestamp 1688980957
transform 1 0 10396 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_108
timestamp 1688980957
transform 1 0 11040 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_116
timestamp 1688980957
transform 1 0 11776 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_120
timestamp 1688980957
transform 1 0 12144 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_124
timestamp 1688980957
transform 1 0 12512 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_131
timestamp 1688980957
transform 1 0 13156 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_135
timestamp 1688980957
transform 1 0 13524 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_9
timestamp 1688980957
transform 1 0 1932 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_13
timestamp 1688980957
transform 1 0 2300 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_17
timestamp 1688980957
transform 1 0 2668 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_21
timestamp 1688980957
transform 1 0 3036 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_36
timestamp 1688980957
transform 1 0 4416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_48
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_57
timestamp 1688980957
transform 1 0 6348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_61
timestamp 1688980957
transform 1 0 6716 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_68
timestamp 1688980957
transform 1 0 7360 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_72
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_76
timestamp 1688980957
transform 1 0 8096 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_80
timestamp 1688980957
transform 1 0 8464 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_92
timestamp 1688980957
transform 1 0 9568 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_96
timestamp 1688980957
transform 1 0 9936 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_100
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_104
timestamp 1688980957
transform 1 0 10672 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_108
timestamp 1688980957
transform 1 0 11040 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_112
timestamp 1688980957
transform 1 0 11408 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_116
timestamp 1688980957
transform 1 0 11776 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_124
timestamp 1688980957
transform 1 0 12512 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_132
timestamp 1688980957
transform 1 0 13248 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_9
timestamp 1688980957
transform 1 0 1932 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_18
timestamp 1688980957
transform 1 0 2760 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_25
timestamp 1688980957
transform 1 0 3404 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_33
timestamp 1688980957
transform 1 0 4140 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_47
timestamp 1688980957
transform 1 0 5428 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_63
timestamp 1688980957
transform 1 0 6900 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_71
timestamp 1688980957
transform 1 0 7636 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_79
timestamp 1688980957
transform 1 0 8372 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_83
timestamp 1688980957
transform 1 0 8740 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_89
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_97
timestamp 1688980957
transform 1 0 10028 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_103
timestamp 1688980957
transform 1 0 10580 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_129
timestamp 1688980957
transform 1 0 12972 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_135
timestamp 1688980957
transform 1 0 13524 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_145
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 9476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 10212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 10948 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 11684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 12420 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input46
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input47
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  input48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 5796 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 6532 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1688980957
transform 1 0 14168 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1688980957
transform 1 0 14168 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1688980957
transform 1 0 14168 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1688980957
transform 1 0 11684 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1688980957
transform 1 0 13616 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1688980957
transform 1 0 14168 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1688980957
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1688980957
transform 1 0 14168 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1688980957
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1688980957
transform 1 0 14168 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1688980957
transform 1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1688980957
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 12328 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 1688980957
transform 1 0 13432 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1688980957
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1688980957
transform 1 0 14260 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1688980957
transform 1 0 14260 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1688980957
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1688980957
transform 1 0 11868 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1688980957
transform 1 0 14260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1688980957
transform 1 0 13616 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access._0_
timestamp 1688980957
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access._1_
timestamp 1688980957
transform 1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access._2_
timestamp 1688980957
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access._3_
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_A_IO_1_bidirectional_frame_config_pass._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_A_IO_1_bidirectional_frame_config_pass._1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_IO_1_bidirectional_frame_config_pass._2_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_A_IO_1_bidirectional_frame_config_pass._3_
timestamp 1688980957
transform 1 0 4968 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access._0_
timestamp 1688980957
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access._1_
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access._2_
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access._3_
timestamp 1688980957
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_B_IO_1_bidirectional_frame_config_pass._0_
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_B_IO_1_bidirectional_frame_config_pass._1_
timestamp 1688980957
transform 1 0 4416 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_IO_1_bidirectional_frame_config_pass._2_
timestamp 1688980957
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_B_IO_1_bidirectional_frame_config_pass._3_
timestamp 1688980957
transform 1 0 5336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 8004 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 5520 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 11684 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 8648 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 9384 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 8004 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 9936 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 7268 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 11592 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 11316 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 6532 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 8464 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 8832 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 9844 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 11224 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 5520 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 6532 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 9476 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 9660 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 11592 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 9844 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 6072 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 6440 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 4232 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 10028 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 5520 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 6624 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 11684 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 11592 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 12052 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 11684 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 6808 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 9384 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 12788 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 9016 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 9936 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 10764 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 9476 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 10856 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 6900 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 7452 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 9476 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 6716 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 12052 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 10028 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 6900 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 4324 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 5888 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 5520 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 6440 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 6440 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 4692 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._2_
timestamp 1688980957
transform 1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 11316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._2_
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._3_
timestamp 1688980957
transform 1 0 5612 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._4_
timestamp 1688980957
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 5888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._2_
timestamp 1688980957
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._3_
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._4_
timestamp 1688980957
transform 1 0 6532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._2_
timestamp 1688980957
transform 1 0 10488 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._3_
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._4_
timestamp 1688980957
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10120 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG1
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG2
timestamp 1688980957
transform 1 0 8004 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG3
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG4
timestamp 1688980957
transform 1 0 12052 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG5
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG6
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEG7
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb0
timestamp 1688980957
transform 1 0 10120 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb1
timestamp 1688980957
transform 1 0 7636 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb2
timestamp 1688980957
transform 1 0 7544 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb3
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb4
timestamp 1688980957
transform 1 0 6900 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb5
timestamp 1688980957
transform 1 0 12512 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb6
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E2BEGb7
timestamp 1688980957
transform 1 0 11592 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG0
timestamp 1688980957
transform 1 0 7820 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG1
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG2
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG3
timestamp 1688980957
transform 1 0 8004 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG5
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG6
timestamp 1688980957
transform 1 0 9200 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG7
timestamp 1688980957
transform 1 0 11592 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG8
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG9
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG10
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_E6BEG11
timestamp 1688980957
transform 1 0 11592 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG0
timestamp 1688980957
transform 1 0 5612 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG1
timestamp 1688980957
transform 1 0 11960 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG2
timestamp 1688980957
transform 1 0 6900 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG3
timestamp 1688980957
transform 1 0 9752 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG4
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG5
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG6
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG7
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG8
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG9
timestamp 1688980957
transform 1 0 6624 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG10
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG11
timestamp 1688980957
transform 1 0 11868 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG12
timestamp 1688980957
transform 1 0 6808 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG13
timestamp 1688980957
transform 1 0 11684 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG14
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix.inst_cus_mux41_buf_EE4BEG15
timestamp 1688980957
transform 1 0 12144 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1_216 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1_218
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 5060 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1_217
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1_219
timestamp 1688980957
transform 1 0 8188 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 10856 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9752 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 8740 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 9384 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  output103 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 1748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 2300 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 1564 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 1564 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 12880 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 13800 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 13248 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 13248 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 13432 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1688980957
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 13984 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1688980957
transform 1 0 14168 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1688980957
transform 1 0 13064 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1688980957
transform 1 0 14168 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1688980957
transform 1 0 14168 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 14168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1688980957
transform 1 0 14168 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1688980957
transform 1 0 14168 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1688980957
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 13248 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 13800 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 13248 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 13800 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 12328 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 12880 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output147
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output148
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1688980957
transform 1 0 14168 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output150
timestamp 1688980957
transform 1 0 13432 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output151
timestamp 1688980957
transform 1 0 13432 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output152
timestamp 1688980957
transform 1 0 13248 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output153
timestamp 1688980957
transform 1 0 13800 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1688980957
transform 1 0 14168 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output155
timestamp 1688980957
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1688980957
transform 1 0 14168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output157
timestamp 1688980957
transform 1 0 13800 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output158
timestamp 1688980957
transform 1 0 13984 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1688980957
transform 1 0 14168 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output160
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output161
timestamp 1688980957
transform 1 0 13984 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output162
timestamp 1688980957
transform 1 0 12328 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output163
timestamp 1688980957
transform 1 0 12880 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output164
timestamp 1688980957
transform 1 0 13248 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output165
timestamp 1688980957
transform 1 0 13800 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output166
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output167
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output168
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output169
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output170
timestamp 1688980957
transform 1 0 13984 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output171
timestamp 1688980957
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1688980957
transform 1 0 14168 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output173
timestamp 1688980957
transform 1 0 13432 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output174
timestamp 1688980957
transform 1 0 13616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1688980957
transform 1 0 14168 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output176
timestamp 1688980957
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output177
timestamp 1688980957
transform 1 0 13248 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output178
timestamp 1688980957
transform 1 0 13800 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1688980957
transform 1 0 14168 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1688980957
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output181
timestamp 1688980957
transform 1 0 13248 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output182
timestamp 1688980957
transform 1 0 13800 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1688980957
transform 1 0 14168 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output184
timestamp 1688980957
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output185
timestamp 1688980957
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output186
timestamp 1688980957
transform 1 0 13248 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output187
timestamp 1688980957
transform 1 0 13800 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output188
timestamp 1688980957
transform 1 0 13064 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1688980957
transform 1 0 14168 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 13248 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 13800 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1688980957
transform 1 0 14168 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 9476 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output201
timestamp 1688980957
transform 1 0 12420 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 13156 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 13616 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 13432 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1688980957
transform 1 0 2116 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 2852 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1688980957
transform 1 0 4324 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 5060 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 6532 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1688980957
transform 1 0 7268 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1688980957
transform 1 0 8004 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output215
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14812 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14812 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14812 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14812 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14812 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 14812 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 14812 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 14812 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 14812 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 14812 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 14812 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 14812 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 14812 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 14812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 14812 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 14812 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 14812 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 14812 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 14812 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 14812 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 14812 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 14812 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 14812 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 14812 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 14812 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 14812 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 14812 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 14812 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 14812 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 14812 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 14812 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 14812 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 14812 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 14812 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 14812 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 14812 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 14812 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 14812 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 14812 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 14812 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 1564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 2116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 2852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 3220 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 4048 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 8464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 9936 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 10672 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 12144 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 12880 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 13984 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 2024 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 2852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 4784 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 5520 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 7912 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 8648 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 9292 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 10120 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 12236 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 12880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 14260 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 14260 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 11160 160 11280 0 FreeSans 480 0 0 0 A_I_top
port 0 nsew signal tristate
flabel metal3 s 0 9528 160 9648 0 FreeSans 480 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s 0 10344 160 10464 0 FreeSans 480 0 0 0 A_T_top
port 2 nsew signal tristate
flabel metal3 s 0 11976 160 12096 0 FreeSans 480 0 0 0 A_config_C_bit0
port 3 nsew signal tristate
flabel metal3 s 0 12792 160 12912 0 FreeSans 480 0 0 0 A_config_C_bit1
port 4 nsew signal tristate
flabel metal3 s 0 13608 160 13728 0 FreeSans 480 0 0 0 A_config_C_bit2
port 5 nsew signal tristate
flabel metal3 s 0 14424 160 14544 0 FreeSans 480 0 0 0 A_config_C_bit3
port 6 nsew signal tristate
flabel metal3 s 0 5448 160 5568 0 FreeSans 480 0 0 0 B_I_top
port 7 nsew signal tristate
flabel metal3 s 0 3816 160 3936 0 FreeSans 480 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s 0 4632 160 4752 0 FreeSans 480 0 0 0 B_T_top
port 9 nsew signal tristate
flabel metal3 s 0 6264 160 6384 0 FreeSans 480 0 0 0 B_config_C_bit0
port 10 nsew signal tristate
flabel metal3 s 0 7080 160 7200 0 FreeSans 480 0 0 0 B_config_C_bit1
port 11 nsew signal tristate
flabel metal3 s 0 7896 160 8016 0 FreeSans 480 0 0 0 B_config_C_bit2
port 12 nsew signal tristate
flabel metal3 s 0 8712 160 8832 0 FreeSans 480 0 0 0 B_config_C_bit3
port 13 nsew signal tristate
flabel metal3 s 15840 17960 16000 18080 0 FreeSans 480 0 0 0 E1BEG[0]
port 14 nsew signal tristate
flabel metal3 s 15840 18232 16000 18352 0 FreeSans 480 0 0 0 E1BEG[1]
port 15 nsew signal tristate
flabel metal3 s 15840 18504 16000 18624 0 FreeSans 480 0 0 0 E1BEG[2]
port 16 nsew signal tristate
flabel metal3 s 15840 18776 16000 18896 0 FreeSans 480 0 0 0 E1BEG[3]
port 17 nsew signal tristate
flabel metal3 s 15840 19048 16000 19168 0 FreeSans 480 0 0 0 E2BEG[0]
port 18 nsew signal tristate
flabel metal3 s 15840 19320 16000 19440 0 FreeSans 480 0 0 0 E2BEG[1]
port 19 nsew signal tristate
flabel metal3 s 15840 19592 16000 19712 0 FreeSans 480 0 0 0 E2BEG[2]
port 20 nsew signal tristate
flabel metal3 s 15840 19864 16000 19984 0 FreeSans 480 0 0 0 E2BEG[3]
port 21 nsew signal tristate
flabel metal3 s 15840 20136 16000 20256 0 FreeSans 480 0 0 0 E2BEG[4]
port 22 nsew signal tristate
flabel metal3 s 15840 20408 16000 20528 0 FreeSans 480 0 0 0 E2BEG[5]
port 23 nsew signal tristate
flabel metal3 s 15840 20680 16000 20800 0 FreeSans 480 0 0 0 E2BEG[6]
port 24 nsew signal tristate
flabel metal3 s 15840 20952 16000 21072 0 FreeSans 480 0 0 0 E2BEG[7]
port 25 nsew signal tristate
flabel metal3 s 15840 21224 16000 21344 0 FreeSans 480 0 0 0 E2BEGb[0]
port 26 nsew signal tristate
flabel metal3 s 15840 21496 16000 21616 0 FreeSans 480 0 0 0 E2BEGb[1]
port 27 nsew signal tristate
flabel metal3 s 15840 21768 16000 21888 0 FreeSans 480 0 0 0 E2BEGb[2]
port 28 nsew signal tristate
flabel metal3 s 15840 22040 16000 22160 0 FreeSans 480 0 0 0 E2BEGb[3]
port 29 nsew signal tristate
flabel metal3 s 15840 22312 16000 22432 0 FreeSans 480 0 0 0 E2BEGb[4]
port 30 nsew signal tristate
flabel metal3 s 15840 22584 16000 22704 0 FreeSans 480 0 0 0 E2BEGb[5]
port 31 nsew signal tristate
flabel metal3 s 15840 22856 16000 22976 0 FreeSans 480 0 0 0 E2BEGb[6]
port 32 nsew signal tristate
flabel metal3 s 15840 23128 16000 23248 0 FreeSans 480 0 0 0 E2BEGb[7]
port 33 nsew signal tristate
flabel metal3 s 15840 27752 16000 27872 0 FreeSans 480 0 0 0 E6BEG[0]
port 34 nsew signal tristate
flabel metal3 s 15840 30472 16000 30592 0 FreeSans 480 0 0 0 E6BEG[10]
port 35 nsew signal tristate
flabel metal3 s 15840 30744 16000 30864 0 FreeSans 480 0 0 0 E6BEG[11]
port 36 nsew signal tristate
flabel metal3 s 15840 28024 16000 28144 0 FreeSans 480 0 0 0 E6BEG[1]
port 37 nsew signal tristate
flabel metal3 s 15840 28296 16000 28416 0 FreeSans 480 0 0 0 E6BEG[2]
port 38 nsew signal tristate
flabel metal3 s 15840 28568 16000 28688 0 FreeSans 480 0 0 0 E6BEG[3]
port 39 nsew signal tristate
flabel metal3 s 15840 28840 16000 28960 0 FreeSans 480 0 0 0 E6BEG[4]
port 40 nsew signal tristate
flabel metal3 s 15840 29112 16000 29232 0 FreeSans 480 0 0 0 E6BEG[5]
port 41 nsew signal tristate
flabel metal3 s 15840 29384 16000 29504 0 FreeSans 480 0 0 0 E6BEG[6]
port 42 nsew signal tristate
flabel metal3 s 15840 29656 16000 29776 0 FreeSans 480 0 0 0 E6BEG[7]
port 43 nsew signal tristate
flabel metal3 s 15840 29928 16000 30048 0 FreeSans 480 0 0 0 E6BEG[8]
port 44 nsew signal tristate
flabel metal3 s 15840 30200 16000 30320 0 FreeSans 480 0 0 0 E6BEG[9]
port 45 nsew signal tristate
flabel metal3 s 15840 23400 16000 23520 0 FreeSans 480 0 0 0 EE4BEG[0]
port 46 nsew signal tristate
flabel metal3 s 15840 26120 16000 26240 0 FreeSans 480 0 0 0 EE4BEG[10]
port 47 nsew signal tristate
flabel metal3 s 15840 26392 16000 26512 0 FreeSans 480 0 0 0 EE4BEG[11]
port 48 nsew signal tristate
flabel metal3 s 15840 26664 16000 26784 0 FreeSans 480 0 0 0 EE4BEG[12]
port 49 nsew signal tristate
flabel metal3 s 15840 26936 16000 27056 0 FreeSans 480 0 0 0 EE4BEG[13]
port 50 nsew signal tristate
flabel metal3 s 15840 27208 16000 27328 0 FreeSans 480 0 0 0 EE4BEG[14]
port 51 nsew signal tristate
flabel metal3 s 15840 27480 16000 27600 0 FreeSans 480 0 0 0 EE4BEG[15]
port 52 nsew signal tristate
flabel metal3 s 15840 23672 16000 23792 0 FreeSans 480 0 0 0 EE4BEG[1]
port 53 nsew signal tristate
flabel metal3 s 15840 23944 16000 24064 0 FreeSans 480 0 0 0 EE4BEG[2]
port 54 nsew signal tristate
flabel metal3 s 15840 24216 16000 24336 0 FreeSans 480 0 0 0 EE4BEG[3]
port 55 nsew signal tristate
flabel metal3 s 15840 24488 16000 24608 0 FreeSans 480 0 0 0 EE4BEG[4]
port 56 nsew signal tristate
flabel metal3 s 15840 24760 16000 24880 0 FreeSans 480 0 0 0 EE4BEG[5]
port 57 nsew signal tristate
flabel metal3 s 15840 25032 16000 25152 0 FreeSans 480 0 0 0 EE4BEG[6]
port 58 nsew signal tristate
flabel metal3 s 15840 25304 16000 25424 0 FreeSans 480 0 0 0 EE4BEG[7]
port 59 nsew signal tristate
flabel metal3 s 15840 25576 16000 25696 0 FreeSans 480 0 0 0 EE4BEG[8]
port 60 nsew signal tristate
flabel metal3 s 15840 25848 16000 25968 0 FreeSans 480 0 0 0 EE4BEG[9]
port 61 nsew signal tristate
flabel metal3 s 0 15240 160 15360 0 FreeSans 480 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal3 s 0 23400 160 23520 0 FreeSans 480 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal3 s 0 24216 160 24336 0 FreeSans 480 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal3 s 0 25032 160 25152 0 FreeSans 480 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal3 s 0 25848 160 25968 0 FreeSans 480 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal3 s 0 26664 160 26784 0 FreeSans 480 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal3 s 0 27480 160 27600 0 FreeSans 480 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal3 s 0 28296 160 28416 0 FreeSans 480 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal3 s 0 29112 160 29232 0 FreeSans 480 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal3 s 0 29928 160 30048 0 FreeSans 480 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal3 s 0 30744 160 30864 0 FreeSans 480 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal3 s 0 16056 160 16176 0 FreeSans 480 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal3 s 0 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal3 s 0 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal3 s 0 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal3 s 0 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal3 s 0 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal3 s 0 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal3 s 0 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal3 s 0 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal3 s 0 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal3 s 0 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal3 s 0 16872 160 16992 0 FreeSans 480 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal3 s 0 39720 160 39840 0 FreeSans 480 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal3 s 0 40536 160 40656 0 FreeSans 480 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal3 s 0 17688 160 17808 0 FreeSans 480 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal3 s 0 18504 160 18624 0 FreeSans 480 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal3 s 0 19320 160 19440 0 FreeSans 480 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal3 s 0 20136 160 20256 0 FreeSans 480 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal3 s 0 20952 160 21072 0 FreeSans 480 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal3 s 0 21768 160 21888 0 FreeSans 480 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal3 s 0 22584 160 22704 0 FreeSans 480 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal3 s 15840 31016 16000 31136 0 FreeSans 480 0 0 0 FrameData_O[0]
port 94 nsew signal tristate
flabel metal3 s 15840 33736 16000 33856 0 FreeSans 480 0 0 0 FrameData_O[10]
port 95 nsew signal tristate
flabel metal3 s 15840 34008 16000 34128 0 FreeSans 480 0 0 0 FrameData_O[11]
port 96 nsew signal tristate
flabel metal3 s 15840 34280 16000 34400 0 FreeSans 480 0 0 0 FrameData_O[12]
port 97 nsew signal tristate
flabel metal3 s 15840 34552 16000 34672 0 FreeSans 480 0 0 0 FrameData_O[13]
port 98 nsew signal tristate
flabel metal3 s 15840 34824 16000 34944 0 FreeSans 480 0 0 0 FrameData_O[14]
port 99 nsew signal tristate
flabel metal3 s 15840 35096 16000 35216 0 FreeSans 480 0 0 0 FrameData_O[15]
port 100 nsew signal tristate
flabel metal3 s 15840 35368 16000 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 101 nsew signal tristate
flabel metal3 s 15840 35640 16000 35760 0 FreeSans 480 0 0 0 FrameData_O[17]
port 102 nsew signal tristate
flabel metal3 s 15840 35912 16000 36032 0 FreeSans 480 0 0 0 FrameData_O[18]
port 103 nsew signal tristate
flabel metal3 s 15840 36184 16000 36304 0 FreeSans 480 0 0 0 FrameData_O[19]
port 104 nsew signal tristate
flabel metal3 s 15840 31288 16000 31408 0 FreeSans 480 0 0 0 FrameData_O[1]
port 105 nsew signal tristate
flabel metal3 s 15840 36456 16000 36576 0 FreeSans 480 0 0 0 FrameData_O[20]
port 106 nsew signal tristate
flabel metal3 s 15840 36728 16000 36848 0 FreeSans 480 0 0 0 FrameData_O[21]
port 107 nsew signal tristate
flabel metal3 s 15840 37000 16000 37120 0 FreeSans 480 0 0 0 FrameData_O[22]
port 108 nsew signal tristate
flabel metal3 s 15840 37272 16000 37392 0 FreeSans 480 0 0 0 FrameData_O[23]
port 109 nsew signal tristate
flabel metal3 s 15840 37544 16000 37664 0 FreeSans 480 0 0 0 FrameData_O[24]
port 110 nsew signal tristate
flabel metal3 s 15840 37816 16000 37936 0 FreeSans 480 0 0 0 FrameData_O[25]
port 111 nsew signal tristate
flabel metal3 s 15840 38088 16000 38208 0 FreeSans 480 0 0 0 FrameData_O[26]
port 112 nsew signal tristate
flabel metal3 s 15840 38360 16000 38480 0 FreeSans 480 0 0 0 FrameData_O[27]
port 113 nsew signal tristate
flabel metal3 s 15840 38632 16000 38752 0 FreeSans 480 0 0 0 FrameData_O[28]
port 114 nsew signal tristate
flabel metal3 s 15840 38904 16000 39024 0 FreeSans 480 0 0 0 FrameData_O[29]
port 115 nsew signal tristate
flabel metal3 s 15840 31560 16000 31680 0 FreeSans 480 0 0 0 FrameData_O[2]
port 116 nsew signal tristate
flabel metal3 s 15840 39176 16000 39296 0 FreeSans 480 0 0 0 FrameData_O[30]
port 117 nsew signal tristate
flabel metal3 s 15840 39448 16000 39568 0 FreeSans 480 0 0 0 FrameData_O[31]
port 118 nsew signal tristate
flabel metal3 s 15840 31832 16000 31952 0 FreeSans 480 0 0 0 FrameData_O[3]
port 119 nsew signal tristate
flabel metal3 s 15840 32104 16000 32224 0 FreeSans 480 0 0 0 FrameData_O[4]
port 120 nsew signal tristate
flabel metal3 s 15840 32376 16000 32496 0 FreeSans 480 0 0 0 FrameData_O[5]
port 121 nsew signal tristate
flabel metal3 s 15840 32648 16000 32768 0 FreeSans 480 0 0 0 FrameData_O[6]
port 122 nsew signal tristate
flabel metal3 s 15840 32920 16000 33040 0 FreeSans 480 0 0 0 FrameData_O[7]
port 123 nsew signal tristate
flabel metal3 s 15840 33192 16000 33312 0 FreeSans 480 0 0 0 FrameData_O[8]
port 124 nsew signal tristate
flabel metal3 s 15840 33464 16000 33584 0 FreeSans 480 0 0 0 FrameData_O[9]
port 125 nsew signal tristate
flabel metal2 s 1306 0 1362 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal2 s 8666 0 8722 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal2 s 9402 0 9458 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal2 s 10138 0 10194 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal2 s 10874 0 10930 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal2 s 11610 0 11666 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal2 s 12346 0 12402 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal2 s 13082 0 13138 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal2 s 13818 0 13874 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal2 s 14554 0 14610 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal2 s 15290 0 15346 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal2 s 2042 0 2098 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal2 s 2778 0 2834 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal2 s 3514 0 3570 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal2 s 4250 0 4306 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal2 s 4986 0 5042 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal2 s 5722 0 5778 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal2 s 6458 0 6514 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal2 s 7194 0 7250 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal2 s 7930 0 7986 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal2 s 1306 44463 1362 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 146 nsew signal tristate
flabel metal2 s 8666 44463 8722 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 147 nsew signal tristate
flabel metal2 s 9402 44463 9458 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 148 nsew signal tristate
flabel metal2 s 10138 44463 10194 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 149 nsew signal tristate
flabel metal2 s 10874 44463 10930 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 150 nsew signal tristate
flabel metal2 s 11610 44463 11666 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 151 nsew signal tristate
flabel metal2 s 12346 44463 12402 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 152 nsew signal tristate
flabel metal2 s 13082 44463 13138 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 153 nsew signal tristate
flabel metal2 s 13818 44463 13874 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 154 nsew signal tristate
flabel metal2 s 14554 44463 14610 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 155 nsew signal tristate
flabel metal2 s 15290 44463 15346 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 156 nsew signal tristate
flabel metal2 s 2042 44463 2098 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 157 nsew signal tristate
flabel metal2 s 2778 44463 2834 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 158 nsew signal tristate
flabel metal2 s 3514 44463 3570 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 159 nsew signal tristate
flabel metal2 s 4250 44463 4306 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 160 nsew signal tristate
flabel metal2 s 4986 44463 5042 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 161 nsew signal tristate
flabel metal2 s 5722 44463 5778 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 162 nsew signal tristate
flabel metal2 s 6458 44463 6514 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 163 nsew signal tristate
flabel metal2 s 7194 44463 7250 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 164 nsew signal tristate
flabel metal2 s 7930 44463 7986 44623 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 165 nsew signal tristate
flabel metal2 s 570 0 626 160 0 FreeSans 224 90 0 0 UserCLK
port 166 nsew signal input
flabel metal2 s 570 44463 626 44623 0 FreeSans 224 90 0 0 UserCLKo
port 167 nsew signal tristate
flabel metal4 s 4370 1040 4690 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 7797 1040 8117 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 11224 1040 11544 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 14651 1040 14971 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 2657 1040 2977 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 6084 1040 6404 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 9511 1040 9831 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 12938 1040 13258 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal3 s 15840 4904 16000 5024 0 FreeSans 480 0 0 0 W1END[0]
port 170 nsew signal input
flabel metal3 s 15840 5176 16000 5296 0 FreeSans 480 0 0 0 W1END[1]
port 171 nsew signal input
flabel metal3 s 15840 5448 16000 5568 0 FreeSans 480 0 0 0 W1END[2]
port 172 nsew signal input
flabel metal3 s 15840 5720 16000 5840 0 FreeSans 480 0 0 0 W1END[3]
port 173 nsew signal input
flabel metal3 s 15840 8168 16000 8288 0 FreeSans 480 0 0 0 W2END[0]
port 174 nsew signal input
flabel metal3 s 15840 8440 16000 8560 0 FreeSans 480 0 0 0 W2END[1]
port 175 nsew signal input
flabel metal3 s 15840 8712 16000 8832 0 FreeSans 480 0 0 0 W2END[2]
port 176 nsew signal input
flabel metal3 s 15840 8984 16000 9104 0 FreeSans 480 0 0 0 W2END[3]
port 177 nsew signal input
flabel metal3 s 15840 9256 16000 9376 0 FreeSans 480 0 0 0 W2END[4]
port 178 nsew signal input
flabel metal3 s 15840 9528 16000 9648 0 FreeSans 480 0 0 0 W2END[5]
port 179 nsew signal input
flabel metal3 s 15840 9800 16000 9920 0 FreeSans 480 0 0 0 W2END[6]
port 180 nsew signal input
flabel metal3 s 15840 10072 16000 10192 0 FreeSans 480 0 0 0 W2END[7]
port 181 nsew signal input
flabel metal3 s 15840 5992 16000 6112 0 FreeSans 480 0 0 0 W2MID[0]
port 182 nsew signal input
flabel metal3 s 15840 6264 16000 6384 0 FreeSans 480 0 0 0 W2MID[1]
port 183 nsew signal input
flabel metal3 s 15840 6536 16000 6656 0 FreeSans 480 0 0 0 W2MID[2]
port 184 nsew signal input
flabel metal3 s 15840 6808 16000 6928 0 FreeSans 480 0 0 0 W2MID[3]
port 185 nsew signal input
flabel metal3 s 15840 7080 16000 7200 0 FreeSans 480 0 0 0 W2MID[4]
port 186 nsew signal input
flabel metal3 s 15840 7352 16000 7472 0 FreeSans 480 0 0 0 W2MID[5]
port 187 nsew signal input
flabel metal3 s 15840 7624 16000 7744 0 FreeSans 480 0 0 0 W2MID[6]
port 188 nsew signal input
flabel metal3 s 15840 7896 16000 8016 0 FreeSans 480 0 0 0 W2MID[7]
port 189 nsew signal input
flabel metal3 s 15840 14696 16000 14816 0 FreeSans 480 0 0 0 W6END[0]
port 190 nsew signal input
flabel metal3 s 15840 17416 16000 17536 0 FreeSans 480 0 0 0 W6END[10]
port 191 nsew signal input
flabel metal3 s 15840 17688 16000 17808 0 FreeSans 480 0 0 0 W6END[11]
port 192 nsew signal input
flabel metal3 s 15840 14968 16000 15088 0 FreeSans 480 0 0 0 W6END[1]
port 193 nsew signal input
flabel metal3 s 15840 15240 16000 15360 0 FreeSans 480 0 0 0 W6END[2]
port 194 nsew signal input
flabel metal3 s 15840 15512 16000 15632 0 FreeSans 480 0 0 0 W6END[3]
port 195 nsew signal input
flabel metal3 s 15840 15784 16000 15904 0 FreeSans 480 0 0 0 W6END[4]
port 196 nsew signal input
flabel metal3 s 15840 16056 16000 16176 0 FreeSans 480 0 0 0 W6END[5]
port 197 nsew signal input
flabel metal3 s 15840 16328 16000 16448 0 FreeSans 480 0 0 0 W6END[6]
port 198 nsew signal input
flabel metal3 s 15840 16600 16000 16720 0 FreeSans 480 0 0 0 W6END[7]
port 199 nsew signal input
flabel metal3 s 15840 16872 16000 16992 0 FreeSans 480 0 0 0 W6END[8]
port 200 nsew signal input
flabel metal3 s 15840 17144 16000 17264 0 FreeSans 480 0 0 0 W6END[9]
port 201 nsew signal input
flabel metal3 s 15840 10344 16000 10464 0 FreeSans 480 0 0 0 WW4END[0]
port 202 nsew signal input
flabel metal3 s 15840 13064 16000 13184 0 FreeSans 480 0 0 0 WW4END[10]
port 203 nsew signal input
flabel metal3 s 15840 13336 16000 13456 0 FreeSans 480 0 0 0 WW4END[11]
port 204 nsew signal input
flabel metal3 s 15840 13608 16000 13728 0 FreeSans 480 0 0 0 WW4END[12]
port 205 nsew signal input
flabel metal3 s 15840 13880 16000 14000 0 FreeSans 480 0 0 0 WW4END[13]
port 206 nsew signal input
flabel metal3 s 15840 14152 16000 14272 0 FreeSans 480 0 0 0 WW4END[14]
port 207 nsew signal input
flabel metal3 s 15840 14424 16000 14544 0 FreeSans 480 0 0 0 WW4END[15]
port 208 nsew signal input
flabel metal3 s 15840 10616 16000 10736 0 FreeSans 480 0 0 0 WW4END[1]
port 209 nsew signal input
flabel metal3 s 15840 10888 16000 11008 0 FreeSans 480 0 0 0 WW4END[2]
port 210 nsew signal input
flabel metal3 s 15840 11160 16000 11280 0 FreeSans 480 0 0 0 WW4END[3]
port 211 nsew signal input
flabel metal3 s 15840 11432 16000 11552 0 FreeSans 480 0 0 0 WW4END[4]
port 212 nsew signal input
flabel metal3 s 15840 11704 16000 11824 0 FreeSans 480 0 0 0 WW4END[5]
port 213 nsew signal input
flabel metal3 s 15840 11976 16000 12096 0 FreeSans 480 0 0 0 WW4END[6]
port 214 nsew signal input
flabel metal3 s 15840 12248 16000 12368 0 FreeSans 480 0 0 0 WW4END[7]
port 215 nsew signal input
flabel metal3 s 15840 12520 16000 12640 0 FreeSans 480 0 0 0 WW4END[8]
port 216 nsew signal input
flabel metal3 s 15840 12792 16000 12912 0 FreeSans 480 0 0 0 WW4END[9]
port 217 nsew signal input
rlabel via1 8037 43520 8037 43520 0 VGND
rlabel metal1 7958 42976 7958 42976 0 VPWR
rlabel metal3 498 11220 498 11220 0 A_I_top
rlabel metal3 544 9588 544 9588 0 A_O_top
rlabel metal3 498 10404 498 10404 0 A_T_top
rlabel metal3 498 12036 498 12036 0 A_config_C_bit0
rlabel metal3 567 12852 567 12852 0 A_config_C_bit1
rlabel metal3 1326 13668 1326 13668 0 A_config_C_bit2
rlabel metal3 498 14484 498 14484 0 A_config_C_bit3
rlabel metal3 498 5508 498 5508 0 B_I_top
rlabel metal3 452 3876 452 3876 0 B_O_top
rlabel metal3 544 4692 544 4692 0 B_T_top
rlabel metal3 498 6324 498 6324 0 B_config_C_bit0
rlabel metal3 498 7140 498 7140 0 B_config_C_bit1
rlabel metal3 567 7956 567 7956 0 B_config_C_bit2
rlabel metal3 475 8772 475 8772 0 B_config_C_bit3
rlabel metal1 13340 17850 13340 17850 0 E1BEG[0]
rlabel metal1 14720 17306 14720 17306 0 E1BEG[1]
rlabel metal1 14766 17850 14766 17850 0 E1BEG[2]
rlabel metal3 15188 18836 15188 18836 0 E1BEG[3]
rlabel metal1 14030 18394 14030 18394 0 E2BEG[0]
rlabel metal1 12236 18938 12236 18938 0 E2BEG[1]
rlabel metal3 15533 19652 15533 19652 0 E2BEG[2]
rlabel metal1 14720 17782 14720 17782 0 E2BEG[3]
rlabel metal2 14398 19839 14398 19839 0 E2BEG[4]
rlabel metal1 14076 19482 14076 19482 0 E2BEG[5]
rlabel metal1 14490 18292 14490 18292 0 E2BEG[6]
rlabel metal3 14866 21012 14866 21012 0 E2BEG[7]
rlabel metal1 14076 20026 14076 20026 0 E2BEGb[0]
rlabel metal3 15096 21556 15096 21556 0 E2BEGb[1]
rlabel metal1 14766 21114 14766 21114 0 E2BEGb[2]
rlabel metal1 14444 21658 14444 21658 0 E2BEGb[3]
rlabel metal3 15418 22372 15418 22372 0 E2BEGb[4]
rlabel metal1 14444 22202 14444 22202 0 E2BEGb[5]
rlabel metal3 15510 22916 15510 22916 0 E2BEGb[6]
rlabel metal3 15142 23188 15142 23188 0 E2BEGb[7]
rlabel metal3 15142 27812 15142 27812 0 E6BEG[0]
rlabel metal3 15510 30532 15510 30532 0 E6BEG[10]
rlabel metal1 13892 31654 13892 31654 0 E6BEG[11]
rlabel metal3 14866 28084 14866 28084 0 E6BEG[1]
rlabel metal3 15510 28356 15510 28356 0 E6BEG[2]
rlabel metal3 15050 28628 15050 28628 0 E6BEG[3]
rlabel metal3 15234 28900 15234 28900 0 E6BEG[4]
rlabel metal3 15096 29172 15096 29172 0 E6BEG[5]
rlabel metal3 15510 29444 15510 29444 0 E6BEG[6]
rlabel metal3 15602 29716 15602 29716 0 E6BEG[7]
rlabel metal3 15073 29988 15073 29988 0 E6BEG[8]
rlabel metal3 14636 30260 14636 30260 0 E6BEG[9]
rlabel metal3 15142 23460 15142 23460 0 EE4BEG[0]
rlabel metal3 15510 26180 15510 26180 0 EE4BEG[10]
rlabel metal3 15418 26452 15418 26452 0 EE4BEG[11]
rlabel metal3 14866 26724 14866 26724 0 EE4BEG[12]
rlabel metal3 14912 26996 14912 26996 0 EE4BEG[13]
rlabel metal3 15510 27268 15510 27268 0 EE4BEG[14]
rlabel metal3 15050 27540 15050 27540 0 EE4BEG[15]
rlabel metal3 15142 23732 15142 23732 0 EE4BEG[1]
rlabel metal3 15510 24004 15510 24004 0 EE4BEG[2]
rlabel metal3 15142 24276 15142 24276 0 EE4BEG[3]
rlabel metal3 15050 24548 15050 24548 0 EE4BEG[4]
rlabel metal3 15510 24820 15510 24820 0 EE4BEG[5]
rlabel metal3 15533 25092 15533 25092 0 EE4BEG[6]
rlabel metal3 14866 25364 14866 25364 0 EE4BEG[7]
rlabel metal3 15602 25636 15602 25636 0 EE4BEG[8]
rlabel metal2 12374 26333 12374 26333 0 EE4BEG[9]
rlabel metal3 498 15300 498 15300 0 FrameData[0]
rlabel metal3 452 23460 452 23460 0 FrameData[10]
rlabel metal3 452 24276 452 24276 0 FrameData[11]
rlabel metal3 452 25092 452 25092 0 FrameData[12]
rlabel metal3 475 25908 475 25908 0 FrameData[13]
rlabel metal3 452 26724 452 26724 0 FrameData[14]
rlabel metal3 820 27540 820 27540 0 FrameData[15]
rlabel metal3 452 28356 452 28356 0 FrameData[16]
rlabel metal3 452 29172 452 29172 0 FrameData[17]
rlabel metal3 452 29988 452 29988 0 FrameData[18]
rlabel metal3 452 30804 452 30804 0 FrameData[19]
rlabel metal3 452 16116 452 16116 0 FrameData[1]
rlabel metal3 774 31620 774 31620 0 FrameData[20]
rlabel metal3 452 32436 452 32436 0 FrameData[21]
rlabel metal3 452 33252 452 33252 0 FrameData[22]
rlabel metal3 475 34068 475 34068 0 FrameData[23]
rlabel metal3 452 34884 452 34884 0 FrameData[24]
rlabel metal3 475 35700 475 35700 0 FrameData[25]
rlabel metal3 452 36516 452 36516 0 FrameData[26]
rlabel metal3 452 37332 452 37332 0 FrameData[27]
rlabel metal3 452 38148 452 38148 0 FrameData[28]
rlabel metal3 452 38964 452 38964 0 FrameData[29]
rlabel metal3 452 16932 452 16932 0 FrameData[2]
rlabel metal3 774 39780 774 39780 0 FrameData[30]
rlabel metal3 452 40596 452 40596 0 FrameData[31]
rlabel metal3 475 17748 475 17748 0 FrameData[3]
rlabel metal3 452 18564 452 18564 0 FrameData[4]
rlabel metal3 452 19380 452 19380 0 FrameData[5]
rlabel metal3 452 20196 452 20196 0 FrameData[6]
rlabel metal3 452 21012 452 21012 0 FrameData[7]
rlabel metal3 452 21828 452 21828 0 FrameData[8]
rlabel metal3 452 22644 452 22644 0 FrameData[9]
rlabel metal1 13340 31654 13340 31654 0 FrameData_O[0]
rlabel metal3 15510 33796 15510 33796 0 FrameData_O[10]
rlabel metal3 15050 34068 15050 34068 0 FrameData_O[11]
rlabel metal3 15142 34340 15142 34340 0 FrameData_O[12]
rlabel metal3 14912 34612 14912 34612 0 FrameData_O[13]
rlabel metal3 15510 34884 15510 34884 0 FrameData_O[14]
rlabel metal3 14866 35156 14866 35156 0 FrameData_O[15]
rlabel metal3 15625 35428 15625 35428 0 FrameData_O[16]
rlabel metal3 14820 35700 14820 35700 0 FrameData_O[17]
rlabel metal3 15510 35972 15510 35972 0 FrameData_O[18]
rlabel metal3 14866 36244 14866 36244 0 FrameData_O[19]
rlabel metal3 14958 31348 14958 31348 0 FrameData_O[1]
rlabel metal3 15142 36516 15142 36516 0 FrameData_O[20]
rlabel metal3 14774 36788 14774 36788 0 FrameData_O[21]
rlabel metal3 15510 37060 15510 37060 0 FrameData_O[22]
rlabel metal3 15050 37332 15050 37332 0 FrameData_O[23]
rlabel metal3 15142 37604 15142 37604 0 FrameData_O[24]
rlabel metal3 14866 37876 14866 37876 0 FrameData_O[25]
rlabel metal3 15510 38148 15510 38148 0 FrameData_O[26]
rlabel metal3 15050 38420 15050 38420 0 FrameData_O[27]
rlabel metal3 15142 38692 15142 38692 0 FrameData_O[28]
rlabel metal3 14912 38964 14912 38964 0 FrameData_O[29]
rlabel metal1 14536 32810 14536 32810 0 FrameData_O[2]
rlabel metal3 15510 39236 15510 39236 0 FrameData_O[30]
rlabel metal3 15050 39508 15050 39508 0 FrameData_O[31]
rlabel metal3 14912 31892 14912 31892 0 FrameData_O[3]
rlabel metal3 15142 32164 15142 32164 0 FrameData_O[4]
rlabel metal3 15096 32436 15096 32436 0 FrameData_O[5]
rlabel metal3 15510 32708 15510 32708 0 FrameData_O[6]
rlabel metal3 15050 32980 15050 32980 0 FrameData_O[7]
rlabel metal3 15142 33252 15142 33252 0 FrameData_O[8]
rlabel metal3 14912 33524 14912 33524 0 FrameData_O[9]
rlabel metal2 1334 704 1334 704 0 FrameStrobe[0]
rlabel metal2 8694 704 8694 704 0 FrameStrobe[10]
rlabel metal2 9430 143 9430 143 0 FrameStrobe[11]
rlabel metal2 10311 68 10311 68 0 FrameStrobe[12]
rlabel metal2 10902 704 10902 704 0 FrameStrobe[13]
rlabel metal2 11638 704 11638 704 0 FrameStrobe[14]
rlabel metal2 12374 704 12374 704 0 FrameStrobe[15]
rlabel metal2 13110 143 13110 143 0 FrameStrobe[16]
rlabel metal2 13899 68 13899 68 0 FrameStrobe[17]
rlabel metal2 14582 704 14582 704 0 FrameStrobe[18]
rlabel metal2 15318 534 15318 534 0 FrameStrobe[19]
rlabel metal2 2123 68 2123 68 0 FrameStrobe[1]
rlabel metal1 2760 1326 2760 1326 0 FrameStrobe[2]
rlabel metal2 3687 68 3687 68 0 FrameStrobe[3]
rlabel metal2 4278 704 4278 704 0 FrameStrobe[4]
rlabel metal2 5014 704 5014 704 0 FrameStrobe[5]
rlabel metal2 5750 704 5750 704 0 FrameStrobe[6]
rlabel metal2 6486 704 6486 704 0 FrameStrobe[7]
rlabel metal2 7367 68 7367 68 0 FrameStrobe[8]
rlabel metal2 8103 68 8103 68 0 FrameStrobe[9]
rlabel metal2 1334 43785 1334 43785 0 FrameStrobe_O[0]
rlabel metal1 8924 43418 8924 43418 0 FrameStrobe_O[10]
rlabel metal2 9430 43972 9430 43972 0 FrameStrobe_O[11]
rlabel metal1 10304 43418 10304 43418 0 FrameStrobe_O[12]
rlabel metal2 10902 43972 10902 43972 0 FrameStrobe_O[13]
rlabel metal1 12006 43078 12006 43078 0 FrameStrobe_O[14]
rlabel metal2 12374 43972 12374 43972 0 FrameStrobe_O[15]
rlabel metal1 13248 43418 13248 43418 0 FrameStrobe_O[16]
rlabel metal1 14076 43418 14076 43418 0 FrameStrobe_O[17]
rlabel metal1 14214 43146 14214 43146 0 FrameStrobe_O[18]
rlabel metal1 14582 42738 14582 42738 0 FrameStrobe_O[19]
rlabel metal1 2208 43146 2208 43146 0 FrameStrobe_O[1]
rlabel metal2 2806 43972 2806 43972 0 FrameStrobe_O[2]
rlabel metal1 3772 43418 3772 43418 0 FrameStrobe_O[3]
rlabel metal1 4416 43418 4416 43418 0 FrameStrobe_O[4]
rlabel metal1 5152 43418 5152 43418 0 FrameStrobe_O[5]
rlabel metal1 5888 43418 5888 43418 0 FrameStrobe_O[6]
rlabel metal1 6624 43418 6624 43418 0 FrameStrobe_O[7]
rlabel metal1 7360 43418 7360 43418 0 FrameStrobe_O[8]
rlabel metal2 8234 43979 8234 43979 0 FrameStrobe_O[9]
rlabel metal1 2162 10710 2162 10710 0 Inst_A_IO_1_bidirectional_frame_config_pass.I
rlabel metal1 6210 17544 6210 17544 0 Inst_A_IO_1_bidirectional_frame_config_pass.O
rlabel metal2 5566 18836 5566 18836 0 Inst_A_IO_1_bidirectional_frame_config_pass.Q
rlabel metal1 1610 9486 1610 9486 0 Inst_A_IO_1_bidirectional_frame_config_pass.T
rlabel metal1 2346 12206 2346 12206 0 Inst_A_config_Config_access.ConfigBits\[0\]
rlabel metal2 2530 12682 2530 12682 0 Inst_A_config_Config_access.ConfigBits\[1\]
rlabel metal1 2346 14382 2346 14382 0 Inst_A_config_Config_access.ConfigBits\[2\]
rlabel metal2 2530 14858 2530 14858 0 Inst_A_config_Config_access.ConfigBits\[3\]
rlabel metal1 2254 6324 2254 6324 0 Inst_B_IO_1_bidirectional_frame_config_pass.I
rlabel via1 6574 19822 6574 19822 0 Inst_B_IO_1_bidirectional_frame_config_pass.O
rlabel metal2 12650 28628 12650 28628 0 Inst_B_IO_1_bidirectional_frame_config_pass.Q
rlabel metal2 4002 7276 4002 7276 0 Inst_B_IO_1_bidirectional_frame_config_pass.T
rlabel metal1 2484 5882 2484 5882 0 Inst_B_config_Config_access.ConfigBits\[0\]
rlabel metal1 2300 6970 2300 6970 0 Inst_B_config_Config_access.ConfigBits\[1\]
rlabel metal1 2392 9554 2392 9554 0 Inst_B_config_Config_access.ConfigBits\[2\]
rlabel metal1 2392 8466 2392 8466 0 Inst_B_config_Config_access.ConfigBits\[3\]
rlabel metal1 10304 5746 10304 5746 0 Inst_W_IO_ConfigMem.ConfigBits\[100\]
rlabel metal2 10994 5950 10994 5950 0 Inst_W_IO_ConfigMem.ConfigBits\[101\]
rlabel metal1 12190 8364 12190 8364 0 Inst_W_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 12558 8058 12558 8058 0 Inst_W_IO_ConfigMem.ConfigBits\[103\]
rlabel metal2 7590 7718 7590 7718 0 Inst_W_IO_ConfigMem.ConfigBits\[104\]
rlabel metal2 9154 6596 9154 6596 0 Inst_W_IO_ConfigMem.ConfigBits\[105\]
rlabel metal1 6164 8466 6164 8466 0 Inst_W_IO_ConfigMem.ConfigBits\[106\]
rlabel metal2 9430 5066 9430 5066 0 Inst_W_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 10488 6222 10488 6222 0 Inst_W_IO_ConfigMem.ConfigBits\[108\]
rlabel metal1 11454 4794 11454 4794 0 Inst_W_IO_ConfigMem.ConfigBits\[109\]
rlabel metal1 6578 20468 6578 20468 0 Inst_W_IO_ConfigMem.ConfigBits\[10\]
rlabel metal2 12788 4794 12788 4794 0 Inst_W_IO_ConfigMem.ConfigBits\[110\]
rlabel metal1 7084 10166 7084 10166 0 Inst_W_IO_ConfigMem.ConfigBits\[111\]
rlabel metal2 8142 10234 8142 10234 0 Inst_W_IO_ConfigMem.ConfigBits\[112\]
rlabel metal1 5014 10064 5014 10064 0 Inst_W_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 9108 20910 9108 20910 0 Inst_W_IO_ConfigMem.ConfigBits\[11\]
rlabel metal1 7406 14926 7406 14926 0 Inst_W_IO_ConfigMem.ConfigBits\[12\]
rlabel metal1 7820 14586 7820 14586 0 Inst_W_IO_ConfigMem.ConfigBits\[13\]
rlabel metal1 7866 15946 7866 15946 0 Inst_W_IO_ConfigMem.ConfigBits\[14\]
rlabel metal2 8694 16388 8694 16388 0 Inst_W_IO_ConfigMem.ConfigBits\[15\]
rlabel metal1 7406 13974 7406 13974 0 Inst_W_IO_ConfigMem.ConfigBits\[16\]
rlabel metal1 6624 13498 6624 13498 0 Inst_W_IO_ConfigMem.ConfigBits\[17\]
rlabel metal1 10258 16218 10258 16218 0 Inst_W_IO_ConfigMem.ConfigBits\[18\]
rlabel metal1 10534 16762 10534 16762 0 Inst_W_IO_ConfigMem.ConfigBits\[19\]
rlabel metal1 13064 12954 13064 12954 0 Inst_W_IO_ConfigMem.ConfigBits\[20\]
rlabel metal2 13294 13209 13294 13209 0 Inst_W_IO_ConfigMem.ConfigBits\[21\]
rlabel metal2 13294 15844 13294 15844 0 Inst_W_IO_ConfigMem.ConfigBits\[22\]
rlabel metal2 13846 15606 13846 15606 0 Inst_W_IO_ConfigMem.ConfigBits\[23\]
rlabel metal1 10120 19278 10120 19278 0 Inst_W_IO_ConfigMem.ConfigBits\[24\]
rlabel metal1 10856 18938 10856 18938 0 Inst_W_IO_ConfigMem.ConfigBits\[25\]
rlabel metal2 12190 17306 12190 17306 0 Inst_W_IO_ConfigMem.ConfigBits\[26\]
rlabel metal2 12742 17612 12742 17612 0 Inst_W_IO_ConfigMem.ConfigBits\[27\]
rlabel metal1 10856 21046 10856 21046 0 Inst_W_IO_ConfigMem.ConfigBits\[28\]
rlabel metal1 11638 20978 11638 20978 0 Inst_W_IO_ConfigMem.ConfigBits\[29\]
rlabel metal1 8280 22542 8280 22542 0 Inst_W_IO_ConfigMem.ConfigBits\[30\]
rlabel metal2 8878 23324 8878 23324 0 Inst_W_IO_ConfigMem.ConfigBits\[31\]
rlabel metal1 8050 12750 8050 12750 0 Inst_W_IO_ConfigMem.ConfigBits\[32\]
rlabel metal2 8786 12988 8786 12988 0 Inst_W_IO_ConfigMem.ConfigBits\[33\]
rlabel metal1 10074 14586 10074 14586 0 Inst_W_IO_ConfigMem.ConfigBits\[34\]
rlabel metal2 10718 15164 10718 15164 0 Inst_W_IO_ConfigMem.ConfigBits\[35\]
rlabel metal1 7130 11322 7130 11322 0 Inst_W_IO_ConfigMem.ConfigBits\[36\]
rlabel metal1 8004 11866 8004 11866 0 Inst_W_IO_ConfigMem.ConfigBits\[37\]
rlabel metal1 13202 10234 13202 10234 0 Inst_W_IO_ConfigMem.ConfigBits\[38\]
rlabel metal1 13800 10778 13800 10778 0 Inst_W_IO_ConfigMem.ConfigBits\[39\]
rlabel metal1 12190 7242 12190 7242 0 Inst_W_IO_ConfigMem.ConfigBits\[40\]
rlabel metal1 13938 3910 13938 3910 0 Inst_W_IO_ConfigMem.ConfigBits\[41\]
rlabel metal1 12144 11322 12144 11322 0 Inst_W_IO_ConfigMem.ConfigBits\[42\]
rlabel metal1 13110 11322 13110 11322 0 Inst_W_IO_ConfigMem.ConfigBits\[43\]
rlabel metal1 5796 23222 5796 23222 0 Inst_W_IO_ConfigMem.ConfigBits\[44\]
rlabel metal1 6670 22202 6670 22202 0 Inst_W_IO_ConfigMem.ConfigBits\[45\]
rlabel metal2 12650 23834 12650 23834 0 Inst_W_IO_ConfigMem.ConfigBits\[46\]
rlabel via1 13202 23715 13202 23715 0 Inst_W_IO_ConfigMem.ConfigBits\[47\]
rlabel metal1 7590 29784 7590 29784 0 Inst_W_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 8096 31926 8096 31926 0 Inst_W_IO_ConfigMem.ConfigBits\[49\]
rlabel metal1 10304 28662 10304 28662 0 Inst_W_IO_ConfigMem.ConfigBits\[50\]
rlabel metal1 10856 28186 10856 28186 0 Inst_W_IO_ConfigMem.ConfigBits\[51\]
rlabel metal2 10534 12517 10534 12517 0 Inst_W_IO_ConfigMem.ConfigBits\[52\]
rlabel metal2 10580 12172 10580 12172 0 Inst_W_IO_ConfigMem.ConfigBits\[53\]
rlabel metal1 12512 9894 12512 9894 0 Inst_W_IO_ConfigMem.ConfigBits\[54\]
rlabel metal1 12742 10064 12742 10064 0 Inst_W_IO_ConfigMem.ConfigBits\[55\]
rlabel metal1 12696 16626 12696 16626 0 Inst_W_IO_ConfigMem.ConfigBits\[56\]
rlabel metal2 13294 17612 13294 17612 0 Inst_W_IO_ConfigMem.ConfigBits\[57\]
rlabel metal1 12006 13838 12006 13838 0 Inst_W_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 12742 14076 12742 14076 0 Inst_W_IO_ConfigMem.ConfigBits\[59\]
rlabel metal1 11684 25738 11684 25738 0 Inst_W_IO_ConfigMem.ConfigBits\[60\]
rlabel metal2 12742 26044 12742 26044 0 Inst_W_IO_ConfigMem.ConfigBits\[61\]
rlabel metal1 7268 26894 7268 26894 0 Inst_W_IO_ConfigMem.ConfigBits\[62\]
rlabel metal1 7682 26554 7682 26554 0 Inst_W_IO_ConfigMem.ConfigBits\[63\]
rlabel metal1 5796 25398 5796 25398 0 Inst_W_IO_ConfigMem.ConfigBits\[64\]
rlabel metal1 7130 25330 7130 25330 0 Inst_W_IO_ConfigMem.ConfigBits\[65\]
rlabel metal1 11086 25432 11086 25432 0 Inst_W_IO_ConfigMem.ConfigBits\[66\]
rlabel metal1 13386 25330 13386 25330 0 Inst_W_IO_ConfigMem.ConfigBits\[67\]
rlabel metal1 7313 29070 7313 29070 0 Inst_W_IO_ConfigMem.ConfigBits\[68\]
rlabel metal1 7866 28730 7866 28730 0 Inst_W_IO_ConfigMem.ConfigBits\[69\]
rlabel metal2 12558 34357 12558 34357 0 Inst_W_IO_ConfigMem.ConfigBits\[70\]
rlabel metal1 12834 28186 12834 28186 0 Inst_W_IO_ConfigMem.ConfigBits\[71\]
rlabel metal1 13340 5338 13340 5338 0 Inst_W_IO_ConfigMem.ConfigBits\[72\]
rlabel metal2 13662 5831 13662 5831 0 Inst_W_IO_ConfigMem.ConfigBits\[73\]
rlabel metal2 12374 5066 12374 5066 0 Inst_W_IO_ConfigMem.ConfigBits\[74\]
rlabel metal1 13202 3706 13202 3706 0 Inst_W_IO_ConfigMem.ConfigBits\[75\]
rlabel metal1 8372 18190 8372 18190 0 Inst_W_IO_ConfigMem.ConfigBits\[76\]
rlabel metal2 9016 18258 9016 18258 0 Inst_W_IO_ConfigMem.ConfigBits\[77\]
rlabel metal2 12742 20162 12742 20162 0 Inst_W_IO_ConfigMem.ConfigBits\[78\]
rlabel metal2 13570 20604 13570 20604 0 Inst_W_IO_ConfigMem.ConfigBits\[79\]
rlabel metal1 8050 21862 8050 21862 0 Inst_W_IO_ConfigMem.ConfigBits\[80\]
rlabel metal1 8602 21114 8602 21114 0 Inst_W_IO_ConfigMem.ConfigBits\[81\]
rlabel metal1 8188 24650 8188 24650 0 Inst_W_IO_ConfigMem.ConfigBits\[82\]
rlabel metal2 9246 25228 9246 25228 0 Inst_W_IO_ConfigMem.ConfigBits\[83\]
rlabel metal1 6072 17034 6072 17034 0 Inst_W_IO_ConfigMem.ConfigBits\[84\]
rlabel metal2 6578 17170 6578 17170 0 Inst_W_IO_ConfigMem.ConfigBits\[85\]
rlabel metal1 12466 22168 12466 22168 0 Inst_W_IO_ConfigMem.ConfigBits\[86\]
rlabel metal1 12880 21658 12880 21658 0 Inst_W_IO_ConfigMem.ConfigBits\[87\]
rlabel metal2 9890 30634 9890 30634 0 Inst_W_IO_ConfigMem.ConfigBits\[88\]
rlabel metal2 10442 31212 10442 31212 0 Inst_W_IO_ConfigMem.ConfigBits\[89\]
rlabel metal1 8970 18700 8970 18700 0 Inst_W_IO_ConfigMem.ConfigBits\[8\]
rlabel metal1 12650 32198 12650 32198 0 Inst_W_IO_ConfigMem.ConfigBits\[90\]
rlabel metal1 12696 33286 12696 33286 0 Inst_W_IO_ConfigMem.ConfigBits\[91\]
rlabel metal2 9246 26945 9246 26945 0 Inst_W_IO_ConfigMem.ConfigBits\[92\]
rlabel metal2 9798 27132 9798 27132 0 Inst_W_IO_ConfigMem.ConfigBits\[93\]
rlabel metal1 10258 23834 10258 23834 0 Inst_W_IO_ConfigMem.ConfigBits\[94\]
rlabel metal2 10902 24412 10902 24412 0 Inst_W_IO_ConfigMem.ConfigBits\[95\]
rlabel metal1 9614 29784 9614 29784 0 Inst_W_IO_ConfigMem.ConfigBits\[96\]
rlabel metal2 9016 32198 9016 32198 0 Inst_W_IO_ConfigMem.ConfigBits\[97\]
rlabel metal2 12282 30430 12282 30430 0 Inst_W_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 13248 34034 13248 34034 0 Inst_W_IO_ConfigMem.ConfigBits\[99\]
rlabel metal1 5704 18734 5704 18734 0 Inst_W_IO_ConfigMem.ConfigBits\[9\]
rlabel metal2 10074 18649 10074 18649 0 Inst_W_IO_switch_matrix.E1BEG0
rlabel metal1 6578 18292 6578 18292 0 Inst_W_IO_switch_matrix.E1BEG1
rlabel metal1 14306 18836 14306 18836 0 Inst_W_IO_switch_matrix.E1BEG2
rlabel metal1 10994 18258 10994 18258 0 Inst_W_IO_switch_matrix.E1BEG3
rlabel metal2 8786 14144 8786 14144 0 Inst_W_IO_switch_matrix.E2BEG0
rlabel metal1 9614 16150 9614 16150 0 Inst_W_IO_switch_matrix.E2BEG1
rlabel metal1 12903 14382 12903 14382 0 Inst_W_IO_switch_matrix.E2BEG2
rlabel metal1 11638 16558 11638 16558 0 Inst_W_IO_switch_matrix.E2BEG3
rlabel metal2 13938 16116 13938 16116 0 Inst_W_IO_switch_matrix.E2BEG4
rlabel metal1 12558 16150 12558 16150 0 Inst_W_IO_switch_matrix.E2BEG5
rlabel metal1 11776 19482 11776 19482 0 Inst_W_IO_switch_matrix.E2BEG6
rlabel metal2 12006 18836 12006 18836 0 Inst_W_IO_switch_matrix.E2BEG7
rlabel metal1 12190 20910 12190 20910 0 Inst_W_IO_switch_matrix.E2BEGb0
rlabel metal2 13892 21998 13892 21998 0 Inst_W_IO_switch_matrix.E2BEGb1
rlabel metal2 9430 16592 9430 16592 0 Inst_W_IO_switch_matrix.E2BEGb2
rlabel metal1 12466 15096 12466 15096 0 Inst_W_IO_switch_matrix.E2BEGb3
rlabel metal1 13294 12104 13294 12104 0 Inst_W_IO_switch_matrix.E2BEGb4
rlabel metal1 14674 22066 14674 22066 0 Inst_W_IO_switch_matrix.E2BEGb5
rlabel metal1 15088 7514 15088 7514 0 Inst_W_IO_switch_matrix.E2BEGb6
rlabel metal3 14007 17204 14007 17204 0 Inst_W_IO_switch_matrix.E2BEGb7
rlabel metal1 12328 23086 12328 23086 0 Inst_W_IO_switch_matrix.E6BEG0
rlabel metal1 13432 20230 13432 20230 0 Inst_W_IO_switch_matrix.E6BEG1
rlabel metal1 10856 29818 10856 29818 0 Inst_W_IO_switch_matrix.E6BEG10
rlabel metal2 13478 30294 13478 30294 0 Inst_W_IO_switch_matrix.E6BEG11
rlabel metal2 12926 29002 12926 29002 0 Inst_W_IO_switch_matrix.E6BEG2
rlabel metal1 15042 31790 15042 31790 0 Inst_W_IO_switch_matrix.E6BEG3
rlabel via2 12926 29155 12926 29155 0 Inst_W_IO_switch_matrix.E6BEG4
rlabel metal1 12972 29070 12972 29070 0 Inst_W_IO_switch_matrix.E6BEG5
rlabel metal1 11546 29648 11546 29648 0 Inst_W_IO_switch_matrix.E6BEG6
rlabel metal1 13616 30362 13616 30362 0 Inst_W_IO_switch_matrix.E6BEG7
rlabel metal1 10764 27098 10764 27098 0 Inst_W_IO_switch_matrix.E6BEG8
rlabel metal1 11730 24378 11730 24378 0 Inst_W_IO_switch_matrix.E6BEG9
rlabel via2 8510 23035 8510 23035 0 Inst_W_IO_switch_matrix.EE4BEG0
rlabel metal1 13340 23086 13340 23086 0 Inst_W_IO_switch_matrix.EE4BEG1
rlabel metal2 12834 26741 12834 26741 0 Inst_W_IO_switch_matrix.EE4BEG10
rlabel metal1 12328 25126 12328 25126 0 Inst_W_IO_switch_matrix.EE4BEG11
rlabel metal1 12006 29172 12006 29172 0 Inst_W_IO_switch_matrix.EE4BEG12
rlabel metal1 13708 28730 13708 28730 0 Inst_W_IO_switch_matrix.EE4BEG13
rlabel metal2 13938 6681 13938 6681 0 Inst_W_IO_switch_matrix.EE4BEG14
rlabel metal1 14076 6426 14076 6426 0 Inst_W_IO_switch_matrix.EE4BEG15
rlabel metal2 13432 32300 13432 32300 0 Inst_W_IO_switch_matrix.EE4BEG2
rlabel metal2 12374 27914 12374 27914 0 Inst_W_IO_switch_matrix.EE4BEG3
rlabel metal1 11086 12104 11086 12104 0 Inst_W_IO_switch_matrix.EE4BEG4
rlabel metal2 13800 21828 13800 21828 0 Inst_W_IO_switch_matrix.EE4BEG5
rlabel metal1 14076 16694 14076 16694 0 Inst_W_IO_switch_matrix.EE4BEG6
rlabel metal1 13524 13974 13524 13974 0 Inst_W_IO_switch_matrix.EE4BEG7
rlabel metal1 12926 26010 12926 26010 0 Inst_W_IO_switch_matrix.EE4BEG8
rlabel metal2 9706 27234 9706 27234 0 Inst_W_IO_switch_matrix.EE4BEG9
rlabel metal1 11684 5542 11684 5542 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out0
rlabel metal1 11546 8500 11546 8500 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out1
rlabel via1 12570 8466 12570 8466 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out2
rlabel metal1 12466 8432 12466 8432 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_A_I.cus_mux41_buf_out3
rlabel metal1 11914 5780 11914 5780 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out0
rlabel metal1 11638 5678 11638 5678 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out1
rlabel via1 12754 5746 12754 5746 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out2
rlabel metal1 12466 5780 12466 5780 0 Inst_W_IO_switch_matrix.inst_cus_mux161_buf_B_I.cus_mux41_buf_out3
rlabel metal1 10534 18258 10534 18258 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN\[0\]
rlabel metal1 9108 18734 9108 18734 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0.AIN\[1\]
rlabel metal1 9844 18394 9844 18394 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._0_
rlabel metal1 9522 18836 9522 18836 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG0._1_
rlabel metal1 5888 18258 5888 18258 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN\[0\]
rlabel metal1 5892 19336 5892 19336 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1.AIN\[1\]
rlabel metal2 5842 18564 5842 18564 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._0_
rlabel metal1 5888 18802 5888 18802 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG1._1_
rlabel metal1 6578 19958 6578 19958 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN\[0\]
rlabel metal1 6854 19788 6854 19788 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2.AIN\[1\]
rlabel metal1 6394 20230 6394 20230 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._0_
rlabel metal1 6808 20026 6808 20026 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG2._1_
rlabel metal1 10718 20434 10718 20434 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN\[0\]
rlabel metal2 9706 21012 9706 21012 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3.AIN\[1\]
rlabel metal1 10258 20570 10258 20570 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._0_
rlabel metal1 9706 21050 9706 21050 0 Inst_W_IO_switch_matrix.inst_cus_mux21_E1BEG3._1_
rlabel metal1 9706 7514 9706 7514 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A0
rlabel metal1 6854 7786 6854 7786 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.A1
rlabel metal1 6578 8058 6578 8058 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN\[0\]
rlabel metal1 6946 7990 6946 7990 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst.AIN\[1\]
rlabel metal1 6670 8330 6670 8330 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._0_
rlabel metal1 6900 8398 6900 8398 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_A_T.cus_mux21_inst._1_
rlabel metal1 8188 9350 8188 9350 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A0
rlabel metal1 6670 9554 6670 9554 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.A1
rlabel metal1 5382 10030 5382 10030 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN\[0\]
rlabel metal1 5796 9690 5796 9690 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst.AIN\[1\]
rlabel metal1 5290 9554 5290 9554 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._0_
rlabel metal1 5336 9486 5336 9486 0 Inst_W_IO_switch_matrix.inst_cus_mux81_buf_B_T.cus_mux21_inst._1_
rlabel metal2 598 9136 598 9136 0 UserCLK
rlabel metal1 1656 43418 1656 43418 0 UserCLKo
rlabel metal3 15096 4964 15096 4964 0 W1END[0]
rlabel metal3 15165 5236 15165 5236 0 W1END[1]
rlabel metal3 15510 5508 15510 5508 0 W1END[2]
rlabel metal3 15372 5780 15372 5780 0 W1END[3]
rlabel metal3 15096 8228 15096 8228 0 W2END[0]
rlabel metal3 14912 8500 14912 8500 0 W2END[1]
rlabel metal3 15510 8772 15510 8772 0 W2END[2]
rlabel metal3 15142 9044 15142 9044 0 W2END[3]
rlabel metal1 13110 8908 13110 8908 0 W2END[4]
rlabel metal3 14314 9588 14314 9588 0 W2END[5]
rlabel metal3 15510 9860 15510 9860 0 W2END[6]
rlabel metal3 14820 10132 14820 10132 0 W2END[7]
rlabel metal3 15050 6052 15050 6052 0 W2MID[0]
rlabel metal3 15625 6324 15625 6324 0 W2MID[1]
rlabel metal1 13708 5202 13708 5202 0 W2MID[2]
rlabel metal3 15510 6868 15510 6868 0 W2MID[3]
rlabel metal3 15096 7140 15096 7140 0 W2MID[4]
rlabel metal3 15234 7412 15234 7412 0 W2MID[5]
rlabel metal3 15533 7684 15533 7684 0 W2MID[6]
rlabel metal3 15096 7956 15096 7956 0 W2MID[7]
rlabel metal3 15372 14756 15372 14756 0 W6END[0]
rlabel metal3 15510 17476 15510 17476 0 W6END[10]
rlabel metal2 11454 17663 11454 17663 0 W6END[11]
rlabel metal3 15096 15028 15096 15028 0 W6END[1]
rlabel metal3 15510 15300 15510 15300 0 W6END[2]
rlabel metal3 15372 15572 15372 15572 0 W6END[3]
rlabel metal3 14820 15844 14820 15844 0 W6END[4]
rlabel metal3 14728 16116 14728 16116 0 W6END[5]
rlabel metal3 15510 16388 15510 16388 0 W6END[6]
rlabel metal3 15096 16660 15096 16660 0 W6END[7]
rlabel metal3 14866 16932 14866 16932 0 W6END[8]
rlabel metal3 15096 17204 15096 17204 0 W6END[9]
rlabel metal3 15280 10404 15280 10404 0 WW4END[0]
rlabel metal3 15556 13124 15556 13124 0 WW4END[10]
rlabel metal3 14912 13396 14912 13396 0 WW4END[11]
rlabel metal3 14958 13668 14958 13668 0 WW4END[12]
rlabel metal3 15533 13940 15533 13940 0 WW4END[13]
rlabel metal3 15510 14212 15510 14212 0 WW4END[14]
rlabel metal3 15050 14484 15050 14484 0 WW4END[15]
rlabel metal3 15050 10676 15050 10676 0 WW4END[1]
rlabel metal3 15556 10948 15556 10948 0 WW4END[2]
rlabel metal3 14130 11220 14130 11220 0 WW4END[3]
rlabel metal3 15096 11492 15096 11492 0 WW4END[4]
rlabel metal3 15004 11764 15004 11764 0 WW4END[5]
rlabel metal3 15533 12036 15533 12036 0 WW4END[6]
rlabel metal2 11822 12563 11822 12563 0 WW4END[7]
rlabel metal3 14981 12580 14981 12580 0 WW4END[8]
rlabel metal3 15188 12852 15188 12852 0 WW4END[9]
rlabel metal1 9338 30090 9338 30090 0 data_inbuf_0.X
rlabel metal1 11178 30668 11178 30668 0 data_inbuf_1.X
rlabel metal1 10350 33082 10350 33082 0 data_inbuf_10.X
rlabel metal2 12650 34085 12650 34085 0 data_inbuf_11.X
rlabel metal2 9614 33796 9614 33796 0 data_inbuf_12.X
rlabel metal2 9890 33762 9890 33762 0 data_inbuf_13.X
rlabel metal1 8786 33626 8786 33626 0 data_inbuf_14.X
rlabel metal1 9476 34102 9476 34102 0 data_inbuf_15.X
rlabel metal1 11868 34714 11868 34714 0 data_inbuf_16.X
rlabel metal1 12650 34476 12650 34476 0 data_inbuf_17.X
rlabel metal1 9246 34714 9246 34714 0 data_inbuf_18.X
rlabel metal1 9062 34544 9062 34544 0 data_inbuf_19.X
rlabel metal1 12282 30804 12282 30804 0 data_inbuf_2.X
rlabel metal1 12650 36006 12650 36006 0 data_inbuf_20.X
rlabel metal1 11822 36652 11822 36652 0 data_inbuf_21.X
rlabel metal1 13110 36550 13110 36550 0 data_inbuf_22.X
rlabel metal1 12558 36856 12558 36856 0 data_inbuf_23.X
rlabel metal2 12742 37519 12742 37519 0 data_inbuf_24.X
rlabel metal1 12650 37366 12650 37366 0 data_inbuf_25.X
rlabel metal1 10488 36890 10488 36890 0 data_inbuf_26.X
rlabel metal1 11638 37434 11638 37434 0 data_inbuf_27.X
rlabel metal1 12972 38522 12972 38522 0 data_inbuf_28.X
rlabel metal1 12236 38930 12236 38930 0 data_inbuf_29.X
rlabel metal2 13110 32402 13110 32402 0 data_inbuf_3.X
rlabel metal1 8326 39440 8326 39440 0 data_inbuf_30.X
rlabel metal1 9430 39372 9430 39372 0 data_inbuf_31.X
rlabel metal1 12558 31994 12558 31994 0 data_inbuf_4.X
rlabel metal2 13294 32963 13294 32963 0 data_inbuf_5.X
rlabel metal1 12558 33864 12558 33864 0 data_inbuf_6.X
rlabel metal1 12190 32912 12190 32912 0 data_inbuf_7.X
rlabel metal1 11086 32912 11086 32912 0 data_inbuf_8.X
rlabel metal1 12558 34612 12558 34612 0 data_inbuf_9.X
rlabel metal1 10534 30736 10534 30736 0 data_outbuf_0.X
rlabel metal1 11086 30906 11086 30906 0 data_outbuf_1.X
rlabel metal1 11178 33524 11178 33524 0 data_outbuf_10.X
rlabel metal1 13386 35122 13386 35122 0 data_outbuf_11.X
rlabel metal1 10994 34000 10994 34000 0 data_outbuf_12.X
rlabel metal1 10672 34170 10672 34170 0 data_outbuf_13.X
rlabel metal1 9292 34170 9292 34170 0 data_outbuf_14.X
rlabel metal1 10718 34612 10718 34612 0 data_outbuf_15.X
rlabel metal1 12236 35054 12236 35054 0 data_outbuf_16.X
rlabel metal1 13110 36176 13110 36176 0 data_outbuf_17.X
rlabel metal1 9982 35258 9982 35258 0 data_outbuf_18.X
rlabel metal1 10258 35190 10258 35190 0 data_outbuf_19.X
rlabel metal1 12650 32878 12650 32878 0 data_outbuf_2.X
rlabel metal1 12420 36142 12420 36142 0 data_outbuf_20.X
rlabel metal2 11638 37604 11638 37604 0 data_outbuf_21.X
rlabel metal1 12834 37808 12834 37808 0 data_outbuf_22.X
rlabel metal2 11914 37060 11914 37060 0 data_outbuf_23.X
rlabel metal1 13064 37978 13064 37978 0 data_outbuf_24.X
rlabel metal2 12558 38131 12558 38131 0 data_outbuf_25.X
rlabel metal2 10810 37638 10810 37638 0 data_outbuf_26.X
rlabel metal2 12466 38182 12466 38182 0 data_outbuf_27.X
rlabel metal1 13064 39406 13064 39406 0 data_outbuf_28.X
rlabel metal2 12742 39236 12742 39236 0 data_outbuf_29.X
rlabel via1 12558 31875 12558 31875 0 data_outbuf_3.X
rlabel metal1 9154 39474 9154 39474 0 data_outbuf_30.X
rlabel metal1 9706 39440 9706 39440 0 data_outbuf_31.X
rlabel metal1 12098 31824 12098 31824 0 data_outbuf_4.X
rlabel metal1 13386 34102 13386 34102 0 data_outbuf_5.X
rlabel metal1 12926 34578 12926 34578 0 data_outbuf_6.X
rlabel metal1 12466 32912 12466 32912 0 data_outbuf_7.X
rlabel metal1 10994 33082 10994 33082 0 data_outbuf_8.X
rlabel metal2 12466 35020 12466 35020 0 data_outbuf_9.X
rlabel metal1 2070 9656 2070 9656 0 net1
rlabel metal1 1885 14994 1885 14994 0 net10
rlabel metal1 6946 14892 6946 14892 0 net100
rlabel metal1 15364 20026 15364 20026 0 net101
rlabel metal1 13846 13838 13846 13838 0 net102
rlabel metal1 1748 10778 1748 10778 0 net103
rlabel metal1 1610 9690 1610 9690 0 net104
rlabel metal1 1794 12138 1794 12138 0 net105
rlabel metal1 2116 12410 2116 12410 0 net106
rlabel metal1 2254 13974 2254 13974 0 net107
rlabel metal1 1932 14314 1932 14314 0 net108
rlabel metal1 1794 4590 1794 4590 0 net109
rlabel metal1 2115 15470 2115 15470 0 net11
rlabel metal1 1978 5270 1978 5270 0 net110
rlabel metal1 1702 6358 1702 6358 0 net111
rlabel metal1 1518 7480 1518 7480 0 net112
rlabel metal1 1932 8534 1932 8534 0 net113
rlabel metal1 1840 7854 1840 7854 0 net114
rlabel metal1 12926 17646 12926 17646 0 net115
rlabel metal2 13662 17119 13662 17119 0 net116
rlabel metal1 14168 17646 14168 17646 0 net117
rlabel metal1 12788 19346 12788 19346 0 net118
rlabel metal1 14260 13498 14260 13498 0 net119
rlabel metal1 1702 5595 1702 5595 0 net12
rlabel metal1 10442 17850 10442 17850 0 net120
rlabel metal1 13616 14586 13616 14586 0 net121
rlabel metal1 11960 16762 11960 16762 0 net122
rlabel metal1 13708 18870 13708 18870 0 net123
rlabel metal1 13754 19312 13754 19312 0 net124
rlabel metal1 13984 18326 13984 18326 0 net125
rlabel metal2 13386 21046 13386 21046 0 net126
rlabel metal1 14214 20808 14214 20808 0 net127
rlabel metal1 13432 21862 13432 21862 0 net128
rlabel metal1 14214 21012 14214 21012 0 net129
rlabel metal2 1610 31008 1610 31008 0 net13
rlabel metal1 14214 20570 14214 20570 0 net130
rlabel metal1 14950 12342 14950 12342 0 net131
rlabel metal1 14122 21998 14122 21998 0 net132
rlabel metal1 13478 22746 13478 22746 0 net133
rlabel metal1 13938 22474 13938 22474 0 net134
rlabel metal1 12650 26928 12650 26928 0 net135
rlabel metal1 13432 30702 13432 30702 0 net136
rlabel metal2 11546 30991 11546 30991 0 net137
rlabel metal1 12742 27642 12742 27642 0 net138
rlabel metal1 13386 29240 13386 29240 0 net139
rlabel metal1 1702 16728 1702 16728 0 net14
rlabel metal2 14214 30430 14214 30430 0 net140
rlabel metal2 12742 29920 12742 29920 0 net141
rlabel metal1 13248 29002 13248 29002 0 net142
rlabel metal1 11776 29818 11776 29818 0 net143
rlabel metal2 14352 32300 14352 32300 0 net144
rlabel metal1 11684 29478 11684 29478 0 net145
rlabel metal1 12834 29240 12834 29240 0 net146
rlabel metal1 13570 23290 13570 23290 0 net147
rlabel metal1 13018 27064 13018 27064 0 net148
rlabel metal1 14214 27506 14214 27506 0 net149
rlabel metal1 1655 10030 1655 10030 0 net15
rlabel metal1 13340 26962 13340 26962 0 net150
rlabel metal1 13846 27438 13846 27438 0 net151
rlabel metal2 12558 27591 12558 27591 0 net152
rlabel metal2 13938 28798 13938 28798 0 net153
rlabel metal1 13386 23222 13386 23222 0 net154
rlabel metal1 14398 33014 14398 33014 0 net155
rlabel metal1 13984 25262 13984 25262 0 net156
rlabel metal1 13938 24718 13938 24718 0 net157
rlabel metal1 13294 24310 13294 24310 0 net158
rlabel metal1 13984 26350 13984 26350 0 net159
rlabel metal1 1647 8912 1647 8912 0 net16
rlabel metal1 13018 24616 13018 24616 0 net160
rlabel metal1 14122 26894 14122 26894 0 net161
rlabel metal1 12558 27030 12558 27030 0 net162
rlabel metal2 10350 31127 10350 31127 0 net163
rlabel metal2 13478 34000 13478 34000 0 net164
rlabel metal1 13938 34680 13938 34680 0 net165
rlabel metal1 12834 33932 12834 33932 0 net166
rlabel via2 13570 35003 13570 35003 0 net167
rlabel metal1 9338 34476 9338 34476 0 net168
rlabel metal1 13570 35598 13570 35598 0 net169
rlabel metal2 6486 34068 6486 34068 0 net17
rlabel metal2 13662 35972 13662 35972 0 net170
rlabel metal1 13248 36074 13248 36074 0 net171
rlabel metal2 13478 35938 13478 35938 0 net172
rlabel metal1 12742 36108 12742 36108 0 net173
rlabel metal2 13754 32147 13754 32147 0 net174
rlabel metal2 12190 36754 12190 36754 0 net175
rlabel metal2 13570 37400 13570 37400 0 net176
rlabel metal1 13110 37910 13110 37910 0 net177
rlabel metal1 13938 37774 13938 37774 0 net178
rlabel metal1 14214 38352 14214 38352 0 net179
rlabel metal1 1610 34680 1610 34680 0 net18
rlabel metal1 13662 38284 13662 38284 0 net180
rlabel metal1 13432 38930 13432 38930 0 net181
rlabel metal1 13386 38998 13386 38998 0 net182
rlabel metal1 14214 39338 14214 39338 0 net183
rlabel metal1 13064 39338 13064 39338 0 net184
rlabel metal1 13202 32810 13202 32810 0 net185
rlabel metal2 13386 39814 13386 39814 0 net186
rlabel metal1 13938 39984 13938 39984 0 net187
rlabel metal2 12190 32198 12190 32198 0 net188
rlabel metal1 12926 31960 12926 31960 0 net189
rlabel metal2 5796 18836 5796 18836 0 net19
rlabel metal2 14122 33898 14122 33898 0 net190
rlabel metal1 13340 33490 13340 33490 0 net191
rlabel metal1 13018 33082 13018 33082 0 net192
rlabel metal1 14214 34068 14214 34068 0 net193
rlabel metal1 13478 33966 13478 33966 0 net194
rlabel metal1 1656 43282 1656 43282 0 net195
rlabel metal1 8786 42874 8786 42874 0 net196
rlabel metal2 9338 43078 9338 43078 0 net197
rlabel metal1 10166 42874 10166 42874 0 net198
rlabel metal1 11224 42874 11224 42874 0 net199
rlabel metal1 4492 20842 4492 20842 0 net2
rlabel via2 12834 37213 12834 37213 0 net20
rlabel metal1 11822 42806 11822 42806 0 net200
rlabel metal2 12558 43078 12558 43078 0 net201
rlabel metal1 13156 42874 13156 42874 0 net202
rlabel metal1 14214 42874 14214 42874 0 net203
rlabel metal1 13202 42806 13202 42806 0 net204
rlabel metal1 13800 42330 13800 42330 0 net205
rlabel metal1 2116 42874 2116 42874 0 net206
rlabel metal1 2944 42874 2944 42874 0 net207
rlabel metal1 3588 42874 3588 42874 0 net208
rlabel metal1 4278 42874 4278 42874 0 net209
rlabel metal1 2185 36550 2185 36550 0 net21
rlabel metal1 5060 39066 5060 39066 0 net210
rlabel metal1 5796 42874 5796 42874 0 net211
rlabel metal1 6532 42874 6532 42874 0 net212
rlabel metal1 7222 42874 7222 42874 0 net213
rlabel metal1 7958 42874 7958 42874 0 net214
rlabel metal2 2622 22100 2622 22100 0 net215
rlabel via1 7970 7922 7970 7922 0 net216
rlabel metal1 8579 10098 8579 10098 0 net217
rlabel metal1 7774 7922 7774 7922 0 net218
rlabel metal2 7866 10336 7866 10336 0 net219
rlabel viali 6753 14352 6753 14352 0 net22
rlabel metal1 1610 38216 1610 38216 0 net23
rlabel metal1 12558 38896 12558 38896 0 net24
rlabel via3 15387 21964 15387 21964 0 net25
rlabel via1 6669 13906 6669 13906 0 net26
rlabel metal1 7589 20910 7589 20910 0 net27
rlabel metal1 2116 18122 2116 18122 0 net28
rlabel via3 12627 31756 12627 31756 0 net29
rlabel metal1 9659 16082 9659 16082 0 net3
rlabel metal2 12742 14943 12742 14943 0 net30
rlabel metal1 1702 20468 1702 20468 0 net31
rlabel metal1 9982 22066 9982 22066 0 net32
rlabel metal3 10925 21964 10925 21964 0 net33
rlabel metal2 1610 22848 1610 22848 0 net34
rlabel metal2 2254 1122 2254 1122 0 net35
rlabel metal1 8786 1530 8786 1530 0 net36
rlabel metal1 9430 1530 9430 1530 0 net37
rlabel metal1 10166 1530 10166 1530 0 net38
rlabel metal1 10902 1530 10902 1530 0 net39
rlabel metal1 1702 23732 1702 23732 0 net4
rlabel metal1 11684 1530 11684 1530 0 net40
rlabel metal1 12374 1530 12374 1530 0 net41
rlabel metal1 13248 1530 13248 1530 0 net42
rlabel metal2 13754 1734 13754 1734 0 net43
rlabel metal2 13478 1768 13478 1768 0 net44
rlabel metal1 13570 1258 13570 1258 0 net45
rlabel metal1 4945 1870 4945 1870 0 net46
rlabel metal1 5014 1224 5014 1224 0 net47
rlabel metal1 1518 5678 1518 5678 0 net48
rlabel metal1 4324 1530 4324 1530 0 net49
rlabel metal2 11132 32300 11132 32300 0 net5
rlabel metal1 5060 1530 5060 1530 0 net50
rlabel metal1 5796 1530 5796 1530 0 net51
rlabel metal1 6532 1530 6532 1530 0 net52
rlabel metal1 7222 1530 7222 1530 0 net53
rlabel metal1 7958 1530 7958 1530 0 net54
rlabel metal2 14398 3859 14398 3859 0 net55
rlabel metal2 14398 6035 14398 6035 0 net56
rlabel metal1 11224 5338 11224 5338 0 net57
rlabel metal1 12558 20332 12558 20332 0 net58
rlabel metal1 9614 7990 9614 7990 0 net59
rlabel metal1 1702 25398 1702 25398 0 net6
rlabel metal1 9430 7820 9430 7820 0 net60
rlabel via1 10454 7854 10454 7854 0 net61
rlabel metal1 7084 7922 7084 7922 0 net62
rlabel metal2 9798 14790 9798 14790 0 net63
rlabel metal1 7314 10098 7314 10098 0 net64
rlabel metal2 6302 21318 6302 21318 0 net65
rlabel metal1 10074 8398 10074 8398 0 net66
rlabel metal1 13202 6630 13202 6630 0 net67
rlabel metal2 9936 19346 9936 19346 0 net68
rlabel metal1 13662 6766 13662 6766 0 net69
rlabel metal1 8556 33354 8556 33354 0 net7
rlabel metal1 13064 6290 13064 6290 0 net70
rlabel metal1 9246 17102 9246 17102 0 net71
rlabel metal1 8786 6256 8786 6256 0 net72
rlabel metal2 7866 16167 7866 16167 0 net73
rlabel metal2 8142 7106 8142 7106 0 net74
rlabel metal2 12650 22865 12650 22865 0 net75
rlabel via1 13398 20366 13398 20366 0 net76
rlabel via1 10718 18343 10718 18343 0 net77
rlabel metal1 14030 14518 14030 14518 0 net78
rlabel metal1 5658 23018 5658 23018 0 net79
rlabel metal1 1748 26758 1748 26758 0 net8
rlabel metal1 6670 26826 6670 26826 0 net80
rlabel metal2 10304 21012 10304 21012 0 net81
rlabel metal1 13110 17000 13110 17000 0 net82
rlabel metal1 13202 15640 13202 15640 0 net83
rlabel metal1 7866 14348 7866 14348 0 net84
rlabel metal1 13041 30158 13041 30158 0 net85
rlabel metal1 14352 17510 14352 17510 0 net86
rlabel metal2 11638 12070 11638 12070 0 net87
rlabel metal2 13708 19822 13708 19822 0 net88
rlabel metal1 7832 12274 7832 12274 0 net89
rlabel metal1 1656 27846 1656 27846 0 net9
rlabel metal1 10350 24038 10350 24038 0 net90
rlabel metal1 13662 11118 13662 11118 0 net91
rlabel metal2 14490 13090 14490 13090 0 net92
rlabel via1 11247 20910 11247 20910 0 net93
rlabel metal3 9039 29036 9039 29036 0 net94
rlabel metal2 11822 21369 11822 21369 0 net95
rlabel metal2 6762 14994 6762 14994 0 net96
rlabel metal1 13984 8806 13984 8806 0 net97
rlabel metal2 13938 12019 13938 12019 0 net98
rlabel metal2 15318 13855 15318 13855 0 net99
rlabel metal1 1794 34170 1794 34170 0 strobe_inbuf_0.X
rlabel metal1 2208 36890 2208 36890 0 strobe_inbuf_1.X
rlabel metal1 5382 14586 5382 14586 0 strobe_inbuf_10.X
rlabel metal2 2392 38998 2392 38998 0 strobe_inbuf_11.X
rlabel metal1 7774 1836 7774 1836 0 strobe_inbuf_12.X
rlabel metal2 10902 2363 10902 2363 0 strobe_inbuf_13.X
rlabel metal2 11730 1785 11730 1785 0 strobe_inbuf_14.X
rlabel metal2 12466 41871 12466 41871 0 strobe_inbuf_15.X
rlabel metal1 13248 2074 13248 2074 0 strobe_inbuf_16.X
rlabel metal1 14490 1938 14490 1938 0 strobe_inbuf_17.X
rlabel metal1 14996 2074 14996 2074 0 strobe_inbuf_18.X
rlabel metal1 14950 1258 14950 1258 0 strobe_inbuf_19.X
rlabel metal1 2990 41786 2990 41786 0 strobe_inbuf_2.X
rlabel metal1 3220 21658 3220 21658 0 strobe_inbuf_3.X
rlabel metal2 4094 2210 4094 2210 0 strobe_inbuf_4.X
rlabel metal1 3680 2006 3680 2006 0 strobe_inbuf_5.X
rlabel via3 5819 2652 5819 2652 0 strobe_inbuf_6.X
rlabel metal1 6624 2074 6624 2074 0 strobe_inbuf_7.X
rlabel metal2 7222 2417 7222 2417 0 strobe_inbuf_8.X
rlabel metal3 7567 2652 7567 2652 0 strobe_inbuf_9.X
rlabel metal1 1886 34714 1886 34714 0 strobe_outbuf_0.X
rlabel metal1 2162 42330 2162 42330 0 strobe_outbuf_1.X
rlabel metal1 8740 42330 8740 42330 0 strobe_outbuf_10.X
rlabel metal1 9430 42330 9430 42330 0 strobe_outbuf_11.X
rlabel metal1 10212 42330 10212 42330 0 strobe_outbuf_12.X
rlabel metal1 10902 42330 10902 42330 0 strobe_outbuf_13.X
rlabel metal1 11638 42330 11638 42330 0 strobe_outbuf_14.X
rlabel metal2 12466 42500 12466 42500 0 strobe_outbuf_15.X
rlabel metal1 13064 42330 13064 42330 0 strobe_outbuf_16.X
rlabel metal1 13938 42058 13938 42058 0 strobe_outbuf_17.X
rlabel metal2 14306 42432 14306 42432 0 strobe_outbuf_18.X
rlabel metal1 14260 41786 14260 41786 0 strobe_outbuf_19.X
rlabel metal1 2944 42330 2944 42330 0 strobe_outbuf_2.X
rlabel metal2 3358 21971 3358 21971 0 strobe_outbuf_3.X
rlabel metal1 2852 2618 2852 2618 0 strobe_outbuf_4.X
rlabel metal1 5014 38522 5014 38522 0 strobe_outbuf_5.X
rlabel metal1 5750 42330 5750 42330 0 strobe_outbuf_6.X
rlabel metal1 6532 42330 6532 42330 0 strobe_outbuf_7.X
rlabel metal1 7222 42330 7222 42330 0 strobe_outbuf_8.X
rlabel metal1 8096 42330 8096 42330 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 16000 44623
<< end >>
