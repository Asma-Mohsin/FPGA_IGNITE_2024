VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO S_term_single
  CLASS BLOCK ;
  FOREIGN S_term_single ;
  ORIGIN 0.000 0.000 ;
  SIZE 231.000 BY 182.000 ;
  PIN Co
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.260 181.300 95.640 182.000 ;
    END
  END Co
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 5.560 0.000 5.940 0.700 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 42.820 0.000 43.200 0.700 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 46.500 0.000 46.880 0.700 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 50.180 0.000 50.560 0.700 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 53.860 0.000 54.240 0.700 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 57.540 0.000 57.920 0.700 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.220 0.000 61.600 0.700 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 64.900 0.000 65.280 0.700 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 68.580 0.000 68.960 0.700 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 72.720 0.000 73.100 0.700 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 76.400 0.000 76.780 0.700 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.240 0.000 9.620 0.700 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 12.920 0.000 13.300 0.700 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 16.600 0.000 16.980 0.700 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.280 0.000 20.660 0.700 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 23.960 0.000 24.340 0.700 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 27.640 0.000 28.020 0.700 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 31.780 0.000 32.160 0.700 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.460 0.000 35.840 0.700 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 39.140 0.000 39.520 0.700 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 188.180 181.300 188.560 182.000 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.120 181.300 206.500 182.000 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 207.960 181.300 208.340 182.000 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 209.340 181.300 209.720 182.000 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 211.180 181.300 211.560 182.000 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 213.020 181.300 213.400 182.000 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 214.860 181.300 215.240 182.000 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 216.700 181.300 217.080 182.000 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 218.080 181.300 218.460 182.000 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 219.920 181.300 220.300 182.000 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 221.760 181.300 222.140 182.000 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.020 181.300 190.400 182.000 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 191.860 181.300 192.240 182.000 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.700 181.300 194.080 182.000 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 195.540 181.300 195.920 182.000 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 197.380 181.300 197.760 182.000 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 198.760 181.300 199.140 182.000 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 200.600 181.300 200.980 182.000 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 202.440 181.300 202.820 182.000 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 204.280 181.300 204.660 182.000 ;
    END
  END FrameStrobe_O[9]
  PIN N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 3.720 181.300 4.100 182.000 ;
    END
  END N1BEG[0]
  PIN N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 5.560 181.300 5.940 182.000 ;
    END
  END N1BEG[1]
  PIN N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 6.940 181.300 7.320 182.000 ;
    END
  END N1BEG[2]
  PIN N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 8.780 181.300 9.160 182.000 ;
    END
  END N1BEG[3]
  PIN N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 10.620 181.300 11.000 182.000 ;
    END
  END N2BEG[0]
  PIN N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 12.460 181.300 12.840 182.000 ;
    END
  END N2BEG[1]
  PIN N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 14.300 181.300 14.680 182.000 ;
    END
  END N2BEG[2]
  PIN N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 15.680 181.300 16.060 182.000 ;
    END
  END N2BEG[3]
  PIN N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 17.520 181.300 17.900 182.000 ;
    END
  END N2BEG[4]
  PIN N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.360 181.300 19.740 182.000 ;
    END
  END N2BEG[5]
  PIN N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 21.200 181.300 21.580 182.000 ;
    END
  END N2BEG[6]
  PIN N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 23.040 181.300 23.420 182.000 ;
    END
  END N2BEG[7]
  PIN N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 24.880 181.300 25.260 182.000 ;
    END
  END N2BEGb[0]
  PIN N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 26.260 181.300 26.640 182.000 ;
    END
  END N2BEGb[1]
  PIN N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 28.100 181.300 28.480 182.000 ;
    END
  END N2BEGb[2]
  PIN N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.940 181.300 30.320 182.000 ;
    END
  END N2BEGb[3]
  PIN N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 31.780 181.300 32.160 182.000 ;
    END
  END N2BEGb[4]
  PIN N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 33.620 181.300 34.000 182.000 ;
    END
  END N2BEGb[5]
  PIN N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.460 181.300 35.840 182.000 ;
    END
  END N2BEGb[6]
  PIN N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 36.840 181.300 37.220 182.000 ;
    END
  END N2BEGb[7]
  PIN N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.680 181.300 39.060 182.000 ;
    END
  END N4BEG[0]
  PIN N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 56.160 181.300 56.540 182.000 ;
    END
  END N4BEG[10]
  PIN N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.000 181.300 58.380 182.000 ;
    END
  END N4BEG[11]
  PIN N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 59.840 181.300 60.220 182.000 ;
    END
  END N4BEG[12]
  PIN N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.680 181.300 62.060 182.000 ;
    END
  END N4BEG[13]
  PIN N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.520 181.300 63.900 182.000 ;
    END
  END N4BEG[14]
  PIN N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 65.360 181.300 65.740 182.000 ;
    END
  END N4BEG[15]
  PIN N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 40.520 181.300 40.900 182.000 ;
    END
  END N4BEG[1]
  PIN N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 42.360 181.300 42.740 182.000 ;
    END
  END N4BEG[2]
  PIN N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 44.200 181.300 44.580 182.000 ;
    END
  END N4BEG[3]
  PIN N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 46.040 181.300 46.420 182.000 ;
    END
  END N4BEG[4]
  PIN N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.420 181.300 47.800 182.000 ;
    END
  END N4BEG[5]
  PIN N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 49.260 181.300 49.640 182.000 ;
    END
  END N4BEG[6]
  PIN N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 51.100 181.300 51.480 182.000 ;
    END
  END N4BEG[7]
  PIN N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.940 181.300 53.320 182.000 ;
    END
  END N4BEG[8]
  PIN N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.780 181.300 55.160 182.000 ;
    END
  END N4BEG[9]
  PIN NN4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 66.740 181.300 67.120 182.000 ;
    END
  END NN4BEG[0]
  PIN NN4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 84.680 181.300 85.060 182.000 ;
    END
  END NN4BEG[10]
  PIN NN4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 86.520 181.300 86.900 182.000 ;
    END
  END NN4BEG[11]
  PIN NN4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.900 181.300 88.280 182.000 ;
    END
  END NN4BEG[12]
  PIN NN4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 89.740 181.300 90.120 182.000 ;
    END
  END NN4BEG[13]
  PIN NN4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.580 181.300 91.960 182.000 ;
    END
  END NN4BEG[14]
  PIN NN4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.420 181.300 93.800 182.000 ;
    END
  END NN4BEG[15]
  PIN NN4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 68.580 181.300 68.960 182.000 ;
    END
  END NN4BEG[1]
  PIN NN4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.420 181.300 70.800 182.000 ;
    END
  END NN4BEG[2]
  PIN NN4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 72.260 181.300 72.640 182.000 ;
    END
  END NN4BEG[3]
  PIN NN4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.100 181.300 74.480 182.000 ;
    END
  END NN4BEG[4]
  PIN NN4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 75.940 181.300 76.320 182.000 ;
    END
  END NN4BEG[5]
  PIN NN4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.320 181.300 77.700 182.000 ;
    END
  END NN4BEG[6]
  PIN NN4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 79.160 181.300 79.540 182.000 ;
    END
  END NN4BEG[7]
  PIN NN4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 81.000 181.300 81.380 182.000 ;
    END
  END NN4BEG[8]
  PIN NN4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 82.840 181.300 83.220 182.000 ;
    END
  END NN4BEG[9]
  PIN S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 96.640 181.300 97.020 182.000 ;
    END
  END S1END[0]
  PIN S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 98.480 181.300 98.860 182.000 ;
    END
  END S1END[1]
  PIN S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 100.320 181.300 100.700 182.000 ;
    END
  END S1END[2]
  PIN S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 102.160 181.300 102.540 182.000 ;
    END
  END S1END[3]
  PIN S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 117.800 181.300 118.180 182.000 ;
    END
  END S2END[0]
  PIN S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 119.640 181.300 120.020 182.000 ;
    END
  END S2END[1]
  PIN S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 121.480 181.300 121.860 182.000 ;
    END
  END S2END[2]
  PIN S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 123.320 181.300 123.700 182.000 ;
    END
  END S2END[3]
  PIN S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 125.160 181.300 125.540 182.000 ;
    END
  END S2END[4]
  PIN S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 127.000 181.300 127.380 182.000 ;
    END
  END S2END[5]
  PIN S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 128.380 181.300 128.760 182.000 ;
    END
  END S2END[6]
  PIN S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 130.220 181.300 130.600 182.000 ;
    END
  END S2END[7]
  PIN S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.000 181.300 104.380 182.000 ;
    END
  END S2MID[0]
  PIN S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 105.840 181.300 106.220 182.000 ;
    END
  END S2MID[1]
  PIN S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 107.220 181.300 107.600 182.000 ;
    END
  END S2MID[2]
  PIN S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 109.060 181.300 109.440 182.000 ;
    END
  END S2MID[3]
  PIN S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.900 181.300 111.280 182.000 ;
    END
  END S2MID[4]
  PIN S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 112.740 181.300 113.120 182.000 ;
    END
  END S2MID[5]
  PIN S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 114.580 181.300 114.960 182.000 ;
    END
  END S2MID[6]
  PIN S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 116.420 181.300 116.800 182.000 ;
    END
  END S2MID[7]
  PIN S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 132.060 181.300 132.440 182.000 ;
    END
  END S4END[0]
  PIN S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 149.540 181.300 149.920 182.000 ;
    END
  END S4END[10]
  PIN S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 151.380 181.300 151.760 182.000 ;
    END
  END S4END[11]
  PIN S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.220 181.300 153.600 182.000 ;
    END
  END S4END[12]
  PIN S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.060 181.300 155.440 182.000 ;
    END
  END S4END[13]
  PIN S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.900 181.300 157.280 182.000 ;
    END
  END S4END[14]
  PIN S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.280 181.300 158.660 182.000 ;
    END
  END S4END[15]
  PIN S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 133.900 181.300 134.280 182.000 ;
    END
  END S4END[1]
  PIN S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 135.740 181.300 136.120 182.000 ;
    END
  END S4END[2]
  PIN S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.393000 ;
    PORT
      LAYER met2 ;
        RECT 137.120 181.300 137.500 182.000 ;
    END
  END S4END[3]
  PIN S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.960 181.300 139.340 182.000 ;
    END
  END S4END[4]
  PIN S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 140.800 181.300 141.180 182.000 ;
    END
  END S4END[5]
  PIN S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 142.640 181.300 143.020 182.000 ;
    END
  END S4END[6]
  PIN S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 144.480 181.300 144.860 182.000 ;
    END
  END S4END[7]
  PIN S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 146.320 181.300 146.700 182.000 ;
    END
  END S4END[8]
  PIN S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 147.700 181.300 148.080 182.000 ;
    END
  END S4END[9]
  PIN SS4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 160.120 181.300 160.500 182.000 ;
    END
  END SS4END[0]
  PIN SS4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.600 181.300 177.980 182.000 ;
    END
  END SS4END[10]
  PIN SS4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 179.440 181.300 179.820 182.000 ;
    END
  END SS4END[11]
  PIN SS4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 181.280 181.300 181.660 182.000 ;
    END
  END SS4END[12]
  PIN SS4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 183.120 181.300 183.500 182.000 ;
    END
  END SS4END[13]
  PIN SS4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 184.960 181.300 185.340 182.000 ;
    END
  END SS4END[14]
  PIN SS4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 186.800 181.300 187.180 182.000 ;
    END
  END SS4END[15]
  PIN SS4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.960 181.300 162.340 182.000 ;
    END
  END SS4END[1]
  PIN SS4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 163.800 181.300 164.180 182.000 ;
    END
  END SS4END[2]
  PIN SS4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.640 181.300 166.020 182.000 ;
    END
  END SS4END[3]
  PIN SS4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 167.480 181.300 167.860 182.000 ;
    END
  END SS4END[4]
  PIN SS4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 168.860 181.300 169.240 182.000 ;
    END
  END SS4END[5]
  PIN SS4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 170.700 181.300 171.080 182.000 ;
    END
  END SS4END[6]
  PIN SS4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 172.540 181.300 172.920 182.000 ;
    END
  END SS4END[7]
  PIN SS4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 174.380 181.300 174.760 182.000 ;
    END
  END SS4END[8]
  PIN SS4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 176.220 181.300 176.600 182.000 ;
    END
  END SS4END[9]
  PIN UIO_BOT_UIN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 154.140 0.000 154.520 0.700 ;
    END
  END UIO_BOT_UIN0
  PIN UIO_BOT_UIN1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 158.280 0.000 158.660 0.700 ;
    END
  END UIO_BOT_UIN1
  PIN UIO_BOT_UIN10
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.960 0.000 162.340 0.700 ;
    END
  END UIO_BOT_UIN10
  PIN UIO_BOT_UIN11
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 165.640 0.000 166.020 0.700 ;
    END
  END UIO_BOT_UIN11
  PIN UIO_BOT_UIN12
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 169.320 0.000 169.700 0.700 ;
    END
  END UIO_BOT_UIN12
  PIN UIO_BOT_UIN13
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 173.000 0.000 173.380 0.700 ;
    END
  END UIO_BOT_UIN13
  PIN UIO_BOT_UIN14
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 176.680 0.000 177.060 0.700 ;
    END
  END UIO_BOT_UIN14
  PIN UIO_BOT_UIN15
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 180.360 0.000 180.740 0.700 ;
    END
  END UIO_BOT_UIN15
  PIN UIO_BOT_UIN16
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 184.040 0.000 184.420 0.700 ;
    END
  END UIO_BOT_UIN16
  PIN UIO_BOT_UIN17
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 187.720 0.000 188.100 0.700 ;
    END
  END UIO_BOT_UIN17
  PIN UIO_BOT_UIN18
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.400 0.000 191.780 0.700 ;
    END
  END UIO_BOT_UIN18
  PIN UIO_BOT_UIN19
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.080 0.000 195.460 0.700 ;
    END
  END UIO_BOT_UIN19
  PIN UIO_BOT_UIN2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.760 0.000 199.140 0.700 ;
    END
  END UIO_BOT_UIN2
  PIN UIO_BOT_UIN3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 202.900 0.000 203.280 0.700 ;
    END
  END UIO_BOT_UIN3
  PIN UIO_BOT_UIN4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 206.580 0.000 206.960 0.700 ;
    END
  END UIO_BOT_UIN4
  PIN UIO_BOT_UIN5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 210.260 0.000 210.640 0.700 ;
    END
  END UIO_BOT_UIN5
  PIN UIO_BOT_UIN6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 213.940 0.000 214.320 0.700 ;
    END
  END UIO_BOT_UIN6
  PIN UIO_BOT_UIN7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.620 0.000 218.000 0.700 ;
    END
  END UIO_BOT_UIN7
  PIN UIO_BOT_UIN8
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 221.300 0.000 221.680 0.700 ;
    END
  END UIO_BOT_UIN8
  PIN UIO_BOT_UIN9
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 224.980 0.000 225.360 0.700 ;
    END
  END UIO_BOT_UIN9
  PIN UIO_BOT_UOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.080 0.000 80.460 0.700 ;
    END
  END UIO_BOT_UOUT0
  PIN UIO_BOT_UOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.760 0.000 84.140 0.700 ;
    END
  END UIO_BOT_UOUT1
  PIN UIO_BOT_UOUT10
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.440 0.000 87.820 0.700 ;
    END
  END UIO_BOT_UOUT10
  PIN UIO_BOT_UOUT11
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.120 0.000 91.500 0.700 ;
    END
  END UIO_BOT_UOUT11
  PIN UIO_BOT_UOUT12
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 94.800 0.000 95.180 0.700 ;
    END
  END UIO_BOT_UOUT12
  PIN UIO_BOT_UOUT13
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.480 0.000 98.860 0.700 ;
    END
  END UIO_BOT_UOUT13
  PIN UIO_BOT_UOUT14
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.160 0.000 102.540 0.700 ;
    END
  END UIO_BOT_UOUT14
  PIN UIO_BOT_UOUT15
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 105.840 0.000 106.220 0.700 ;
    END
  END UIO_BOT_UOUT15
  PIN UIO_BOT_UOUT16
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.520 0.000 109.900 0.700 ;
    END
  END UIO_BOT_UOUT16
  PIN UIO_BOT_UOUT17
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 113.200 0.000 113.580 0.700 ;
    END
  END UIO_BOT_UOUT17
  PIN UIO_BOT_UOUT18
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.340 0.000 117.720 0.700 ;
    END
  END UIO_BOT_UOUT18
  PIN UIO_BOT_UOUT19
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.020 0.000 121.400 0.700 ;
    END
  END UIO_BOT_UOUT19
  PIN UIO_BOT_UOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.700 0.000 125.080 0.700 ;
    END
  END UIO_BOT_UOUT2
  PIN UIO_BOT_UOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.380 0.000 128.760 0.700 ;
    END
  END UIO_BOT_UOUT3
  PIN UIO_BOT_UOUT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.060 0.000 132.440 0.700 ;
    END
  END UIO_BOT_UOUT4
  PIN UIO_BOT_UOUT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.740 0.000 136.120 0.700 ;
    END
  END UIO_BOT_UOUT5
  PIN UIO_BOT_UOUT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 139.420 0.000 139.800 0.700 ;
    END
  END UIO_BOT_UOUT6
  PIN UIO_BOT_UOUT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.100 0.000 143.480 0.700 ;
    END
  END UIO_BOT_UOUT7
  PIN UIO_BOT_UOUT8
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.780 0.000 147.160 0.700 ;
    END
  END UIO_BOT_UOUT8
  PIN UIO_BOT_UOUT9
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 150.460 0.000 150.840 0.700 ;
    END
  END UIO_BOT_UOUT9
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 0.700 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 0.700 ;
    END
  END UserCLKo
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -12.040 -11.660 -8.940 193.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 -11.660 242.960 -8.560 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.040 190.800 242.960 193.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 239.860 -11.660 242.960 193.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 20.580 -16.460 22.180 198.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 -16.460 175.780 198.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 21.290 247.760 22.890 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 174.470 247.760 176.070 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.840 -16.460 -13.740 198.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 -16.460 247.760 -13.360 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 195.600 247.760 198.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.660 -16.460 247.760 198.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.880 -16.460 25.480 198.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.480 -16.460 179.080 198.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.840 24.590 247.760 26.190 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 4.870 5.355 226.050 176.990 ;
      LAYER li1 ;
        RECT 5.060 5.355 225.860 176.885 ;
      LAYER met1 ;
        RECT 3.750 3.100 225.860 177.040 ;
      LAYER met2 ;
        RECT 4.380 181.020 5.280 181.300 ;
        RECT 6.220 181.020 6.660 181.300 ;
        RECT 7.600 181.020 8.500 181.300 ;
        RECT 9.440 181.020 10.340 181.300 ;
        RECT 11.280 181.020 12.180 181.300 ;
        RECT 13.120 181.020 14.020 181.300 ;
        RECT 14.960 181.020 15.400 181.300 ;
        RECT 16.340 181.020 17.240 181.300 ;
        RECT 18.180 181.020 19.080 181.300 ;
        RECT 20.020 181.020 20.920 181.300 ;
        RECT 21.860 181.020 22.760 181.300 ;
        RECT 23.700 181.020 24.600 181.300 ;
        RECT 25.540 181.020 25.980 181.300 ;
        RECT 26.920 181.020 27.820 181.300 ;
        RECT 28.760 181.020 29.660 181.300 ;
        RECT 30.600 181.020 31.500 181.300 ;
        RECT 32.440 181.020 33.340 181.300 ;
        RECT 34.280 181.020 35.180 181.300 ;
        RECT 36.120 181.020 36.560 181.300 ;
        RECT 37.500 181.020 38.400 181.300 ;
        RECT 39.340 181.020 40.240 181.300 ;
        RECT 41.180 181.020 42.080 181.300 ;
        RECT 43.020 181.020 43.920 181.300 ;
        RECT 44.860 181.020 45.760 181.300 ;
        RECT 46.700 181.020 47.140 181.300 ;
        RECT 48.080 181.020 48.980 181.300 ;
        RECT 49.920 181.020 50.820 181.300 ;
        RECT 51.760 181.020 52.660 181.300 ;
        RECT 53.600 181.020 54.500 181.300 ;
        RECT 55.440 181.020 55.880 181.300 ;
        RECT 56.820 181.020 57.720 181.300 ;
        RECT 58.660 181.020 59.560 181.300 ;
        RECT 60.500 181.020 61.400 181.300 ;
        RECT 62.340 181.020 63.240 181.300 ;
        RECT 64.180 181.020 65.080 181.300 ;
        RECT 66.020 181.020 66.460 181.300 ;
        RECT 67.400 181.020 68.300 181.300 ;
        RECT 69.240 181.020 70.140 181.300 ;
        RECT 71.080 181.020 71.980 181.300 ;
        RECT 72.920 181.020 73.820 181.300 ;
        RECT 74.760 181.020 75.660 181.300 ;
        RECT 76.600 181.020 77.040 181.300 ;
        RECT 77.980 181.020 78.880 181.300 ;
        RECT 79.820 181.020 80.720 181.300 ;
        RECT 81.660 181.020 82.560 181.300 ;
        RECT 83.500 181.020 84.400 181.300 ;
        RECT 85.340 181.020 86.240 181.300 ;
        RECT 87.180 181.020 87.620 181.300 ;
        RECT 88.560 181.020 89.460 181.300 ;
        RECT 90.400 181.020 91.300 181.300 ;
        RECT 92.240 181.020 93.140 181.300 ;
        RECT 94.080 181.020 94.980 181.300 ;
        RECT 95.920 181.020 96.360 181.300 ;
        RECT 97.300 181.020 98.200 181.300 ;
        RECT 99.140 181.020 100.040 181.300 ;
        RECT 100.980 181.020 101.880 181.300 ;
        RECT 102.820 181.020 103.720 181.300 ;
        RECT 104.660 181.020 105.560 181.300 ;
        RECT 106.500 181.020 106.940 181.300 ;
        RECT 107.880 181.020 108.780 181.300 ;
        RECT 109.720 181.020 110.620 181.300 ;
        RECT 111.560 181.020 112.460 181.300 ;
        RECT 113.400 181.020 114.300 181.300 ;
        RECT 115.240 181.020 116.140 181.300 ;
        RECT 117.080 181.020 117.520 181.300 ;
        RECT 118.460 181.020 119.360 181.300 ;
        RECT 120.300 181.020 121.200 181.300 ;
        RECT 122.140 181.020 123.040 181.300 ;
        RECT 123.980 181.020 124.880 181.300 ;
        RECT 125.820 181.020 126.720 181.300 ;
        RECT 127.660 181.020 128.100 181.300 ;
        RECT 129.040 181.020 129.940 181.300 ;
        RECT 130.880 181.020 131.780 181.300 ;
        RECT 132.720 181.020 133.620 181.300 ;
        RECT 134.560 181.020 135.460 181.300 ;
        RECT 136.400 181.020 136.840 181.300 ;
        RECT 137.780 181.020 138.680 181.300 ;
        RECT 139.620 181.020 140.520 181.300 ;
        RECT 141.460 181.020 142.360 181.300 ;
        RECT 143.300 181.020 144.200 181.300 ;
        RECT 145.140 181.020 146.040 181.300 ;
        RECT 146.980 181.020 147.420 181.300 ;
        RECT 148.360 181.020 149.260 181.300 ;
        RECT 150.200 181.020 151.100 181.300 ;
        RECT 152.040 181.020 152.940 181.300 ;
        RECT 153.880 181.020 154.780 181.300 ;
        RECT 155.720 181.020 156.620 181.300 ;
        RECT 157.560 181.020 158.000 181.300 ;
        RECT 158.940 181.020 159.840 181.300 ;
        RECT 160.780 181.020 161.680 181.300 ;
        RECT 162.620 181.020 163.520 181.300 ;
        RECT 164.460 181.020 165.360 181.300 ;
        RECT 166.300 181.020 167.200 181.300 ;
        RECT 168.140 181.020 168.580 181.300 ;
        RECT 169.520 181.020 170.420 181.300 ;
        RECT 171.360 181.020 172.260 181.300 ;
        RECT 173.200 181.020 174.100 181.300 ;
        RECT 175.040 181.020 175.940 181.300 ;
        RECT 176.880 181.020 177.320 181.300 ;
        RECT 178.260 181.020 179.160 181.300 ;
        RECT 180.100 181.020 181.000 181.300 ;
        RECT 181.940 181.020 182.840 181.300 ;
        RECT 183.780 181.020 184.680 181.300 ;
        RECT 185.620 181.020 186.520 181.300 ;
        RECT 187.460 181.020 187.900 181.300 ;
        RECT 188.840 181.020 189.740 181.300 ;
        RECT 190.680 181.020 191.580 181.300 ;
        RECT 192.520 181.020 193.420 181.300 ;
        RECT 194.360 181.020 195.260 181.300 ;
        RECT 196.200 181.020 197.100 181.300 ;
        RECT 198.040 181.020 198.480 181.300 ;
        RECT 199.420 181.020 200.320 181.300 ;
        RECT 201.260 181.020 202.160 181.300 ;
        RECT 203.100 181.020 204.000 181.300 ;
        RECT 204.940 181.020 205.840 181.300 ;
        RECT 206.780 181.020 207.680 181.300 ;
        RECT 208.620 181.020 209.060 181.300 ;
        RECT 210.000 181.020 210.900 181.300 ;
        RECT 211.840 181.020 212.740 181.300 ;
        RECT 213.680 181.020 214.580 181.300 ;
        RECT 215.520 181.020 216.420 181.300 ;
        RECT 217.360 181.020 217.800 181.300 ;
        RECT 218.740 181.020 219.640 181.300 ;
        RECT 220.580 181.020 221.480 181.300 ;
        RECT 222.420 181.020 225.300 181.300 ;
        RECT 3.780 0.980 225.300 181.020 ;
        RECT 3.780 0.270 5.280 0.980 ;
        RECT 6.220 0.270 8.960 0.980 ;
        RECT 9.900 0.270 12.640 0.980 ;
        RECT 13.580 0.270 16.320 0.980 ;
        RECT 17.260 0.270 20.000 0.980 ;
        RECT 20.940 0.270 23.680 0.980 ;
        RECT 24.620 0.270 27.360 0.980 ;
        RECT 28.300 0.270 31.500 0.980 ;
        RECT 32.440 0.270 35.180 0.980 ;
        RECT 36.120 0.270 38.860 0.980 ;
        RECT 39.800 0.270 42.540 0.980 ;
        RECT 43.480 0.270 46.220 0.980 ;
        RECT 47.160 0.270 49.900 0.980 ;
        RECT 50.840 0.270 53.580 0.980 ;
        RECT 54.520 0.270 57.260 0.980 ;
        RECT 58.200 0.270 60.940 0.980 ;
        RECT 61.880 0.270 64.620 0.980 ;
        RECT 65.560 0.270 68.300 0.980 ;
        RECT 69.240 0.270 72.440 0.980 ;
        RECT 73.380 0.270 76.120 0.980 ;
        RECT 77.060 0.270 79.800 0.980 ;
        RECT 80.740 0.270 83.480 0.980 ;
        RECT 84.420 0.270 87.160 0.980 ;
        RECT 88.100 0.270 90.840 0.980 ;
        RECT 91.780 0.270 94.520 0.980 ;
        RECT 95.460 0.270 98.200 0.980 ;
        RECT 99.140 0.270 99.630 0.980 ;
        RECT 100.470 0.270 101.880 0.980 ;
        RECT 102.820 0.270 102.850 0.980 ;
        RECT 103.690 0.270 105.560 0.980 ;
        RECT 106.500 0.270 109.240 0.980 ;
        RECT 110.180 0.270 112.920 0.980 ;
        RECT 113.860 0.270 117.060 0.980 ;
        RECT 118.000 0.270 120.740 0.980 ;
        RECT 121.680 0.270 124.420 0.980 ;
        RECT 125.360 0.270 128.100 0.980 ;
        RECT 129.040 0.270 131.780 0.980 ;
        RECT 132.720 0.270 135.460 0.980 ;
        RECT 136.400 0.270 139.140 0.980 ;
        RECT 140.080 0.270 142.820 0.980 ;
        RECT 143.760 0.270 146.500 0.980 ;
        RECT 147.440 0.270 150.180 0.980 ;
        RECT 151.120 0.270 153.860 0.980 ;
        RECT 154.800 0.270 158.000 0.980 ;
        RECT 158.940 0.270 161.680 0.980 ;
        RECT 162.620 0.270 165.360 0.980 ;
        RECT 166.300 0.270 169.040 0.980 ;
        RECT 169.980 0.270 172.720 0.980 ;
        RECT 173.660 0.270 176.400 0.980 ;
        RECT 177.340 0.270 180.080 0.980 ;
        RECT 181.020 0.270 183.760 0.980 ;
        RECT 184.700 0.270 187.440 0.980 ;
        RECT 188.380 0.270 191.120 0.980 ;
        RECT 192.060 0.270 194.800 0.980 ;
        RECT 195.740 0.270 198.480 0.980 ;
        RECT 199.420 0.270 202.620 0.980 ;
        RECT 203.560 0.270 206.300 0.980 ;
        RECT 207.240 0.270 209.980 0.980 ;
        RECT 210.920 0.270 213.660 0.980 ;
        RECT 214.600 0.270 217.340 0.980 ;
        RECT 218.280 0.270 221.020 0.980 ;
        RECT 221.960 0.270 224.700 0.980 ;
      LAYER met3 ;
        RECT 11.565 5.275 221.195 176.965 ;
      LAYER met4 ;
        RECT 101.495 6.295 128.505 173.225 ;
  END
END S_term_single
END LIBRARY

