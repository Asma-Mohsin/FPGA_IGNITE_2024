VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_IO
  CLASS BLOCK ;
  FOREIGN W_IO ;
  ORIGIN 0.000 0.000 ;
  SIZE 80.000 BY 223.115 ;
  PIN A_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 0.800 46.200 ;
    END
  END A_I_top
  PIN A_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 0.800 36.000 ;
    END
  END A_O_top
  PIN A_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 0.800 41.440 ;
    END
  END A_T_top
  PIN A_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 0.800 50.960 ;
    END
  END A_config_C_bit0
  PIN A_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 0.800 55.720 ;
    END
  END A_config_C_bit1
  PIN A_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 0.800 60.480 ;
    END
  END A_config_C_bit2
  PIN A_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 0.800 65.240 ;
    END
  END A_config_C_bit3
  PIN B_I_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 0.800 12.200 ;
    END
  END B_I_top
  PIN B_O_top
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 0.800 2.680 ;
    END
  END B_O_top
  PIN B_T_top
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 0.800 7.440 ;
    END
  END B_T_top
  PIN B_config_C_bit0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 0.800 16.960 ;
    END
  END B_config_C_bit0
  PIN B_config_C_bit1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 0.800 21.720 ;
    END
  END B_config_C_bit1
  PIN B_config_C_bit2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 0.800 26.480 ;
    END
  END B_config_C_bit2
  PIN B_config_C_bit3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 0.800 31.240 ;
    END
  END B_config_C_bit3
  PIN E1BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 84.360 80.000 84.960 ;
    END
  END E1BEG[0]
  PIN E1BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 85.720 80.000 86.320 ;
    END
  END E1BEG[1]
  PIN E1BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 87.760 80.000 88.360 ;
    END
  END E1BEG[2]
  PIN E1BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 89.120 80.000 89.720 ;
    END
  END E1BEG[3]
  PIN E2BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 91.160 80.000 91.760 ;
    END
  END E2BEG[0]
  PIN E2BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 92.520 80.000 93.120 ;
    END
  END E2BEG[1]
  PIN E2BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 94.560 80.000 95.160 ;
    END
  END E2BEG[2]
  PIN E2BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 95.920 80.000 96.520 ;
    END
  END E2BEG[3]
  PIN E2BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 97.960 80.000 98.560 ;
    END
  END E2BEG[4]
  PIN E2BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 100.000 80.000 100.600 ;
    END
  END E2BEG[5]
  PIN E2BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 101.360 80.000 101.960 ;
    END
  END E2BEG[6]
  PIN E2BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 103.400 80.000 104.000 ;
    END
  END E2BEG[7]
  PIN E2BEGb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 104.760 80.000 105.360 ;
    END
  END E2BEGb[0]
  PIN E2BEGb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 106.800 80.000 107.400 ;
    END
  END E2BEGb[1]
  PIN E2BEGb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 108.160 80.000 108.760 ;
    END
  END E2BEGb[2]
  PIN E2BEGb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 110.200 80.000 110.800 ;
    END
  END E2BEGb[3]
  PIN E2BEGb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 112.240 80.000 112.840 ;
    END
  END E2BEGb[4]
  PIN E2BEGb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 113.600 80.000 114.200 ;
    END
  END E2BEGb[5]
  PIN E2BEGb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 115.640 80.000 116.240 ;
    END
  END E2BEGb[6]
  PIN E2BEGb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 117.000 80.000 117.600 ;
    END
  END E2BEGb[7]
  PIN E6BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 146.920 80.000 147.520 ;
    END
  END E6BEG[0]
  PIN E6BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 163.920 80.000 164.520 ;
    END
  END E6BEG[10]
  PIN E6BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 165.960 80.000 166.560 ;
    END
  END E6BEG[11]
  PIN E6BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 148.280 80.000 148.880 ;
    END
  END E6BEG[1]
  PIN E6BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 150.320 80.000 150.920 ;
    END
  END E6BEG[2]
  PIN E6BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 151.680 80.000 152.280 ;
    END
  END E6BEG[3]
  PIN E6BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 153.720 80.000 154.320 ;
    END
  END E6BEG[4]
  PIN E6BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 155.760 80.000 156.360 ;
    END
  END E6BEG[5]
  PIN E6BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 157.120 80.000 157.720 ;
    END
  END E6BEG[6]
  PIN E6BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 159.160 80.000 159.760 ;
    END
  END E6BEG[7]
  PIN E6BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 160.520 80.000 161.120 ;
    END
  END E6BEG[8]
  PIN E6BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 162.560 80.000 163.160 ;
    END
  END E6BEG[9]
  PIN EE4BEG[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 119.040 80.000 119.640 ;
    END
  END EE4BEG[0]
  PIN EE4BEG[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 136.040 80.000 136.640 ;
    END
  END EE4BEG[10]
  PIN EE4BEG[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 138.080 80.000 138.680 ;
    END
  END EE4BEG[11]
  PIN EE4BEG[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 140.120 80.000 140.720 ;
    END
  END EE4BEG[12]
  PIN EE4BEG[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 141.480 80.000 142.080 ;
    END
  END EE4BEG[13]
  PIN EE4BEG[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 143.520 80.000 144.120 ;
    END
  END EE4BEG[14]
  PIN EE4BEG[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 144.880 80.000 145.480 ;
    END
  END EE4BEG[15]
  PIN EE4BEG[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 120.400 80.000 121.000 ;
    END
  END EE4BEG[1]
  PIN EE4BEG[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 122.440 80.000 123.040 ;
    END
  END EE4BEG[2]
  PIN EE4BEG[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 123.800 80.000 124.400 ;
    END
  END EE4BEG[3]
  PIN EE4BEG[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 125.840 80.000 126.440 ;
    END
  END EE4BEG[4]
  PIN EE4BEG[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 127.880 80.000 128.480 ;
    END
  END EE4BEG[5]
  PIN EE4BEG[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 129.240 80.000 129.840 ;
    END
  END EE4BEG[6]
  PIN EE4BEG[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 131.280 80.000 131.880 ;
    END
  END EE4BEG[7]
  PIN EE4BEG[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 132.640 80.000 133.240 ;
    END
  END EE4BEG[8]
  PIN EE4BEG[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 134.680 80.000 135.280 ;
    END
  END EE4BEG[9]
  PIN FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 0.800 70.000 ;
    END
  END FrameData[0]
  PIN FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 0.800 118.960 ;
    END
  END FrameData[10]
  PIN FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 0.800 123.720 ;
    END
  END FrameData[11]
  PIN FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 0.800 128.480 ;
    END
  END FrameData[12]
  PIN FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 0.800 133.240 ;
    END
  END FrameData[13]
  PIN FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 0.800 138.000 ;
    END
  END FrameData[14]
  PIN FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 0.800 142.760 ;
    END
  END FrameData[15]
  PIN FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 0.800 147.520 ;
    END
  END FrameData[16]
  PIN FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 0.800 152.960 ;
    END
  END FrameData[17]
  PIN FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 0.800 157.720 ;
    END
  END FrameData[18]
  PIN FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 0.800 162.480 ;
    END
  END FrameData[19]
  PIN FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.160 0.800 74.760 ;
    END
  END FrameData[1]
  PIN FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 0.800 167.240 ;
    END
  END FrameData[20]
  PIN FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 0.800 172.000 ;
    END
  END FrameData[21]
  PIN FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 0.800 176.760 ;
    END
  END FrameData[22]
  PIN FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 0.800 181.520 ;
    END
  END FrameData[23]
  PIN FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 0.800 186.280 ;
    END
  END FrameData[24]
  PIN FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 0.800 191.720 ;
    END
  END FrameData[25]
  PIN FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 0.800 196.480 ;
    END
  END FrameData[26]
  PIN FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 0.800 201.240 ;
    END
  END FrameData[27]
  PIN FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 0.800 206.000 ;
    END
  END FrameData[28]
  PIN FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.160 0.800 210.760 ;
    END
  END FrameData[29]
  PIN FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 0.800 80.200 ;
    END
  END FrameData[2]
  PIN FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 0.800 215.520 ;
    END
  END FrameData[30]
  PIN FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 0.800 220.280 ;
    END
  END FrameData[31]
  PIN FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 0.800 84.960 ;
    END
  END FrameData[3]
  PIN FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 0.800 89.720 ;
    END
  END FrameData[4]
  PIN FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 0.800 94.480 ;
    END
  END FrameData[5]
  PIN FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 0.800 99.240 ;
    END
  END FrameData[6]
  PIN FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 0.800 104.000 ;
    END
  END FrameData[7]
  PIN FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 0.800 108.760 ;
    END
  END FrameData[8]
  PIN FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 0.800 114.200 ;
    END
  END FrameData[9]
  PIN FrameData_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 168.000 80.000 168.600 ;
    END
  END FrameData_O[0]
  PIN FrameData_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 185.000 80.000 185.600 ;
    END
  END FrameData_O[10]
  PIN FrameData_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 187.040 80.000 187.640 ;
    END
  END FrameData_O[11]
  PIN FrameData_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 188.400 80.000 189.000 ;
    END
  END FrameData_O[12]
  PIN FrameData_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 190.440 80.000 191.040 ;
    END
  END FrameData_O[13]
  PIN FrameData_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 191.800 80.000 192.400 ;
    END
  END FrameData_O[14]
  PIN FrameData_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 193.840 80.000 194.440 ;
    END
  END FrameData_O[15]
  PIN FrameData_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 195.880 80.000 196.480 ;
    END
  END FrameData_O[16]
  PIN FrameData_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 197.240 80.000 197.840 ;
    END
  END FrameData_O[17]
  PIN FrameData_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 199.280 80.000 199.880 ;
    END
  END FrameData_O[18]
  PIN FrameData_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 200.640 80.000 201.240 ;
    END
  END FrameData_O[19]
  PIN FrameData_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 169.360 80.000 169.960 ;
    END
  END FrameData_O[1]
  PIN FrameData_O[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 202.680 80.000 203.280 ;
    END
  END FrameData_O[20]
  PIN FrameData_O[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 204.040 80.000 204.640 ;
    END
  END FrameData_O[21]
  PIN FrameData_O[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 206.080 80.000 206.680 ;
    END
  END FrameData_O[22]
  PIN FrameData_O[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 207.440 80.000 208.040 ;
    END
  END FrameData_O[23]
  PIN FrameData_O[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 209.480 80.000 210.080 ;
    END
  END FrameData_O[24]
  PIN FrameData_O[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 211.520 80.000 212.120 ;
    END
  END FrameData_O[25]
  PIN FrameData_O[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 212.880 80.000 213.480 ;
    END
  END FrameData_O[26]
  PIN FrameData_O[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 214.920 80.000 215.520 ;
    END
  END FrameData_O[27]
  PIN FrameData_O[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 216.280 80.000 216.880 ;
    END
  END FrameData_O[28]
  PIN FrameData_O[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 218.320 80.000 218.920 ;
    END
  END FrameData_O[29]
  PIN FrameData_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 171.400 80.000 172.000 ;
    END
  END FrameData_O[2]
  PIN FrameData_O[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 219.680 80.000 220.280 ;
    END
  END FrameData_O[30]
  PIN FrameData_O[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 221.720 80.000 222.320 ;
    END
  END FrameData_O[31]
  PIN FrameData_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 172.760 80.000 173.360 ;
    END
  END FrameData_O[3]
  PIN FrameData_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 174.800 80.000 175.400 ;
    END
  END FrameData_O[4]
  PIN FrameData_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 176.160 80.000 176.760 ;
    END
  END FrameData_O[5]
  PIN FrameData_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 178.200 80.000 178.800 ;
    END
  END FrameData_O[6]
  PIN FrameData_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 179.560 80.000 180.160 ;
    END
  END FrameData_O[7]
  PIN FrameData_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 181.600 80.000 182.200 ;
    END
  END FrameData_O[8]
  PIN FrameData_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 183.640 80.000 184.240 ;
    END
  END FrameData_O[9]
  PIN FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 0.000 5.890 0.800 ;
    END
  END FrameStrobe[0]
  PIN FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 0.800 ;
    END
  END FrameStrobe[10]
  PIN FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 0.800 ;
    END
  END FrameStrobe[11]
  PIN FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 0.800 ;
    END
  END FrameStrobe[12]
  PIN FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 0.800 ;
    END
  END FrameStrobe[13]
  PIN FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 0.800 ;
    END
  END FrameStrobe[14]
  PIN FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 0.800 ;
    END
  END FrameStrobe[15]
  PIN FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 0.800 ;
    END
  END FrameStrobe[16]
  PIN FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 0.800 ;
    END
  END FrameStrobe[17]
  PIN FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 0.800 ;
    END
  END FrameStrobe[18]
  PIN FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 0.800 ;
    END
  END FrameStrobe[19]
  PIN FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 0.800 ;
    END
  END FrameStrobe[1]
  PIN FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 0.800 ;
    END
  END FrameStrobe[2]
  PIN FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 0.800 ;
    END
  END FrameStrobe[3]
  PIN FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 0.800 ;
    END
  END FrameStrobe[4]
  PIN FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 0.800 ;
    END
  END FrameStrobe[5]
  PIN FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 0.800 ;
    END
  END FrameStrobe[6]
  PIN FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 0.800 ;
    END
  END FrameStrobe[7]
  PIN FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 0.800 ;
    END
  END FrameStrobe[8]
  PIN FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 0.800 ;
    END
  END FrameStrobe[9]
  PIN FrameStrobe_O[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 222.315 5.890 223.115 ;
    END
  END FrameStrobe_O[0]
  PIN FrameStrobe_O[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 222.315 44.070 223.115 ;
    END
  END FrameStrobe_O[10]
  PIN FrameStrobe_O[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.470 222.315 47.750 223.115 ;
    END
  END FrameStrobe_O[11]
  PIN FrameStrobe_O[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 222.315 51.430 223.115 ;
    END
  END FrameStrobe_O[12]
  PIN FrameStrobe_O[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 222.315 55.570 223.115 ;
    END
  END FrameStrobe_O[13]
  PIN FrameStrobe_O[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 222.315 59.250 223.115 ;
    END
  END FrameStrobe_O[14]
  PIN FrameStrobe_O[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 222.315 62.930 223.115 ;
    END
  END FrameStrobe_O[15]
  PIN FrameStrobe_O[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 222.315 66.610 223.115 ;
    END
  END FrameStrobe_O[16]
  PIN FrameStrobe_O[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 222.315 70.750 223.115 ;
    END
  END FrameStrobe_O[17]
  PIN FrameStrobe_O[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 222.315 74.430 223.115 ;
    END
  END FrameStrobe_O[18]
  PIN FrameStrobe_O[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 222.315 78.110 223.115 ;
    END
  END FrameStrobe_O[19]
  PIN FrameStrobe_O[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 222.315 9.570 223.115 ;
    END
  END FrameStrobe_O[1]
  PIN FrameStrobe_O[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 222.315 13.250 223.115 ;
    END
  END FrameStrobe_O[2]
  PIN FrameStrobe_O[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 222.315 17.390 223.115 ;
    END
  END FrameStrobe_O[3]
  PIN FrameStrobe_O[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 222.315 21.070 223.115 ;
    END
  END FrameStrobe_O[4]
  PIN FrameStrobe_O[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 222.315 24.750 223.115 ;
    END
  END FrameStrobe_O[5]
  PIN FrameStrobe_O[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 222.315 28.890 223.115 ;
    END
  END FrameStrobe_O[6]
  PIN FrameStrobe_O[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 222.315 32.570 223.115 ;
    END
  END FrameStrobe_O[7]
  PIN FrameStrobe_O[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 222.315 36.250 223.115 ;
    END
  END FrameStrobe_O[8]
  PIN FrameStrobe_O[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 222.315 39.930 223.115 ;
    END
  END FrameStrobe_O[9]
  PIN UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 0.800 ;
    END
  END UserCLK
  PIN UserCLKo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 222.315 2.210 223.115 ;
    END
  END UserCLKo
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 27.705 5.200 29.305 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.690 5.200 52.290 217.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.215 5.200 17.815 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.200 5.200 40.800 217.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.185 5.200 63.785 217.840 ;
    END
  END VPWR
  PIN W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 0.720 80.000 1.320 ;
    END
  END W1END[0]
  PIN W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 2.080 80.000 2.680 ;
    END
  END W1END[1]
  PIN W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 4.120 80.000 4.720 ;
    END
  END W1END[2]
  PIN W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 5.480 80.000 6.080 ;
    END
  END W1END[3]
  PIN W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 21.120 80.000 21.720 ;
    END
  END W2END[0]
  PIN W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 23.160 80.000 23.760 ;
    END
  END W2END[1]
  PIN W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 24.520 80.000 25.120 ;
    END
  END W2END[2]
  PIN W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 26.560 80.000 27.160 ;
    END
  END W2END[3]
  PIN W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 28.600 80.000 29.200 ;
    END
  END W2END[4]
  PIN W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 29.960 80.000 30.560 ;
    END
  END W2END[5]
  PIN W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 32.000 80.000 32.600 ;
    END
  END W2END[6]
  PIN W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 33.360 80.000 33.960 ;
    END
  END W2END[7]
  PIN W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 7.520 80.000 8.120 ;
    END
  END W2MID[0]
  PIN W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 8.880 80.000 9.480 ;
    END
  END W2MID[1]
  PIN W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 10.920 80.000 11.520 ;
    END
  END W2MID[2]
  PIN W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 12.280 80.000 12.880 ;
    END
  END W2MID[3]
  PIN W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 14.320 80.000 14.920 ;
    END
  END W2MID[4]
  PIN W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 16.360 80.000 16.960 ;
    END
  END W2MID[5]
  PIN W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 17.720 80.000 18.320 ;
    END
  END W2MID[6]
  PIN W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 19.760 80.000 20.360 ;
    END
  END W2MID[7]
  PIN W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 63.280 80.000 63.880 ;
    END
  END W6END[0]
  PIN W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 80.280 80.000 80.880 ;
    END
  END W6END[10]
  PIN W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 82.320 80.000 82.920 ;
    END
  END W6END[11]
  PIN W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 64.640 80.000 65.240 ;
    END
  END W6END[1]
  PIN W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 66.680 80.000 67.280 ;
    END
  END W6END[2]
  PIN W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 68.040 80.000 68.640 ;
    END
  END W6END[3]
  PIN W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 70.080 80.000 70.680 ;
    END
  END W6END[4]
  PIN W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 72.120 80.000 72.720 ;
    END
  END W6END[5]
  PIN W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 73.480 80.000 74.080 ;
    END
  END W6END[6]
  PIN W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 75.520 80.000 76.120 ;
    END
  END W6END[7]
  PIN W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 76.880 80.000 77.480 ;
    END
  END W6END[8]
  PIN W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 78.920 80.000 79.520 ;
    END
  END W6END[9]
  PIN WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 35.400 80.000 36.000 ;
    END
  END WW4END[0]
  PIN WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 52.400 80.000 53.000 ;
    END
  END WW4END[10]
  PIN WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 54.440 80.000 55.040 ;
    END
  END WW4END[11]
  PIN WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 56.480 80.000 57.080 ;
    END
  END WW4END[12]
  PIN WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 57.840 80.000 58.440 ;
    END
  END WW4END[13]
  PIN WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 59.880 80.000 60.480 ;
    END
  END WW4END[14]
  PIN WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 61.240 80.000 61.840 ;
    END
  END WW4END[15]
  PIN WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 36.760 80.000 37.360 ;
    END
  END WW4END[1]
  PIN WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 38.800 80.000 39.400 ;
    END
  END WW4END[2]
  PIN WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 40.160 80.000 40.760 ;
    END
  END WW4END[3]
  PIN WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 42.200 80.000 42.800 ;
    END
  END WW4END[4]
  PIN WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 44.240 80.000 44.840 ;
    END
  END WW4END[5]
  PIN WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 45.600 80.000 46.200 ;
    END
  END WW4END[6]
  PIN WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 47.640 80.000 48.240 ;
    END
  END WW4END[7]
  PIN WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 49.000 80.000 49.600 ;
    END
  END WW4END[8]
  PIN WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 79.200 51.040 80.000 51.640 ;
    END
  END WW4END[9]
  OBS
      LAYER li1 ;
        RECT 5.520 2.465 79.895 217.685 ;
      LAYER met1 ;
        RECT 1.910 2.080 79.970 218.920 ;
      LAYER met2 ;
        RECT 2.490 222.035 5.330 222.770 ;
        RECT 6.170 222.035 9.010 222.770 ;
        RECT 9.850 222.035 12.690 222.770 ;
        RECT 13.530 222.035 16.830 222.770 ;
        RECT 17.670 222.035 20.510 222.770 ;
        RECT 21.350 222.035 24.190 222.770 ;
        RECT 25.030 222.035 28.330 222.770 ;
        RECT 29.170 222.035 32.010 222.770 ;
        RECT 32.850 222.035 35.690 222.770 ;
        RECT 36.530 222.035 39.370 222.770 ;
        RECT 40.210 222.035 43.510 222.770 ;
        RECT 44.350 222.035 47.190 222.770 ;
        RECT 48.030 222.035 50.870 222.770 ;
        RECT 51.710 222.035 55.010 222.770 ;
        RECT 55.850 222.035 58.690 222.770 ;
        RECT 59.530 222.035 62.370 222.770 ;
        RECT 63.210 222.035 66.050 222.770 ;
        RECT 66.890 222.035 70.190 222.770 ;
        RECT 71.030 222.035 73.870 222.770 ;
        RECT 74.710 222.035 77.550 222.770 ;
        RECT 78.390 222.035 79.940 222.770 ;
        RECT 1.940 1.080 79.940 222.035 ;
        RECT 2.490 0.270 5.330 1.080 ;
        RECT 6.170 0.270 9.010 1.080 ;
        RECT 9.850 0.270 12.690 1.080 ;
        RECT 13.530 0.270 16.830 1.080 ;
        RECT 17.670 0.270 20.510 1.080 ;
        RECT 21.350 0.270 24.190 1.080 ;
        RECT 25.030 0.270 28.330 1.080 ;
        RECT 29.170 0.270 32.010 1.080 ;
        RECT 32.850 0.270 35.690 1.080 ;
        RECT 36.530 0.270 39.370 1.080 ;
        RECT 40.210 0.270 43.510 1.080 ;
        RECT 44.350 0.270 47.190 1.080 ;
        RECT 48.030 0.270 50.870 1.080 ;
        RECT 51.710 0.270 55.010 1.080 ;
        RECT 55.850 0.270 58.690 1.080 ;
        RECT 59.530 0.270 62.370 1.080 ;
        RECT 63.210 0.270 66.050 1.080 ;
        RECT 66.890 0.270 70.190 1.080 ;
        RECT 71.030 0.270 73.870 1.080 ;
        RECT 74.710 0.270 77.550 1.080 ;
        RECT 78.390 0.270 79.940 1.080 ;
      LAYER met3 ;
        RECT 0.800 221.320 78.800 222.185 ;
        RECT 0.800 220.680 79.200 221.320 ;
        RECT 1.200 219.280 78.800 220.680 ;
        RECT 0.800 217.920 78.800 219.280 ;
        RECT 0.800 217.280 79.200 217.920 ;
        RECT 0.800 215.920 78.800 217.280 ;
        RECT 1.200 214.520 78.800 215.920 ;
        RECT 0.800 213.880 79.200 214.520 ;
        RECT 0.800 211.160 78.800 213.880 ;
        RECT 1.200 211.120 78.800 211.160 ;
        RECT 1.200 210.480 79.200 211.120 ;
        RECT 1.200 209.760 78.800 210.480 ;
        RECT 0.800 209.080 78.800 209.760 ;
        RECT 0.800 208.440 79.200 209.080 ;
        RECT 0.800 206.400 78.800 208.440 ;
        RECT 1.200 205.680 78.800 206.400 ;
        RECT 1.200 205.040 79.200 205.680 ;
        RECT 1.200 205.000 78.800 205.040 ;
        RECT 0.800 202.280 78.800 205.000 ;
        RECT 0.800 201.640 79.200 202.280 ;
        RECT 1.200 200.240 78.800 201.640 ;
        RECT 0.800 198.880 78.800 200.240 ;
        RECT 0.800 198.240 79.200 198.880 ;
        RECT 0.800 196.880 78.800 198.240 ;
        RECT 1.200 195.480 78.800 196.880 ;
        RECT 0.800 194.840 79.200 195.480 ;
        RECT 0.800 193.440 78.800 194.840 ;
        RECT 0.800 192.800 79.200 193.440 ;
        RECT 0.800 192.120 78.800 192.800 ;
        RECT 1.200 190.720 78.800 192.120 ;
        RECT 0.800 190.040 78.800 190.720 ;
        RECT 0.800 189.400 79.200 190.040 ;
        RECT 0.800 186.680 78.800 189.400 ;
        RECT 1.200 186.640 78.800 186.680 ;
        RECT 1.200 186.000 79.200 186.640 ;
        RECT 1.200 185.280 78.800 186.000 ;
        RECT 0.800 183.240 78.800 185.280 ;
        RECT 0.800 182.600 79.200 183.240 ;
        RECT 0.800 181.920 78.800 182.600 ;
        RECT 1.200 181.200 78.800 181.920 ;
        RECT 1.200 180.560 79.200 181.200 ;
        RECT 1.200 180.520 78.800 180.560 ;
        RECT 0.800 177.800 78.800 180.520 ;
        RECT 0.800 177.160 79.200 177.800 ;
        RECT 1.200 175.760 78.800 177.160 ;
        RECT 0.800 174.400 78.800 175.760 ;
        RECT 0.800 173.760 79.200 174.400 ;
        RECT 0.800 172.400 78.800 173.760 ;
        RECT 1.200 171.000 78.800 172.400 ;
        RECT 0.800 170.360 79.200 171.000 ;
        RECT 0.800 167.640 78.800 170.360 ;
        RECT 1.200 167.600 78.800 167.640 ;
        RECT 1.200 166.960 79.200 167.600 ;
        RECT 1.200 166.240 78.800 166.960 ;
        RECT 0.800 165.560 78.800 166.240 ;
        RECT 0.800 164.920 79.200 165.560 ;
        RECT 0.800 162.880 78.800 164.920 ;
        RECT 1.200 162.160 78.800 162.880 ;
        RECT 1.200 161.520 79.200 162.160 ;
        RECT 1.200 161.480 78.800 161.520 ;
        RECT 0.800 158.760 78.800 161.480 ;
        RECT 0.800 158.120 79.200 158.760 ;
        RECT 1.200 156.720 78.800 158.120 ;
        RECT 0.800 155.360 78.800 156.720 ;
        RECT 0.800 154.720 79.200 155.360 ;
        RECT 0.800 153.360 78.800 154.720 ;
        RECT 1.200 153.320 78.800 153.360 ;
        RECT 1.200 152.680 79.200 153.320 ;
        RECT 1.200 151.960 78.800 152.680 ;
        RECT 0.800 149.920 78.800 151.960 ;
        RECT 0.800 149.280 79.200 149.920 ;
        RECT 0.800 147.920 78.800 149.280 ;
        RECT 1.200 146.520 78.800 147.920 ;
        RECT 0.800 145.880 79.200 146.520 ;
        RECT 0.800 143.160 78.800 145.880 ;
        RECT 1.200 143.120 78.800 143.160 ;
        RECT 1.200 142.480 79.200 143.120 ;
        RECT 1.200 141.760 78.800 142.480 ;
        RECT 0.800 139.720 78.800 141.760 ;
        RECT 0.800 139.080 79.200 139.720 ;
        RECT 0.800 138.400 78.800 139.080 ;
        RECT 1.200 137.680 78.800 138.400 ;
        RECT 1.200 137.040 79.200 137.680 ;
        RECT 1.200 137.000 78.800 137.040 ;
        RECT 0.800 134.280 78.800 137.000 ;
        RECT 0.800 133.640 79.200 134.280 ;
        RECT 1.200 132.240 78.800 133.640 ;
        RECT 0.800 130.880 78.800 132.240 ;
        RECT 0.800 130.240 79.200 130.880 ;
        RECT 0.800 128.880 78.800 130.240 ;
        RECT 1.200 127.480 78.800 128.880 ;
        RECT 0.800 126.840 79.200 127.480 ;
        RECT 0.800 125.440 78.800 126.840 ;
        RECT 0.800 124.800 79.200 125.440 ;
        RECT 0.800 124.120 78.800 124.800 ;
        RECT 1.200 122.720 78.800 124.120 ;
        RECT 0.800 122.040 78.800 122.720 ;
        RECT 0.800 121.400 79.200 122.040 ;
        RECT 0.800 119.360 78.800 121.400 ;
        RECT 1.200 118.640 78.800 119.360 ;
        RECT 1.200 118.000 79.200 118.640 ;
        RECT 1.200 117.960 78.800 118.000 ;
        RECT 0.800 115.240 78.800 117.960 ;
        RECT 0.800 114.600 79.200 115.240 ;
        RECT 1.200 113.200 78.800 114.600 ;
        RECT 0.800 111.840 78.800 113.200 ;
        RECT 0.800 111.200 79.200 111.840 ;
        RECT 0.800 109.800 78.800 111.200 ;
        RECT 0.800 109.160 79.200 109.800 ;
        RECT 1.200 107.760 78.800 109.160 ;
        RECT 0.800 106.400 78.800 107.760 ;
        RECT 0.800 105.760 79.200 106.400 ;
        RECT 0.800 104.400 78.800 105.760 ;
        RECT 1.200 103.000 78.800 104.400 ;
        RECT 0.800 102.360 79.200 103.000 ;
        RECT 0.800 99.640 78.800 102.360 ;
        RECT 1.200 99.600 78.800 99.640 ;
        RECT 1.200 98.960 79.200 99.600 ;
        RECT 1.200 98.240 78.800 98.960 ;
        RECT 0.800 97.560 78.800 98.240 ;
        RECT 0.800 96.920 79.200 97.560 ;
        RECT 0.800 94.880 78.800 96.920 ;
        RECT 1.200 94.160 78.800 94.880 ;
        RECT 1.200 93.520 79.200 94.160 ;
        RECT 1.200 93.480 78.800 93.520 ;
        RECT 0.800 90.760 78.800 93.480 ;
        RECT 0.800 90.120 79.200 90.760 ;
        RECT 1.200 88.720 78.800 90.120 ;
        RECT 0.800 87.360 78.800 88.720 ;
        RECT 0.800 86.720 79.200 87.360 ;
        RECT 0.800 85.360 78.800 86.720 ;
        RECT 1.200 83.960 78.800 85.360 ;
        RECT 0.800 83.320 79.200 83.960 ;
        RECT 0.800 81.920 78.800 83.320 ;
        RECT 0.800 81.280 79.200 81.920 ;
        RECT 0.800 80.600 78.800 81.280 ;
        RECT 1.200 79.200 78.800 80.600 ;
        RECT 0.800 78.520 78.800 79.200 ;
        RECT 0.800 77.880 79.200 78.520 ;
        RECT 0.800 75.160 78.800 77.880 ;
        RECT 1.200 75.120 78.800 75.160 ;
        RECT 1.200 74.480 79.200 75.120 ;
        RECT 1.200 73.760 78.800 74.480 ;
        RECT 0.800 71.720 78.800 73.760 ;
        RECT 0.800 71.080 79.200 71.720 ;
        RECT 0.800 70.400 78.800 71.080 ;
        RECT 1.200 69.680 78.800 70.400 ;
        RECT 1.200 69.040 79.200 69.680 ;
        RECT 1.200 69.000 78.800 69.040 ;
        RECT 0.800 66.280 78.800 69.000 ;
        RECT 0.800 65.640 79.200 66.280 ;
        RECT 1.200 64.240 78.800 65.640 ;
        RECT 0.800 62.880 78.800 64.240 ;
        RECT 0.800 62.240 79.200 62.880 ;
        RECT 0.800 60.880 78.800 62.240 ;
        RECT 1.200 59.480 78.800 60.880 ;
        RECT 0.800 58.840 79.200 59.480 ;
        RECT 0.800 56.120 78.800 58.840 ;
        RECT 1.200 56.080 78.800 56.120 ;
        RECT 1.200 55.440 79.200 56.080 ;
        RECT 1.200 54.720 78.800 55.440 ;
        RECT 0.800 54.040 78.800 54.720 ;
        RECT 0.800 53.400 79.200 54.040 ;
        RECT 0.800 51.360 78.800 53.400 ;
        RECT 1.200 50.640 78.800 51.360 ;
        RECT 1.200 50.000 79.200 50.640 ;
        RECT 1.200 49.960 78.800 50.000 ;
        RECT 0.800 47.240 78.800 49.960 ;
        RECT 0.800 46.600 79.200 47.240 ;
        RECT 1.200 45.200 78.800 46.600 ;
        RECT 0.800 43.840 78.800 45.200 ;
        RECT 0.800 43.200 79.200 43.840 ;
        RECT 0.800 41.840 78.800 43.200 ;
        RECT 1.200 41.800 78.800 41.840 ;
        RECT 1.200 41.160 79.200 41.800 ;
        RECT 1.200 40.440 78.800 41.160 ;
        RECT 0.800 38.400 78.800 40.440 ;
        RECT 0.800 37.760 79.200 38.400 ;
        RECT 0.800 36.400 78.800 37.760 ;
        RECT 1.200 35.000 78.800 36.400 ;
        RECT 0.800 34.360 79.200 35.000 ;
        RECT 0.800 31.640 78.800 34.360 ;
        RECT 1.200 31.600 78.800 31.640 ;
        RECT 1.200 30.960 79.200 31.600 ;
        RECT 1.200 30.240 78.800 30.960 ;
        RECT 0.800 28.200 78.800 30.240 ;
        RECT 0.800 27.560 79.200 28.200 ;
        RECT 0.800 26.880 78.800 27.560 ;
        RECT 1.200 26.160 78.800 26.880 ;
        RECT 1.200 25.520 79.200 26.160 ;
        RECT 1.200 25.480 78.800 25.520 ;
        RECT 0.800 22.760 78.800 25.480 ;
        RECT 0.800 22.120 79.200 22.760 ;
        RECT 1.200 20.720 78.800 22.120 ;
        RECT 0.800 19.360 78.800 20.720 ;
        RECT 0.800 18.720 79.200 19.360 ;
        RECT 0.800 17.360 78.800 18.720 ;
        RECT 1.200 15.960 78.800 17.360 ;
        RECT 0.800 15.320 79.200 15.960 ;
        RECT 0.800 13.920 78.800 15.320 ;
        RECT 0.800 13.280 79.200 13.920 ;
        RECT 0.800 12.600 78.800 13.280 ;
        RECT 1.200 11.200 78.800 12.600 ;
        RECT 0.800 10.520 78.800 11.200 ;
        RECT 0.800 9.880 79.200 10.520 ;
        RECT 0.800 7.840 78.800 9.880 ;
        RECT 1.200 7.120 78.800 7.840 ;
        RECT 1.200 6.480 79.200 7.120 ;
        RECT 1.200 6.440 78.800 6.480 ;
        RECT 0.800 3.720 78.800 6.440 ;
        RECT 0.800 3.080 79.200 3.720 ;
        RECT 1.200 1.680 78.800 3.080 ;
        RECT 0.800 0.855 78.800 1.680 ;
      LAYER met4 ;
        RECT 18.215 5.200 27.305 217.840 ;
        RECT 29.705 5.200 38.800 217.840 ;
        RECT 41.200 5.200 50.290 217.840 ;
        RECT 52.690 5.200 61.785 217.840 ;
        RECT 64.185 5.200 67.785 217.840 ;
  END
END W_IO
END LIBRARY

