`timescale 1ns/1ps
module User_project_IO(UIN0, UIN1, UIN2, UIN3, UIN4, UIN5, UIN6, UIN7, UIN8, UIN9, UIN10, UIN11, UIN12, UIN13, UIN14, UIN15, UIN16, UIN17, UIN18, UIN19, UOUT0, UOUT1, UOUT2, UOUT3, UOUT4, UOUT5, UOUT6, UOUT7, UOUT8, UOUT9, UOUT10, UOUT11, UOUT12, UOUT13, UOUT14, UOUT15, UOUT16, UOUT17, UOUT18, UOUT19, FIN0, FIN1, FIN2, FIN3, FIN4, FIN5, FIN6, FIN7, FIN8, FIN9, FIN10, FIN11, FIN12, FIN13, FIN14, FIN15, FIN16, FIN17, FIN18, FIN19, FOUT0, FOUT1, FOUT2, FOUT3, FOUT4, FOUT5, FOUT6, FOUT7, FOUT8, FOUT9, FOUT10, FOUT11, FOUT12, FOUT13, FOUT14, FOUT15, FOUT16, FOUT17, FOUT18, FOUT19);
(* FABulous, EXTERNAL *) input UIN0; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT0; // EXTERNAL
input FIN0;
output FOUT0;
(* FABulous, EXTERNAL *) input UIN1; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT1; // EXTERNAL
input FIN1;
output FOUT1;
(* FABulous, EXTERNAL *) input UIN2; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT2; // EXTERNAL
input FIN2;
output FOUT2;
(* FABulous, EXTERNAL *) input UIN3; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT3; // EXTERNAL
input FIN3;
output FOUT3;
(* FABulous, EXTERNAL *) input UIN4; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT4; // EXTERNAL
input FIN4;
output FOUT4;
(* FABulous, EXTERNAL *) input UIN5; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT5; // EXTERNAL
input FIN5;
output FOUT5;
(* FABulous, EXTERNAL *) input UIN6; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT6; // EXTERNAL
input FIN6;
output FOUT6;
(* FABulous, EXTERNAL *) input UIN7; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT7; // EXTERNAL
input FIN7;
output FOUT7;
(* FABulous, EXTERNAL *) input UIN8; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT8; // EXTERNAL
input FIN8;
output FOUT8;
(* FABulous, EXTERNAL *) input UIN9; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT9; // EXTERNAL
input FIN9;
output FOUT9;
(* FABulous, EXTERNAL *) input UIN10; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT10; // EXTERNAL
input FIN10;
output FOUT10;
(* FABulous, EXTERNAL *) input UIN11; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT11; // EXTERNAL
input FIN11;
output FOUT11;
(* FABulous, EXTERNAL *) input UIN12; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT12; // EXTERNAL
input FIN12;
output FOUT12;
(* FABulous, EXTERNAL *) input UIN13; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT13; // EXTERNAL
input FIN13;
output FOUT13;
(* FABulous, EXTERNAL *) input UIN14; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT14; // EXTERNAL
input FIN14;
output FOUT14;
(* FABulous, EXTERNAL *) input UIN15; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT15; // EXTERNAL
input FIN15;
output FOUT15;
(* FABulous, EXTERNAL *) input UIN16; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT16; // EXTERNAL
input FIN16;
output FOUT16;
(* FABulous, EXTERNAL *) input UIN17; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT17; // EXTERNAL
input FIN17;
output FOUT17;
(* FABulous, EXTERNAL *) input UIN18; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT18; // EXTERNAL
input FIN18;
output FOUT18;
(* FABulous, EXTERNAL *) input UIN19; // EXTERNAL
(* FABulous, EXTERNAL *) output UOUT19; // EXTERNAL
input FIN19;
output FOUT19;
   assign UOUT0 = FIN0;
   assign FOUT0 = UIN0;
   assign UOUT1 = FIN1;
   assign FOUT1 = UIN1;
   assign UOUT2 = FIN2;
   assign FOUT2 = UIN2;
   assign UOUT3 = FIN3;
   assign FOUT3 = UIN3;
   assign UOUT4 = FIN4;
   assign FOUT4 = UIN4;
   assign UOUT5 = FIN5;
   assign FOUT5 = UIN5;
   assign UOUT6 = FIN6;
   assign FOUT6 = UIN6;
   assign UOUT7 = FIN7;
   assign FOUT7 = UIN7;
   assign UOUT8 = FIN8;
   assign FOUT8 = UIN8;
   assign UOUT9 = FIN9;
   assign FOUT9 = UIN9;
   assign UOUT10 = FIN10;
   assign FOUT10 = UIN10;
   assign UOUT11 = FIN11;
   assign FOUT11 = UIN11;
   assign UOUT12 = FIN12;
   assign FOUT12 = UIN12;
   assign UOUT13 = FIN13;
   assign FOUT13 = UIN13;
   assign UOUT14 = FIN14;
   assign FOUT14 = UIN14;
   assign UOUT15 = FIN15;
   assign FOUT15 = UIN15;
   assign UOUT16 = FIN16;
   assign FOUT16 = UIN16;
   assign UOUT17 = FIN17;
   assign FOUT17 = UIN17;
   assign UOUT18 = FIN18;
   assign FOUT18 = UIN18;
   assign UOUT19 = FIN19;
   assign FOUT19 = UIN19;
endmodule
